
module addr_sel ( clk, addr_serial_num, sram_raddr_w0, sram_raddr_w1, 
        sram_raddr_d0, sram_raddr_d1 );
  input [6:0] addr_serial_num;
  output [9:0] sram_raddr_w0;
  output [9:0] sram_raddr_w1;
  output [9:0] sram_raddr_d0;
  output [9:0] sram_raddr_d1;
  input clk;
  wire   sram_raddr_w0_nx_4_, sram_raddr_w0_nx_3_, sram_raddr_w0_nx_2_, N9,
         N10, N11, N12, N13, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68;
  wire   [6:0] sram_raddr_w1_nx;
  wire   [6:4] sub_34_carry;

  DFF_X1 sram_raddr_w0_reg_6_ ( .D(n32), .CK(clk), .Q(sram_raddr_w0[6]) );
  DFF_X1 sram_raddr_w0_reg_5_ ( .D(n36), .CK(clk), .Q(sram_raddr_w0[5]) );
  DFF_X1 sram_raddr_w0_reg_4_ ( .D(sram_raddr_w0_nx_4_), .CK(clk), .Q(
        sram_raddr_w0[4]) );
  DFF_X1 sram_raddr_w0_reg_3_ ( .D(sram_raddr_w0_nx_3_), .CK(clk), .Q(
        sram_raddr_w0[3]) );
  DFF_X1 sram_raddr_w0_reg_2_ ( .D(sram_raddr_w0_nx_2_), .CK(clk), .Q(
        sram_raddr_w0[2]) );
  DFF_X1 sram_raddr_w1_reg_6_ ( .D(sram_raddr_w1_nx[6]), .CK(clk), .Q(
        sram_raddr_w1[6]) );
  DFF_X1 sram_raddr_w1_reg_5_ ( .D(sram_raddr_w1_nx[5]), .CK(clk), .Q(
        sram_raddr_w1[5]) );
  DFF_X1 sram_raddr_w1_reg_4_ ( .D(sram_raddr_w1_nx[4]), .CK(clk), .Q(
        sram_raddr_w1[4]) );
  DFF_X1 sram_raddr_w1_reg_3_ ( .D(sram_raddr_w1_nx[3]), .CK(clk), .Q(
        sram_raddr_w1[3]) );
  DFF_X1 sram_raddr_w1_reg_2_ ( .D(sram_raddr_w1_nx[2]), .CK(clk), .Q(
        sram_raddr_w1[2]) );
  DFF_X1 sram_raddr_w1_reg_1_ ( .D(sram_raddr_w1_nx[1]), .CK(clk), .Q(
        sram_raddr_w1[1]) );
  DFF_X1 sram_raddr_w1_reg_0_ ( .D(sram_raddr_w1_nx[0]), .CK(clk), .Q(
        sram_raddr_w1[0]) );
  DFF_X1 sram_raddr_d0_reg_6_ ( .D(n30), .CK(clk), .Q(sram_raddr_d0[6]) );
  DFF_X1 sram_raddr_d0_reg_5_ ( .D(n34), .CK(clk), .Q(sram_raddr_d0[5]) );
  DFF_X1 sram_raddr_d0_reg_4_ ( .D(sram_raddr_w0_nx_4_), .CK(clk), .Q(
        sram_raddr_d0[4]) );
  DFF_X1 sram_raddr_d0_reg_3_ ( .D(sram_raddr_w0_nx_3_), .CK(clk), .Q(
        sram_raddr_d0[3]) );
  DFF_X1 sram_raddr_d0_reg_2_ ( .D(sram_raddr_w0_nx_2_), .CK(clk), .Q(
        sram_raddr_d0[2]) );
  DFF_X1 sram_raddr_d1_reg_6_ ( .D(sram_raddr_w1_nx[6]), .CK(clk), .Q(
        sram_raddr_d1[6]) );
  DFF_X1 sram_raddr_d1_reg_5_ ( .D(sram_raddr_w1_nx[5]), .CK(clk), .Q(
        sram_raddr_d1[5]) );
  DFF_X1 sram_raddr_d1_reg_4_ ( .D(sram_raddr_w1_nx[4]), .CK(clk), .Q(
        sram_raddr_d1[4]) );
  DFF_X1 sram_raddr_d1_reg_3_ ( .D(sram_raddr_w1_nx[3]), .CK(clk), .Q(
        sram_raddr_d1[3]) );
  DFF_X1 sram_raddr_d1_reg_2_ ( .D(sram_raddr_w1_nx[2]), .CK(clk), .Q(
        sram_raddr_d1[2]) );
  DFF_X1 sram_raddr_d1_reg_1_ ( .D(sram_raddr_w1_nx[1]), .CK(clk), .Q(
        sram_raddr_d1[1]) );
  DFF_X1 sram_raddr_d1_reg_0_ ( .D(sram_raddr_w1_nx[0]), .CK(clk), .Q(
        sram_raddr_d1[0]) );
  DFF_X1 sram_raddr_w0_reg_1_ ( .D(n55), .CK(clk), .Q(sram_raddr_w0[1]) );
  DFF_X1 sram_raddr_w0_reg_0_ ( .D(n54), .CK(clk), .Q(sram_raddr_w0[0]) );
  DFF_X1 sram_raddr_d0_reg_1_ ( .D(n55), .CK(clk), .Q(sram_raddr_d0[1]) );
  DFF_X1 sram_raddr_d0_reg_0_ ( .D(n54), .CK(clk), .Q(sram_raddr_d0[0]) );
  INV_X1 U6 ( .A(1'b1), .ZN(sram_raddr_d1[7]) );
  INV_X1 U8 ( .A(1'b1), .ZN(sram_raddr_d1[8]) );
  INV_X1 U10 ( .A(1'b1), .ZN(sram_raddr_d1[9]) );
  INV_X1 U12 ( .A(1'b1), .ZN(sram_raddr_d0[7]) );
  INV_X1 U20 ( .A(1'b1), .ZN(sram_raddr_d0[8]) );
  INV_X1 U25 ( .A(1'b1), .ZN(sram_raddr_d0[9]) );
  INV_X1 U27 ( .A(1'b1), .ZN(sram_raddr_w1[7]) );
  INV_X1 U29 ( .A(1'b1), .ZN(sram_raddr_w1[8]) );
  INV_X1 U31 ( .A(1'b1), .ZN(sram_raddr_w1[9]) );
  INV_X1 U33 ( .A(1'b1), .ZN(sram_raddr_w0[7]) );
  INV_X1 U35 ( .A(1'b1), .ZN(sram_raddr_w0[8]) );
  INV_X1 U37 ( .A(1'b1), .ZN(sram_raddr_w0[9]) );
  INV_X1 U39 ( .A(n64), .ZN(n25) );
  INV_X1 U40 ( .A(n63), .ZN(n26) );
  INV_X1 U41 ( .A(N9), .ZN(n27) );
  BUF_X1 U42 ( .A(addr_serial_num[1]), .Z(n28) );
  BUF_X1 U43 ( .A(addr_serial_num[0]), .Z(n29) );
  BUF_X1 U44 ( .A(n31), .Z(n30) );
  BUF_X1 U45 ( .A(addr_serial_num[6]), .Z(n31) );
  BUF_X1 U46 ( .A(addr_serial_num[6]), .Z(n32) );
  INV_X1 U47 ( .A(addr_serial_num[5]), .ZN(n33) );
  INV_X1 U48 ( .A(n33), .ZN(n34) );
  INV_X1 U49 ( .A(n33), .ZN(n35) );
  INV_X1 U50 ( .A(n56), .ZN(n36) );
  CLKBUF_X1 U51 ( .A(n58), .Z(n37) );
  CLKBUF_X1 U52 ( .A(n40), .Z(n38) );
  INV_X1 U53 ( .A(n37), .ZN(n39) );
  INV_X1 U54 ( .A(n58), .ZN(n40) );
  INV_X1 U55 ( .A(n64), .ZN(n41) );
  INV_X1 U56 ( .A(n41), .ZN(n42) );
  INV_X1 U57 ( .A(n41), .ZN(n43) );
  INV_X1 U58 ( .A(n63), .ZN(n44) );
  INV_X1 U59 ( .A(n44), .ZN(n45) );
  INV_X1 U60 ( .A(n44), .ZN(n46) );
  INV_X1 U61 ( .A(N9), .ZN(n47) );
  INV_X1 U62 ( .A(n47), .ZN(n48) );
  INV_X1 U63 ( .A(n47), .ZN(n49) );
  INV_X1 U64 ( .A(n66), .ZN(n50) );
  INV_X1 U65 ( .A(n50), .ZN(n51) );
  INV_X1 U66 ( .A(n50), .ZN(n52) );
  INV_X1 U67 ( .A(n37), .ZN(n53) );
  OR2_X1 U68 ( .A1(n68), .A2(n29), .ZN(n54) );
  OR2_X1 U69 ( .A1(n68), .A2(n28), .ZN(n55) );
  INV_X1 U70 ( .A(sub_34_carry[5]), .ZN(n57) );
  XNOR2_X1 U71 ( .A(n35), .B(sub_34_carry[5]), .ZN(N12) );
  XNOR2_X1 U72 ( .A(n30), .B(sub_34_carry[6]), .ZN(N13) );
  NAND2_X1 U73 ( .A1(n56), .A2(n57), .ZN(sub_34_carry[6]) );
  INV_X1 U74 ( .A(addr_serial_num[5]), .ZN(n56) );
  OR2_X1 U75 ( .A1(n26), .A2(n27), .ZN(sub_34_carry[4]) );
  OR2_X1 U76 ( .A1(n25), .A2(sub_34_carry[4]), .ZN(sub_34_carry[5]) );
  XNOR2_X1 U77 ( .A(addr_serial_num[3]), .B(addr_serial_num[2]), .ZN(N10) );
  XNOR2_X1 U78 ( .A(addr_serial_num[4]), .B(sub_34_carry[4]), .ZN(N11) );
  INV_X1 U79 ( .A(addr_serial_num[2]), .ZN(N9) );
  OR2_X1 U80 ( .A1(N13), .A2(n39), .ZN(sram_raddr_w1_nx[6]) );
  OR2_X1 U81 ( .A1(N12), .A2(n38), .ZN(sram_raddr_w1_nx[5]) );
  OR2_X1 U82 ( .A1(N11), .A2(n53), .ZN(sram_raddr_w1_nx[4]) );
  OR2_X1 U83 ( .A1(N10), .A2(n40), .ZN(sram_raddr_w1_nx[3]) );
  OR2_X1 U84 ( .A1(n48), .A2(n38), .ZN(sram_raddr_w1_nx[2]) );
  OR2_X1 U85 ( .A1(n28), .A2(n53), .ZN(sram_raddr_w1_nx[1]) );
  OR2_X1 U86 ( .A1(n29), .A2(n39), .ZN(sram_raddr_w1_nx[0]) );
  MUX2_X1 U87 ( .A(n59), .B(n60), .S(n32), .Z(n58) );
  NAND2_X1 U88 ( .A1(n36), .A2(n61), .ZN(n60) );
  OAI211_X1 U89 ( .C1(n62), .C2(n49), .A(n46), .B(n43), .ZN(n61) );
  OR2_X1 U90 ( .A1(n65), .A2(n34), .ZN(n59) );
  NAND2_X1 U91 ( .A1(n42), .A2(n52), .ZN(sram_raddr_w0_nx_4_) );
  NAND2_X1 U92 ( .A1(n45), .A2(n51), .ZN(sram_raddr_w0_nx_3_) );
  NAND2_X1 U93 ( .A1(n49), .A2(n52), .ZN(sram_raddr_w0_nx_2_) );
  INV_X1 U94 ( .A(n51), .ZN(n68) );
  OAI211_X1 U95 ( .C1(n67), .C2(n65), .A(n31), .B(n35), .ZN(n66) );
  NAND3_X1 U96 ( .A1(n45), .A2(n42), .A3(n48), .ZN(n65) );
  INV_X1 U97 ( .A(addr_serial_num[4]), .ZN(n64) );
  INV_X1 U98 ( .A(addr_serial_num[3]), .ZN(n63) );
  INV_X1 U99 ( .A(n62), .ZN(n67) );
  NAND2_X1 U100 ( .A1(addr_serial_num[1]), .A2(addr_serial_num[0]), .ZN(n62)
         );
endmodule



    module quantize_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_OUTPUT_DATA_WIDTH16 ( 
        ori_data, quantized_data );
  input [167:0] ori_data;
  output [127:0] quantized_data;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432;

  INV_X1 U3 ( .A(n389), .ZN(n1) );
  INV_X1 U4 ( .A(n412), .ZN(n2) );
  INV_X1 U5 ( .A(n266), .ZN(n3) );
  INV_X1 U6 ( .A(n290), .ZN(n4) );
  INV_X1 U7 ( .A(n313), .ZN(n5) );
  INV_X1 U8 ( .A(n337), .ZN(n6) );
  INV_X1 U9 ( .A(n360), .ZN(n7) );
  INV_X1 U10 ( .A(n384), .ZN(n8) );
  CLKBUF_X1 U11 ( .A(n257), .Z(n9) );
  CLKBUF_X1 U12 ( .A(n56), .Z(n10) );
  CLKBUF_X1 U13 ( .A(n361), .Z(n11) );
  CLKBUF_X1 U14 ( .A(n59), .Z(n12) );
  CLKBUF_X1 U15 ( .A(n390), .Z(n13) );
  CLKBUF_X1 U16 ( .A(n62), .Z(n14) );
  CLKBUF_X1 U17 ( .A(n314), .Z(n15) );
  CLKBUF_X1 U18 ( .A(n65), .Z(n16) );
  CLKBUF_X1 U19 ( .A(n338), .Z(n17) );
  CLKBUF_X1 U20 ( .A(n68), .Z(n18) );
  CLKBUF_X1 U21 ( .A(n267), .Z(n19) );
  CLKBUF_X1 U22 ( .A(n71), .Z(n20) );
  CLKBUF_X1 U23 ( .A(n291), .Z(n21) );
  CLKBUF_X1 U24 ( .A(n74), .Z(n22) );
  CLKBUF_X1 U25 ( .A(n317), .Z(n23) );
  CLKBUF_X1 U26 ( .A(n77), .Z(n24) );
  CLKBUF_X1 U27 ( .A(n341), .Z(n25) );
  CLKBUF_X1 U28 ( .A(n80), .Z(n26) );
  CLKBUF_X1 U29 ( .A(n393), .Z(n27) );
  CLKBUF_X1 U30 ( .A(n87), .Z(n28) );
  CLKBUF_X1 U31 ( .A(n294), .Z(n29) );
  CLKBUF_X1 U32 ( .A(n90), .Z(n30) );
  CLKBUF_X1 U33 ( .A(n364), .Z(n31) );
  CLKBUF_X1 U34 ( .A(n93), .Z(n32) );
  CLKBUF_X1 U35 ( .A(n259), .Z(n33) );
  CLKBUF_X1 U36 ( .A(n96), .Z(n34) );
  CLKBUF_X1 U37 ( .A(n270), .Z(n35) );
  CLKBUF_X1 U38 ( .A(n99), .Z(n36) );
  CLKBUF_X1 U39 ( .A(n9), .Z(n37) );
  CLKBUF_X1 U40 ( .A(n11), .Z(n38) );
  CLKBUF_X1 U41 ( .A(n13), .Z(n39) );
  CLKBUF_X1 U42 ( .A(n15), .Z(n40) );
  CLKBUF_X1 U43 ( .A(n17), .Z(n41) );
  CLKBUF_X1 U44 ( .A(n19), .Z(n42) );
  CLKBUF_X1 U45 ( .A(n21), .Z(n43) );
  CLKBUF_X1 U46 ( .A(n23), .Z(n44) );
  CLKBUF_X1 U47 ( .A(n25), .Z(n45) );
  CLKBUF_X1 U48 ( .A(n83), .Z(n46) );
  CLKBUF_X1 U49 ( .A(n27), .Z(n47) );
  CLKBUF_X1 U50 ( .A(n29), .Z(n48) );
  CLKBUF_X1 U51 ( .A(n31), .Z(n49) );
  CLKBUF_X1 U52 ( .A(n33), .Z(n50) );
  CLKBUF_X1 U53 ( .A(n35), .Z(n51) );
  CLKBUF_X1 U54 ( .A(n229), .Z(n52) );
  INV_X1 U55 ( .A(n232), .ZN(n53) );
  INV_X1 U56 ( .A(n53), .ZN(n54) );
  INV_X1 U57 ( .A(n53), .ZN(n55) );
  INV_X1 U58 ( .A(n9), .ZN(n56) );
  INV_X1 U59 ( .A(n10), .ZN(n57) );
  INV_X1 U60 ( .A(n10), .ZN(n58) );
  INV_X1 U61 ( .A(n11), .ZN(n59) );
  INV_X1 U62 ( .A(n12), .ZN(n60) );
  INV_X1 U63 ( .A(n12), .ZN(n61) );
  INV_X1 U64 ( .A(n13), .ZN(n62) );
  INV_X1 U65 ( .A(n14), .ZN(n63) );
  INV_X1 U66 ( .A(n14), .ZN(n64) );
  INV_X1 U67 ( .A(n15), .ZN(n65) );
  INV_X1 U68 ( .A(n16), .ZN(n66) );
  INV_X1 U69 ( .A(n16), .ZN(n67) );
  INV_X1 U70 ( .A(n17), .ZN(n68) );
  INV_X1 U71 ( .A(n18), .ZN(n69) );
  INV_X1 U72 ( .A(n18), .ZN(n70) );
  INV_X1 U73 ( .A(n19), .ZN(n71) );
  INV_X1 U74 ( .A(n20), .ZN(n72) );
  INV_X1 U75 ( .A(n20), .ZN(n73) );
  INV_X1 U76 ( .A(n21), .ZN(n74) );
  INV_X1 U77 ( .A(n22), .ZN(n75) );
  INV_X1 U78 ( .A(n22), .ZN(n76) );
  INV_X1 U79 ( .A(n23), .ZN(n77) );
  INV_X1 U80 ( .A(n24), .ZN(n78) );
  INV_X1 U81 ( .A(n24), .ZN(n79) );
  INV_X1 U82 ( .A(n25), .ZN(n80) );
  INV_X1 U83 ( .A(n26), .ZN(n81) );
  INV_X1 U84 ( .A(n26), .ZN(n82) );
  INV_X1 U85 ( .A(n242), .ZN(n83) );
  INV_X1 U86 ( .A(n83), .ZN(n84) );
  INV_X1 U87 ( .A(n242), .ZN(n85) );
  INV_X1 U88 ( .A(n84), .ZN(n86) );
  INV_X1 U89 ( .A(n27), .ZN(n87) );
  INV_X1 U90 ( .A(n28), .ZN(n88) );
  INV_X1 U91 ( .A(n28), .ZN(n89) );
  INV_X1 U92 ( .A(n29), .ZN(n90) );
  INV_X1 U93 ( .A(n30), .ZN(n91) );
  INV_X1 U94 ( .A(n30), .ZN(n92) );
  INV_X1 U95 ( .A(n31), .ZN(n93) );
  INV_X1 U96 ( .A(n32), .ZN(n94) );
  INV_X1 U97 ( .A(n32), .ZN(n95) );
  INV_X1 U98 ( .A(n33), .ZN(n96) );
  INV_X1 U99 ( .A(n34), .ZN(n97) );
  INV_X1 U100 ( .A(n34), .ZN(n98) );
  INV_X1 U101 ( .A(n35), .ZN(n99) );
  INV_X1 U102 ( .A(n36), .ZN(n100) );
  INV_X1 U103 ( .A(n36), .ZN(n101) );
  CLKBUF_X1 U104 ( .A(n260), .Z(n102) );
  INV_X1 U105 ( .A(n54), .ZN(n103) );
  INV_X1 U106 ( .A(n103), .ZN(n104) );
  INV_X1 U107 ( .A(n103), .ZN(n105) );
  INV_X1 U108 ( .A(n232), .ZN(n106) );
  INV_X1 U109 ( .A(n106), .ZN(n107) );
  INV_X1 U110 ( .A(n106), .ZN(n108) );
  CLKBUF_X1 U111 ( .A(n110), .Z(n109) );
  CLKBUF_X1 U112 ( .A(n257), .Z(n110) );
  INV_X1 U113 ( .A(n110), .ZN(n111) );
  INV_X1 U114 ( .A(n111), .ZN(n112) );
  INV_X1 U115 ( .A(n111), .ZN(n113) );
  INV_X1 U116 ( .A(n57), .ZN(n114) );
  INV_X1 U117 ( .A(n114), .ZN(n115) );
  INV_X1 U118 ( .A(n114), .ZN(n116) );
  CLKBUF_X1 U119 ( .A(n118), .Z(n117) );
  CLKBUF_X1 U120 ( .A(n361), .Z(n118) );
  INV_X1 U121 ( .A(n60), .ZN(n119) );
  INV_X1 U122 ( .A(n119), .ZN(n120) );
  INV_X1 U123 ( .A(n119), .ZN(n121) );
  INV_X1 U124 ( .A(n118), .ZN(n122) );
  INV_X1 U125 ( .A(n122), .ZN(n123) );
  INV_X1 U126 ( .A(n122), .ZN(n124) );
  CLKBUF_X1 U127 ( .A(n126), .Z(n125) );
  CLKBUF_X1 U128 ( .A(n390), .Z(n126) );
  INV_X1 U129 ( .A(n63), .ZN(n127) );
  INV_X1 U130 ( .A(n127), .ZN(n128) );
  INV_X1 U131 ( .A(n127), .ZN(n129) );
  INV_X1 U132 ( .A(n126), .ZN(n130) );
  INV_X1 U133 ( .A(n130), .ZN(n131) );
  INV_X1 U134 ( .A(n130), .ZN(n132) );
  CLKBUF_X1 U135 ( .A(n134), .Z(n133) );
  CLKBUF_X1 U136 ( .A(n314), .Z(n134) );
  INV_X1 U137 ( .A(n66), .ZN(n135) );
  INV_X1 U138 ( .A(n135), .ZN(n136) );
  INV_X1 U139 ( .A(n135), .ZN(n137) );
  INV_X1 U140 ( .A(n134), .ZN(n138) );
  INV_X1 U141 ( .A(n138), .ZN(n139) );
  INV_X1 U142 ( .A(n138), .ZN(n140) );
  CLKBUF_X1 U143 ( .A(n142), .Z(n141) );
  CLKBUF_X1 U144 ( .A(n338), .Z(n142) );
  INV_X1 U145 ( .A(n69), .ZN(n143) );
  INV_X1 U146 ( .A(n143), .ZN(n144) );
  INV_X1 U147 ( .A(n143), .ZN(n145) );
  INV_X1 U148 ( .A(n142), .ZN(n146) );
  INV_X1 U149 ( .A(n146), .ZN(n147) );
  INV_X1 U150 ( .A(n146), .ZN(n148) );
  CLKBUF_X1 U151 ( .A(n150), .Z(n149) );
  CLKBUF_X1 U152 ( .A(n267), .Z(n150) );
  INV_X1 U153 ( .A(n150), .ZN(n151) );
  INV_X1 U154 ( .A(n151), .ZN(n152) );
  INV_X1 U155 ( .A(n151), .ZN(n153) );
  INV_X1 U156 ( .A(n72), .ZN(n154) );
  INV_X1 U157 ( .A(n154), .ZN(n155) );
  INV_X1 U158 ( .A(n154), .ZN(n156) );
  CLKBUF_X1 U159 ( .A(n158), .Z(n157) );
  CLKBUF_X1 U160 ( .A(n291), .Z(n158) );
  INV_X1 U161 ( .A(n75), .ZN(n159) );
  INV_X1 U162 ( .A(n159), .ZN(n160) );
  INV_X1 U163 ( .A(n159), .ZN(n161) );
  INV_X1 U164 ( .A(n158), .ZN(n162) );
  INV_X1 U165 ( .A(n162), .ZN(n163) );
  INV_X1 U166 ( .A(n162), .ZN(n164) );
  CLKBUF_X1 U167 ( .A(n166), .Z(n165) );
  CLKBUF_X1 U168 ( .A(n317), .Z(n166) );
  INV_X1 U169 ( .A(n44), .ZN(n167) );
  INV_X1 U170 ( .A(n167), .ZN(n168) );
  INV_X1 U171 ( .A(n167), .ZN(n169) );
  INV_X1 U172 ( .A(n166), .ZN(n170) );
  INV_X1 U173 ( .A(n170), .ZN(n171) );
  INV_X1 U174 ( .A(n170), .ZN(n172) );
  CLKBUF_X1 U175 ( .A(n174), .Z(n173) );
  CLKBUF_X1 U176 ( .A(n341), .Z(n174) );
  INV_X1 U177 ( .A(n45), .ZN(n175) );
  INV_X1 U178 ( .A(n175), .ZN(n176) );
  INV_X1 U179 ( .A(n175), .ZN(n177) );
  INV_X1 U180 ( .A(n174), .ZN(n178) );
  INV_X1 U181 ( .A(n178), .ZN(n179) );
  INV_X1 U182 ( .A(n178), .ZN(n180) );
  CLKBUF_X1 U183 ( .A(n182), .Z(n181) );
  CLKBUF_X1 U184 ( .A(n262), .Z(n182) );
  INV_X1 U185 ( .A(n182), .ZN(n183) );
  INV_X1 U186 ( .A(n183), .ZN(n184) );
  INV_X1 U187 ( .A(n183), .ZN(n185) );
  INV_X1 U188 ( .A(n46), .ZN(n186) );
  INV_X1 U189 ( .A(n186), .ZN(n187) );
  INV_X1 U190 ( .A(n186), .ZN(n188) );
  CLKBUF_X1 U191 ( .A(n190), .Z(n189) );
  CLKBUF_X1 U192 ( .A(n393), .Z(n190) );
  INV_X1 U193 ( .A(n47), .ZN(n191) );
  INV_X1 U194 ( .A(n191), .ZN(n192) );
  INV_X1 U195 ( .A(n191), .ZN(n193) );
  INV_X1 U196 ( .A(n190), .ZN(n194) );
  INV_X1 U197 ( .A(n194), .ZN(n195) );
  INV_X1 U198 ( .A(n194), .ZN(n196) );
  CLKBUF_X1 U199 ( .A(n198), .Z(n197) );
  CLKBUF_X1 U200 ( .A(n294), .Z(n198) );
  INV_X1 U201 ( .A(n48), .ZN(n199) );
  INV_X1 U202 ( .A(n199), .ZN(n200) );
  INV_X1 U203 ( .A(n199), .ZN(n201) );
  INV_X1 U204 ( .A(n198), .ZN(n202) );
  INV_X1 U205 ( .A(n202), .ZN(n203) );
  INV_X1 U206 ( .A(n202), .ZN(n204) );
  CLKBUF_X1 U207 ( .A(n206), .Z(n205) );
  CLKBUF_X1 U208 ( .A(n364), .Z(n206) );
  INV_X1 U209 ( .A(n49), .ZN(n207) );
  INV_X1 U210 ( .A(n207), .ZN(n208) );
  INV_X1 U211 ( .A(n207), .ZN(n209) );
  INV_X1 U212 ( .A(n206), .ZN(n210) );
  INV_X1 U213 ( .A(n210), .ZN(n211) );
  INV_X1 U214 ( .A(n210), .ZN(n212) );
  CLKBUF_X1 U215 ( .A(n214), .Z(n213) );
  CLKBUF_X1 U216 ( .A(n259), .Z(n214) );
  INV_X1 U217 ( .A(n214), .ZN(n215) );
  INV_X1 U218 ( .A(n215), .ZN(n216) );
  INV_X1 U219 ( .A(n215), .ZN(n217) );
  INV_X1 U220 ( .A(n50), .ZN(n218) );
  INV_X1 U221 ( .A(n218), .ZN(n219) );
  INV_X1 U222 ( .A(n218), .ZN(n220) );
  CLKBUF_X1 U223 ( .A(n222), .Z(n221) );
  CLKBUF_X1 U224 ( .A(n270), .Z(n222) );
  INV_X1 U225 ( .A(n222), .ZN(n223) );
  INV_X1 U226 ( .A(n223), .ZN(n224) );
  INV_X1 U227 ( .A(n223), .ZN(n225) );
  INV_X1 U228 ( .A(n51), .ZN(n226) );
  INV_X1 U229 ( .A(n226), .ZN(n227) );
  INV_X1 U230 ( .A(n226), .ZN(n228) );
  INV_X1 U231 ( .A(n260), .ZN(n229) );
  INV_X1 U232 ( .A(n52), .ZN(n230) );
  INV_X1 U233 ( .A(n52), .ZN(n231) );
  INV_X1 U234 ( .A(n229), .ZN(n232) );
  INV_X1 U235 ( .A(n56), .ZN(n233) );
  INV_X1 U236 ( .A(n59), .ZN(n234) );
  INV_X1 U237 ( .A(n62), .ZN(n235) );
  INV_X1 U238 ( .A(n65), .ZN(n236) );
  INV_X1 U239 ( .A(n68), .ZN(n237) );
  INV_X1 U240 ( .A(n71), .ZN(n238) );
  INV_X1 U241 ( .A(n74), .ZN(n239) );
  INV_X1 U242 ( .A(n77), .ZN(n240) );
  INV_X1 U243 ( .A(n80), .ZN(n241) );
  INV_X1 U244 ( .A(n262), .ZN(n242) );
  INV_X1 U245 ( .A(n84), .ZN(n243) );
  INV_X1 U246 ( .A(n87), .ZN(n244) );
  INV_X1 U247 ( .A(n90), .ZN(n245) );
  INV_X1 U248 ( .A(n93), .ZN(n246) );
  INV_X1 U249 ( .A(n96), .ZN(n247) );
  INV_X1 U250 ( .A(n99), .ZN(n248) );
  OR2_X1 U251 ( .A1(n249), .A2(ori_data[20]), .ZN(n259) );
  NOR4_X1 U252 ( .A1(n8), .A2(ori_data[16]), .A3(n430), .A4(ori_data[17]), 
        .ZN(n249) );
  OR2_X1 U253 ( .A1(n250), .A2(ori_data[125]), .ZN(n270) );
  NOR4_X1 U254 ( .A1(n3), .A2(ori_data[121]), .A3(n286), .A4(ori_data[122]), 
        .ZN(n250) );
  OR2_X1 U255 ( .A1(n251), .A2(ori_data[104]), .ZN(n294) );
  NOR4_X1 U256 ( .A1(ori_data[100]), .A2(ori_data[101]), .A3(n310), .A4(
        ori_data[102]), .ZN(n251) );
  OR2_X1 U257 ( .A1(n252), .A2(ori_data[41]), .ZN(n364) );
  NOR4_X1 U258 ( .A1(n7), .A2(ori_data[37]), .A3(n381), .A4(ori_data[38]), 
        .ZN(n252) );
  OR2_X1 U259 ( .A1(n253), .A2(ori_data[146]), .ZN(n262) );
  NOR4_X1 U260 ( .A1(n2), .A2(ori_data[142]), .A3(n426), .A4(ori_data[143]), 
        .ZN(n253) );
  OR2_X1 U261 ( .A1(n254), .A2(ori_data[167]), .ZN(n393) );
  NOR4_X1 U262 ( .A1(n1), .A2(ori_data[163]), .A3(n409), .A4(ori_data[164]), 
        .ZN(n254) );
  OR2_X1 U263 ( .A1(n255), .A2(ori_data[83]), .ZN(n317) );
  NOR4_X1 U264 ( .A1(n5), .A2(ori_data[79]), .A3(n334), .A4(ori_data[80]), 
        .ZN(n255) );
  OR2_X1 U265 ( .A1(n256), .A2(ori_data[62]), .ZN(n341) );
  NOR4_X1 U266 ( .A1(n6), .A2(ori_data[58]), .A3(n357), .A4(ori_data[59]), 
        .ZN(n256) );
  OAI21_X1 U267 ( .B1(n115), .B2(n258), .A(n219), .ZN(quantized_data[9]) );
  INV_X1 U268 ( .A(ori_data[9]), .ZN(n258) );
  OAI21_X1 U269 ( .B1(n55), .B2(n261), .A(n188), .ZN(quantized_data[99]) );
  INV_X1 U270 ( .A(ori_data[129]), .ZN(n261) );
  OAI21_X1 U271 ( .B1(n54), .B2(n263), .A(n46), .ZN(quantized_data[98]) );
  INV_X1 U272 ( .A(ori_data[128]), .ZN(n263) );
  OAI21_X1 U273 ( .B1(n102), .B2(n264), .A(n185), .ZN(quantized_data[97]) );
  INV_X1 U274 ( .A(ori_data[127]), .ZN(n264) );
  OAI21_X1 U275 ( .B1(n107), .B2(n265), .A(n86), .ZN(quantized_data[96]) );
  INV_X1 U276 ( .A(ori_data[126]), .ZN(n265) );
  OAI21_X1 U277 ( .B1(n266), .B2(n42), .A(n268), .ZN(quantized_data[95]) );
  INV_X1 U278 ( .A(ori_data[120]), .ZN(n266) );
  OAI21_X1 U279 ( .B1(n238), .B2(n269), .A(n221), .ZN(quantized_data[94]) );
  INV_X1 U280 ( .A(ori_data[119]), .ZN(n269) );
  OAI21_X1 U281 ( .B1(n149), .B2(n271), .A(n248), .ZN(quantized_data[93]) );
  INV_X1 U282 ( .A(ori_data[118]), .ZN(n271) );
  OAI21_X1 U283 ( .B1(n155), .B2(n272), .A(n227), .ZN(quantized_data[92]) );
  INV_X1 U284 ( .A(ori_data[117]), .ZN(n272) );
  OAI21_X1 U285 ( .B1(n156), .B2(n273), .A(n228), .ZN(quantized_data[91]) );
  INV_X1 U286 ( .A(ori_data[116]), .ZN(n273) );
  OAI21_X1 U287 ( .B1(n152), .B2(n274), .A(n225), .ZN(quantized_data[90]) );
  INV_X1 U288 ( .A(ori_data[115]), .ZN(n274) );
  OAI21_X1 U289 ( .B1(n113), .B2(n275), .A(n217), .ZN(quantized_data[8]) );
  INV_X1 U290 ( .A(ori_data[8]), .ZN(n275) );
  OAI21_X1 U291 ( .B1(n155), .B2(n276), .A(n228), .ZN(quantized_data[89]) );
  INV_X1 U292 ( .A(ori_data[114]), .ZN(n276) );
  OAI21_X1 U293 ( .B1(n152), .B2(n277), .A(n224), .ZN(quantized_data[88]) );
  INV_X1 U294 ( .A(ori_data[113]), .ZN(n277) );
  OAI21_X1 U295 ( .B1(n153), .B2(n278), .A(n224), .ZN(quantized_data[87]) );
  INV_X1 U296 ( .A(ori_data[112]), .ZN(n278) );
  OAI21_X1 U297 ( .B1(n238), .B2(n279), .A(n51), .ZN(quantized_data[86]) );
  INV_X1 U298 ( .A(ori_data[111]), .ZN(n279) );
  OAI21_X1 U299 ( .B1(n149), .B2(n280), .A(n101), .ZN(quantized_data[85]) );
  INV_X1 U300 ( .A(ori_data[110]), .ZN(n280) );
  OAI21_X1 U301 ( .B1(n42), .B2(n281), .A(n248), .ZN(quantized_data[84]) );
  INV_X1 U302 ( .A(ori_data[109]), .ZN(n281) );
  OAI21_X1 U303 ( .B1(n73), .B2(n282), .A(n100), .ZN(quantized_data[83]) );
  INV_X1 U304 ( .A(ori_data[108]), .ZN(n282) );
  OAI21_X1 U305 ( .B1(n156), .B2(n283), .A(n227), .ZN(quantized_data[82]) );
  INV_X1 U306 ( .A(ori_data[107]), .ZN(n283) );
  OAI21_X1 U307 ( .B1(n153), .B2(n284), .A(n225), .ZN(quantized_data[81]) );
  INV_X1 U308 ( .A(ori_data[106]), .ZN(n284) );
  OAI21_X1 U309 ( .B1(n72), .B2(n285), .A(n221), .ZN(quantized_data[80]) );
  INV_X1 U310 ( .A(ori_data[105]), .ZN(n285) );
  NAND2_X1 U311 ( .A1(n268), .A2(n100), .ZN(n267) );
  OR2_X1 U312 ( .A1(ori_data[124]), .A2(ori_data[123]), .ZN(n286) );
  OAI21_X1 U313 ( .B1(n287), .B2(n288), .A(ori_data[125]), .ZN(n268) );
  NAND2_X1 U314 ( .A1(ori_data[124]), .A2(ori_data[123]), .ZN(n288) );
  NAND3_X1 U315 ( .A1(ori_data[121]), .A2(ori_data[120]), .A3(ori_data[122]), 
        .ZN(n287) );
  OAI21_X1 U316 ( .B1(n58), .B2(n289), .A(n213), .ZN(quantized_data[7]) );
  INV_X1 U317 ( .A(ori_data[7]), .ZN(n289) );
  OAI21_X1 U318 ( .B1(n290), .B2(n43), .A(n292), .ZN(quantized_data[79]) );
  INV_X1 U319 ( .A(ori_data[99]), .ZN(n290) );
  OAI21_X1 U320 ( .B1(n163), .B2(n293), .A(n203), .ZN(quantized_data[78]) );
  INV_X1 U321 ( .A(ori_data[98]), .ZN(n293) );
  OAI21_X1 U322 ( .B1(n157), .B2(n295), .A(n91), .ZN(quantized_data[77]) );
  INV_X1 U323 ( .A(ori_data[97]), .ZN(n295) );
  OAI21_X1 U324 ( .B1(n164), .B2(n296), .A(n204), .ZN(quantized_data[76]) );
  INV_X1 U325 ( .A(ori_data[96]), .ZN(n296) );
  OAI21_X1 U326 ( .B1(n161), .B2(n297), .A(n201), .ZN(quantized_data[75]) );
  INV_X1 U327 ( .A(ori_data[95]), .ZN(n297) );
  OAI21_X1 U328 ( .B1(n43), .B2(n298), .A(n92), .ZN(quantized_data[74]) );
  INV_X1 U329 ( .A(ori_data[94]), .ZN(n298) );
  OAI21_X1 U330 ( .B1(n161), .B2(n299), .A(n201), .ZN(quantized_data[73]) );
  INV_X1 U331 ( .A(ori_data[93]), .ZN(n299) );
  OAI21_X1 U332 ( .B1(n239), .B2(n300), .A(n48), .ZN(quantized_data[72]) );
  INV_X1 U333 ( .A(ori_data[92]), .ZN(n300) );
  OAI21_X1 U334 ( .B1(n75), .B2(n301), .A(n197), .ZN(quantized_data[71]) );
  INV_X1 U335 ( .A(ori_data[91]), .ZN(n301) );
  OAI21_X1 U336 ( .B1(n163), .B2(n302), .A(n203), .ZN(quantized_data[70]) );
  INV_X1 U337 ( .A(ori_data[90]), .ZN(n302) );
  OAI21_X1 U338 ( .B1(n37), .B2(n303), .A(n213), .ZN(quantized_data[6]) );
  INV_X1 U339 ( .A(ori_data[6]), .ZN(n303) );
  OAI21_X1 U340 ( .B1(n239), .B2(n304), .A(n245), .ZN(quantized_data[69]) );
  INV_X1 U341 ( .A(ori_data[89]), .ZN(n304) );
  OAI21_X1 U342 ( .B1(n164), .B2(n305), .A(n204), .ZN(quantized_data[68]) );
  INV_X1 U343 ( .A(ori_data[88]), .ZN(n305) );
  OAI21_X1 U344 ( .B1(n160), .B2(n306), .A(n200), .ZN(quantized_data[67]) );
  INV_X1 U345 ( .A(ori_data[87]), .ZN(n306) );
  OAI21_X1 U346 ( .B1(n76), .B2(n307), .A(n245), .ZN(quantized_data[66]) );
  INV_X1 U347 ( .A(ori_data[86]), .ZN(n307) );
  OAI21_X1 U348 ( .B1(n160), .B2(n308), .A(n200), .ZN(quantized_data[65]) );
  INV_X1 U349 ( .A(ori_data[85]), .ZN(n308) );
  OAI21_X1 U350 ( .B1(n157), .B2(n309), .A(n197), .ZN(quantized_data[64]) );
  INV_X1 U351 ( .A(ori_data[84]), .ZN(n309) );
  NAND2_X1 U352 ( .A1(n292), .A2(n91), .ZN(n291) );
  OR2_X1 U353 ( .A1(n4), .A2(ori_data[103]), .ZN(n310) );
  OAI21_X1 U354 ( .B1(n311), .B2(n312), .A(ori_data[104]), .ZN(n292) );
  NAND2_X1 U355 ( .A1(ori_data[99]), .A2(ori_data[103]), .ZN(n312) );
  NAND3_X1 U356 ( .A1(ori_data[101]), .A2(ori_data[100]), .A3(ori_data[102]), 
        .ZN(n311) );
  OAI21_X1 U357 ( .B1(n313), .B2(n40), .A(n315), .ZN(quantized_data[63]) );
  INV_X1 U358 ( .A(ori_data[78]), .ZN(n313) );
  OAI21_X1 U359 ( .B1(n137), .B2(n316), .A(n165), .ZN(quantized_data[62]) );
  INV_X1 U360 ( .A(ori_data[77]), .ZN(n316) );
  OAI21_X1 U361 ( .B1(n137), .B2(n318), .A(n171), .ZN(quantized_data[61]) );
  INV_X1 U362 ( .A(ori_data[76]), .ZN(n318) );
  OAI21_X1 U363 ( .B1(n236), .B2(n319), .A(n172), .ZN(quantized_data[60]) );
  INV_X1 U364 ( .A(ori_data[75]), .ZN(n319) );
  OAI21_X1 U365 ( .B1(n116), .B2(n320), .A(n220), .ZN(quantized_data[5]) );
  INV_X1 U366 ( .A(ori_data[5]), .ZN(n320) );
  OAI21_X1 U367 ( .B1(n139), .B2(n321), .A(n169), .ZN(quantized_data[59]) );
  INV_X1 U368 ( .A(ori_data[74]), .ZN(n321) );
  OAI21_X1 U369 ( .B1(n136), .B2(n322), .A(n168), .ZN(quantized_data[58]) );
  INV_X1 U370 ( .A(ori_data[73]), .ZN(n322) );
  OAI21_X1 U371 ( .B1(n67), .B2(n323), .A(n165), .ZN(quantized_data[57]) );
  INV_X1 U372 ( .A(ori_data[72]), .ZN(n323) );
  OAI21_X1 U373 ( .B1(n139), .B2(n324), .A(n79), .ZN(quantized_data[56]) );
  INV_X1 U374 ( .A(ori_data[71]), .ZN(n324) );
  OAI21_X1 U375 ( .B1(n40), .B2(n325), .A(n78), .ZN(quantized_data[55]) );
  INV_X1 U376 ( .A(ori_data[70]), .ZN(n325) );
  OAI21_X1 U377 ( .B1(n133), .B2(n326), .A(n171), .ZN(quantized_data[54]) );
  INV_X1 U378 ( .A(ori_data[69]), .ZN(n326) );
  OAI21_X1 U379 ( .B1(n140), .B2(n327), .A(n169), .ZN(quantized_data[53]) );
  INV_X1 U380 ( .A(ori_data[68]), .ZN(n327) );
  OAI21_X1 U381 ( .B1(n136), .B2(n328), .A(n44), .ZN(quantized_data[52]) );
  INV_X1 U382 ( .A(ori_data[67]), .ZN(n328) );
  OAI21_X1 U383 ( .B1(n236), .B2(n329), .A(n240), .ZN(quantized_data[51]) );
  INV_X1 U384 ( .A(ori_data[66]), .ZN(n329) );
  OAI21_X1 U385 ( .B1(n66), .B2(n330), .A(n172), .ZN(quantized_data[50]) );
  INV_X1 U386 ( .A(ori_data[65]), .ZN(n330) );
  OAI21_X1 U387 ( .B1(n109), .B2(n331), .A(n97), .ZN(quantized_data[4]) );
  INV_X1 U388 ( .A(ori_data[4]), .ZN(n331) );
  OAI21_X1 U389 ( .B1(n133), .B2(n332), .A(n168), .ZN(quantized_data[49]) );
  INV_X1 U390 ( .A(ori_data[64]), .ZN(n332) );
  OAI21_X1 U391 ( .B1(n140), .B2(n333), .A(n240), .ZN(quantized_data[48]) );
  INV_X1 U392 ( .A(ori_data[63]), .ZN(n333) );
  NAND2_X1 U393 ( .A1(n315), .A2(n78), .ZN(n314) );
  OR2_X1 U394 ( .A1(ori_data[82]), .A2(ori_data[81]), .ZN(n334) );
  OAI21_X1 U395 ( .B1(n335), .B2(n336), .A(ori_data[83]), .ZN(n315) );
  NAND2_X1 U396 ( .A1(ori_data[82]), .A2(ori_data[81]), .ZN(n336) );
  NAND3_X1 U397 ( .A1(ori_data[79]), .A2(ori_data[78]), .A3(ori_data[80]), 
        .ZN(n335) );
  OAI21_X1 U398 ( .B1(n337), .B2(n41), .A(n339), .ZN(quantized_data[47]) );
  INV_X1 U399 ( .A(ori_data[57]), .ZN(n337) );
  OAI21_X1 U400 ( .B1(n70), .B2(n340), .A(n241), .ZN(quantized_data[46]) );
  INV_X1 U401 ( .A(ori_data[56]), .ZN(n340) );
  OAI21_X1 U402 ( .B1(n141), .B2(n342), .A(n180), .ZN(quantized_data[45]) );
  INV_X1 U403 ( .A(ori_data[55]), .ZN(n342) );
  OAI21_X1 U404 ( .B1(n237), .B2(n343), .A(n179), .ZN(quantized_data[44]) );
  INV_X1 U405 ( .A(ori_data[54]), .ZN(n343) );
  OAI21_X1 U406 ( .B1(n148), .B2(n344), .A(n177), .ZN(quantized_data[43]) );
  INV_X1 U407 ( .A(ori_data[53]), .ZN(n344) );
  OAI21_X1 U408 ( .B1(n141), .B2(n345), .A(n176), .ZN(quantized_data[42]) );
  INV_X1 U409 ( .A(ori_data[52]), .ZN(n345) );
  OAI21_X1 U410 ( .B1(n144), .B2(n346), .A(n81), .ZN(quantized_data[41]) );
  INV_X1 U411 ( .A(ori_data[51]), .ZN(n346) );
  OAI21_X1 U412 ( .B1(n237), .B2(n347), .A(n82), .ZN(quantized_data[40]) );
  INV_X1 U413 ( .A(ori_data[50]), .ZN(n347) );
  OAI21_X1 U414 ( .B1(n112), .B2(n348), .A(n216), .ZN(quantized_data[3]) );
  INV_X1 U415 ( .A(ori_data[3]), .ZN(n348) );
  OAI21_X1 U416 ( .B1(n145), .B2(n349), .A(n45), .ZN(quantized_data[39]) );
  INV_X1 U417 ( .A(ori_data[49]), .ZN(n349) );
  OAI21_X1 U418 ( .B1(n148), .B2(n350), .A(n180), .ZN(quantized_data[38]) );
  INV_X1 U419 ( .A(ori_data[48]), .ZN(n350) );
  OAI21_X1 U420 ( .B1(n145), .B2(n351), .A(n176), .ZN(quantized_data[37]) );
  INV_X1 U421 ( .A(ori_data[47]), .ZN(n351) );
  OAI21_X1 U422 ( .B1(n41), .B2(n352), .A(n173), .ZN(quantized_data[36]) );
  INV_X1 U423 ( .A(ori_data[46]), .ZN(n352) );
  OAI21_X1 U424 ( .B1(n147), .B2(n353), .A(n173), .ZN(quantized_data[35]) );
  INV_X1 U425 ( .A(ori_data[45]), .ZN(n353) );
  OAI21_X1 U426 ( .B1(n69), .B2(n354), .A(n179), .ZN(quantized_data[34]) );
  INV_X1 U427 ( .A(ori_data[44]), .ZN(n354) );
  OAI21_X1 U428 ( .B1(n144), .B2(n355), .A(n177), .ZN(quantized_data[33]) );
  INV_X1 U429 ( .A(ori_data[43]), .ZN(n355) );
  OAI21_X1 U430 ( .B1(n147), .B2(n356), .A(n241), .ZN(quantized_data[32]) );
  INV_X1 U431 ( .A(ori_data[42]), .ZN(n356) );
  NAND2_X1 U432 ( .A1(n339), .A2(n81), .ZN(n338) );
  OR2_X1 U433 ( .A1(ori_data[61]), .A2(ori_data[60]), .ZN(n357) );
  OAI21_X1 U434 ( .B1(n358), .B2(n359), .A(ori_data[62]), .ZN(n339) );
  NAND2_X1 U435 ( .A1(ori_data[61]), .A2(ori_data[60]), .ZN(n359) );
  NAND3_X1 U436 ( .A1(ori_data[58]), .A2(ori_data[57]), .A3(ori_data[59]), 
        .ZN(n358) );
  OAI21_X1 U437 ( .B1(n360), .B2(n38), .A(n362), .ZN(quantized_data[31]) );
  INV_X1 U438 ( .A(ori_data[36]), .ZN(n360) );
  OAI21_X1 U439 ( .B1(n117), .B2(n363), .A(n211), .ZN(quantized_data[30]) );
  INV_X1 U440 ( .A(ori_data[35]), .ZN(n363) );
  OAI21_X1 U441 ( .B1(n233), .B2(n365), .A(n50), .ZN(quantized_data[2]) );
  INV_X1 U442 ( .A(ori_data[2]), .ZN(n365) );
  OAI21_X1 U443 ( .B1(n117), .B2(n366), .A(n208), .ZN(quantized_data[29]) );
  INV_X1 U444 ( .A(ori_data[34]), .ZN(n366) );
  OAI21_X1 U445 ( .B1(n234), .B2(n367), .A(n49), .ZN(quantized_data[28]) );
  INV_X1 U446 ( .A(ori_data[33]), .ZN(n367) );
  OAI21_X1 U447 ( .B1(n124), .B2(n368), .A(n205), .ZN(quantized_data[27]) );
  INV_X1 U448 ( .A(ori_data[32]), .ZN(n368) );
  OAI21_X1 U449 ( .B1(n120), .B2(n369), .A(n212), .ZN(quantized_data[26]) );
  INV_X1 U450 ( .A(ori_data[31]), .ZN(n369) );
  OAI21_X1 U451 ( .B1(n120), .B2(n370), .A(n94), .ZN(quantized_data[25]) );
  INV_X1 U452 ( .A(ori_data[30]), .ZN(n370) );
  OAI21_X1 U453 ( .B1(n234), .B2(n371), .A(n209), .ZN(quantized_data[24]) );
  INV_X1 U454 ( .A(ori_data[29]), .ZN(n371) );
  OAI21_X1 U455 ( .B1(n121), .B2(n372), .A(n95), .ZN(quantized_data[23]) );
  INV_X1 U456 ( .A(ori_data[28]), .ZN(n372) );
  OAI21_X1 U457 ( .B1(n61), .B2(n373), .A(n205), .ZN(quantized_data[22]) );
  INV_X1 U458 ( .A(ori_data[27]), .ZN(n373) );
  OAI21_X1 U459 ( .B1(n121), .B2(n374), .A(n246), .ZN(quantized_data[21]) );
  INV_X1 U460 ( .A(ori_data[26]), .ZN(n374) );
  OAI21_X1 U461 ( .B1(n38), .B2(n375), .A(n208), .ZN(quantized_data[20]) );
  INV_X1 U462 ( .A(ori_data[25]), .ZN(n375) );
  OAI21_X1 U463 ( .B1(n233), .B2(n376), .A(n247), .ZN(quantized_data[1]) );
  INV_X1 U464 ( .A(ori_data[1]), .ZN(n376) );
  OAI21_X1 U465 ( .B1(n124), .B2(n377), .A(n246), .ZN(quantized_data[19]) );
  INV_X1 U466 ( .A(ori_data[24]), .ZN(n377) );
  OAI21_X1 U467 ( .B1(n60), .B2(n378), .A(n212), .ZN(quantized_data[18]) );
  INV_X1 U468 ( .A(ori_data[23]), .ZN(n378) );
  OAI21_X1 U469 ( .B1(n123), .B2(n379), .A(n211), .ZN(quantized_data[17]) );
  INV_X1 U470 ( .A(ori_data[22]), .ZN(n379) );
  OAI21_X1 U471 ( .B1(n123), .B2(n380), .A(n209), .ZN(quantized_data[16]) );
  INV_X1 U472 ( .A(ori_data[21]), .ZN(n380) );
  NAND2_X1 U473 ( .A1(n362), .A2(n94), .ZN(n361) );
  OR2_X1 U474 ( .A1(ori_data[40]), .A2(ori_data[39]), .ZN(n381) );
  OAI21_X1 U475 ( .B1(n382), .B2(n383), .A(ori_data[41]), .ZN(n362) );
  NAND2_X1 U476 ( .A1(ori_data[40]), .A2(ori_data[39]), .ZN(n383) );
  NAND3_X1 U477 ( .A1(ori_data[37]), .A2(ori_data[36]), .A3(ori_data[38]), 
        .ZN(n382) );
  OAI21_X1 U478 ( .B1(n384), .B2(n37), .A(n385), .ZN(quantized_data[15]) );
  INV_X1 U479 ( .A(ori_data[15]), .ZN(n384) );
  OAI21_X1 U480 ( .B1(n116), .B2(n386), .A(n220), .ZN(quantized_data[14]) );
  INV_X1 U481 ( .A(ori_data[14]), .ZN(n386) );
  OAI21_X1 U482 ( .B1(n115), .B2(n387), .A(n219), .ZN(quantized_data[13]) );
  INV_X1 U483 ( .A(ori_data[13]), .ZN(n387) );
  OAI21_X1 U484 ( .B1(n112), .B2(n388), .A(n216), .ZN(quantized_data[12]) );
  INV_X1 U485 ( .A(ori_data[12]), .ZN(n388) );
  OAI21_X1 U486 ( .B1(n389), .B2(n235), .A(n391), .ZN(quantized_data[127]) );
  INV_X1 U487 ( .A(ori_data[162]), .ZN(n389) );
  OAI21_X1 U488 ( .B1(n132), .B2(n392), .A(n195), .ZN(quantized_data[126]) );
  INV_X1 U489 ( .A(ori_data[161]), .ZN(n392) );
  OAI21_X1 U490 ( .B1(n129), .B2(n394), .A(n192), .ZN(quantized_data[125]) );
  INV_X1 U491 ( .A(ori_data[160]), .ZN(n394) );
  OAI21_X1 U492 ( .B1(n39), .B2(n395), .A(n88), .ZN(quantized_data[124]) );
  INV_X1 U493 ( .A(ori_data[159]), .ZN(n395) );
  OAI21_X1 U494 ( .B1(n125), .B2(n396), .A(n189), .ZN(quantized_data[123]) );
  INV_X1 U495 ( .A(ori_data[158]), .ZN(n396) );
  OAI21_X1 U496 ( .B1(n131), .B2(n397), .A(n196), .ZN(quantized_data[122]) );
  INV_X1 U497 ( .A(ori_data[157]), .ZN(n397) );
  OAI21_X1 U498 ( .B1(n63), .B2(n398), .A(n244), .ZN(quantized_data[121]) );
  INV_X1 U499 ( .A(ori_data[156]), .ZN(n398) );
  OAI21_X1 U500 ( .B1(n128), .B2(n399), .A(n193), .ZN(quantized_data[120]) );
  INV_X1 U501 ( .A(ori_data[155]), .ZN(n399) );
  OAI21_X1 U502 ( .B1(n113), .B2(n400), .A(n217), .ZN(quantized_data[11]) );
  INV_X1 U503 ( .A(ori_data[11]), .ZN(n400) );
  OAI21_X1 U504 ( .B1(n235), .B2(n401), .A(n47), .ZN(quantized_data[119]) );
  INV_X1 U505 ( .A(ori_data[154]), .ZN(n401) );
  OAI21_X1 U506 ( .B1(n39), .B2(n402), .A(n189), .ZN(quantized_data[118]) );
  INV_X1 U507 ( .A(ori_data[153]), .ZN(n402) );
  OAI21_X1 U508 ( .B1(n125), .B2(n403), .A(n89), .ZN(quantized_data[117]) );
  INV_X1 U509 ( .A(ori_data[152]), .ZN(n403) );
  OAI21_X1 U510 ( .B1(n128), .B2(n404), .A(n192), .ZN(quantized_data[116]) );
  INV_X1 U511 ( .A(ori_data[151]), .ZN(n404) );
  OAI21_X1 U512 ( .B1(n64), .B2(n405), .A(n244), .ZN(quantized_data[115]) );
  INV_X1 U513 ( .A(ori_data[150]), .ZN(n405) );
  OAI21_X1 U514 ( .B1(n132), .B2(n406), .A(n195), .ZN(quantized_data[114]) );
  INV_X1 U515 ( .A(ori_data[149]), .ZN(n406) );
  OAI21_X1 U516 ( .B1(n131), .B2(n407), .A(n196), .ZN(quantized_data[113]) );
  INV_X1 U517 ( .A(ori_data[148]), .ZN(n407) );
  OAI21_X1 U518 ( .B1(n129), .B2(n408), .A(n193), .ZN(quantized_data[112]) );
  INV_X1 U519 ( .A(ori_data[147]), .ZN(n408) );
  NAND2_X1 U520 ( .A1(n391), .A2(n88), .ZN(n390) );
  OR2_X1 U521 ( .A1(ori_data[166]), .A2(ori_data[165]), .ZN(n409) );
  OAI21_X1 U522 ( .B1(n410), .B2(n411), .A(ori_data[167]), .ZN(n391) );
  NAND2_X1 U523 ( .A1(ori_data[166]), .A2(ori_data[165]), .ZN(n411) );
  NAND3_X1 U524 ( .A1(ori_data[163]), .A2(ori_data[162]), .A3(ori_data[164]), 
        .ZN(n410) );
  OAI21_X1 U525 ( .B1(n412), .B2(n231), .A(n413), .ZN(quantized_data[111]) );
  INV_X1 U526 ( .A(ori_data[141]), .ZN(n412) );
  OAI21_X1 U527 ( .B1(n107), .B2(n414), .A(n181), .ZN(quantized_data[110]) );
  INV_X1 U528 ( .A(ori_data[140]), .ZN(n414) );
  OAI21_X1 U529 ( .B1(n57), .B2(n415), .A(n98), .ZN(quantized_data[10]) );
  INV_X1 U530 ( .A(ori_data[10]), .ZN(n415) );
  OAI21_X1 U531 ( .B1(n102), .B2(n416), .A(n181), .ZN(quantized_data[109]) );
  INV_X1 U532 ( .A(ori_data[139]), .ZN(n416) );
  OAI21_X1 U533 ( .B1(n230), .B2(n417), .A(n243), .ZN(quantized_data[108]) );
  INV_X1 U534 ( .A(ori_data[138]), .ZN(n417) );
  OAI21_X1 U535 ( .B1(n108), .B2(n418), .A(n187), .ZN(quantized_data[107]) );
  INV_X1 U536 ( .A(ori_data[137]), .ZN(n418) );
  OAI21_X1 U537 ( .B1(n108), .B2(n419), .A(n185), .ZN(quantized_data[106]) );
  INV_X1 U538 ( .A(ori_data[136]), .ZN(n419) );
  OAI21_X1 U539 ( .B1(n104), .B2(n420), .A(n187), .ZN(quantized_data[105]) );
  INV_X1 U540 ( .A(ori_data[135]), .ZN(n420) );
  OAI21_X1 U541 ( .B1(n230), .B2(n421), .A(n184), .ZN(quantized_data[104]) );
  INV_X1 U542 ( .A(ori_data[134]), .ZN(n421) );
  OAI21_X1 U543 ( .B1(n105), .B2(n422), .A(n188), .ZN(quantized_data[103]) );
  INV_X1 U544 ( .A(ori_data[133]), .ZN(n422) );
  OAI21_X1 U545 ( .B1(n104), .B2(n423), .A(n243), .ZN(quantized_data[102]) );
  INV_X1 U546 ( .A(ori_data[132]), .ZN(n423) );
  OAI21_X1 U547 ( .B1(n105), .B2(n424), .A(n184), .ZN(quantized_data[101]) );
  INV_X1 U548 ( .A(ori_data[131]), .ZN(n424) );
  OAI21_X1 U549 ( .B1(n231), .B2(n425), .A(n85), .ZN(quantized_data[100]) );
  INV_X1 U550 ( .A(ori_data[130]), .ZN(n425) );
  NAND2_X1 U551 ( .A1(n413), .A2(n85), .ZN(n260) );
  OR2_X1 U552 ( .A1(ori_data[145]), .A2(ori_data[144]), .ZN(n426) );
  OAI21_X1 U553 ( .B1(n427), .B2(n428), .A(ori_data[146]), .ZN(n413) );
  NAND2_X1 U554 ( .A1(ori_data[145]), .A2(ori_data[144]), .ZN(n428) );
  NAND3_X1 U555 ( .A1(ori_data[142]), .A2(ori_data[141]), .A3(ori_data[143]), 
        .ZN(n427) );
  OAI21_X1 U556 ( .B1(n109), .B2(n429), .A(n247), .ZN(quantized_data[0]) );
  INV_X1 U557 ( .A(ori_data[0]), .ZN(n429) );
  NAND2_X1 U558 ( .A1(n385), .A2(n97), .ZN(n257) );
  OR2_X1 U559 ( .A1(ori_data[19]), .A2(ori_data[18]), .ZN(n430) );
  OAI21_X1 U560 ( .B1(n431), .B2(n432), .A(ori_data[20]), .ZN(n385) );
  NAND2_X1 U561 ( .A1(ori_data[19]), .A2(ori_data[18]), .ZN(n432) );
  NAND3_X1 U562 ( .A1(ori_data[16]), .A2(ori_data[15]), .A3(ori_data[17]), 
        .ZN(n431) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_1 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_2 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_3 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_4 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_5 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_6 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_7 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_8 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_9 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_10 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_11 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_12 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_13 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_14 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_15 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_16 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_17 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_18 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_19 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_20 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_21 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_22 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_23 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_24 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_25 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_26 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_27 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_28 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_29 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_30 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_31 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_32 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_33 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_34 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_35 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_36 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_37 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_38 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_39 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_40 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_41 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_42 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_43 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_44 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_45 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_46 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_47 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_48 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_49 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_50 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_51 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_52 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_53 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_54 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_55 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_56 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_57 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_58 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_59 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_60 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_61 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_62 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_63 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_64 ( A, B, 
        SUM );
  input [20:0] A;
  input [20:0] B;
  output [20:0] SUM;
  wire   n2, n3;
  wire   [20:2] carry;

  FA_X1 U1_20 ( .A(A[20]), .B(B[20]), .CI(carry[20]), .S(SUM[20]) );
  FA_X1 U1_19 ( .A(A[19]), .B(B[19]), .CI(carry[19]), .CO(carry[20]), .S(
        SUM[19]) );
  FA_X1 U1_18 ( .A(A[18]), .B(B[18]), .CI(carry[18]), .CO(carry[19]), .S(
        SUM[18]) );
  FA_X1 U1_17 ( .A(A[17]), .B(B[17]), .CI(carry[17]), .CO(carry[18]), .S(
        SUM[17]) );
  FA_X1 U1_16 ( .A(A[16]), .B(B[16]), .CI(carry[16]), .CO(carry[17]), .S(
        SUM[16]) );
  FA_X1 U1_15 ( .A(A[15]), .B(B[15]), .CI(carry[15]), .CO(carry[16]), .S(
        SUM[15]) );
  FA_X1 U1_14 ( .A(A[14]), .B(B[14]), .CI(carry[14]), .CO(carry[15]), .S(
        SUM[14]) );
  FA_X1 U1_13 ( .A(A[13]), .B(B[13]), .CI(carry[13]), .CO(carry[14]), .S(
        SUM[13]) );
  FA_X1 U1_12 ( .A(A[12]), .B(B[12]), .CI(carry[12]), .CO(carry[13]), .S(
        SUM[12]) );
  FA_X1 U1_11 ( .A(A[11]), .B(B[11]), .CI(carry[11]), .CO(carry[12]), .S(
        SUM[11]) );
  FA_X1 U1_10 ( .A(A[10]), .B(B[10]), .CI(carry[10]), .CO(carry[11]), .S(
        SUM[10]) );
  FA_X1 U1_9 ( .A(A[9]), .B(B[9]), .CI(carry[9]), .CO(carry[10]), .S(SUM[9])
         );
  FA_X1 U1_8 ( .A(A[8]), .B(B[8]), .CI(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  FA_X1 U1_7 ( .A(A[7]), .B(B[7]), .CI(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  FA_X1 U1_6 ( .A(A[6]), .B(B[6]), .CI(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  FA_X1 U1_5 ( .A(A[5]), .B(B[5]), .CI(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  FA_X1 U1_4 ( .A(A[4]), .B(B[4]), .CI(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  FA_X1 U1_3 ( .A(A[3]), .B(B[3]), .CI(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  FA_X1 U1_2 ( .A(A[2]), .B(B[2]), .CI(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  FA_X1 U1_1 ( .A(A[1]), .B(B[1]), .CI(n3), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(n2), .B(A[0]), .Z(SUM[0]) );
  BUF_X1 U2 ( .A(B[0]), .Z(n2) );
  AND2_X1 U3 ( .A1(n2), .A2(A[0]), .ZN(n3) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_128 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  INV_X1 U13 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U14 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U15 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U16 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U17 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U18 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_63 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n91), .B(n94), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_128 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n92), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n134), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n132), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n134), .ZN(n96) );
  INV_X1 U96 ( .A(n31), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(B[7]), .ZN(n132) );
  INV_X1 U132 ( .A(B[0]), .ZN(n133) );
  INV_X1 U133 ( .A(A[0]), .ZN(n137) );
  INV_X1 U134 ( .A(A[3]), .ZN(n136) );
  INV_X1 U135 ( .A(A[5]), .ZN(n135) );
  INV_X1 U136 ( .A(A[7]), .ZN(n134) );
  NOR2_X1 U137 ( .A1(n116), .A2(n114), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n113), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n92), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n114), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n113), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n91), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n115), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n95), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n95), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n116), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n115), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n94), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_127 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  INV_X1 U13 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U14 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U15 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U16 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U17 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U18 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_62 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n91), .B(n94), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_127 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n92), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n134), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n132), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n134), .ZN(n96) );
  INV_X1 U96 ( .A(n31), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(B[7]), .ZN(n132) );
  INV_X1 U132 ( .A(B[0]), .ZN(n133) );
  INV_X1 U133 ( .A(A[0]), .ZN(n137) );
  INV_X1 U134 ( .A(A[3]), .ZN(n136) );
  INV_X1 U135 ( .A(A[5]), .ZN(n135) );
  INV_X1 U136 ( .A(A[7]), .ZN(n134) );
  NOR2_X1 U137 ( .A1(n116), .A2(n114), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n113), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n92), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n114), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n113), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n91), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n115), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n95), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n95), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n116), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n115), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n94), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_126 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  INV_X1 U13 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U14 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U15 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U16 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U17 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U18 ( .A(A[4]), .Z(SUM[4]) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_61 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n91), .B(n94), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_126 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n92), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n134), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n132), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n134), .ZN(n96) );
  INV_X1 U96 ( .A(n31), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(B[7]), .ZN(n132) );
  INV_X1 U132 ( .A(B[0]), .ZN(n133) );
  INV_X1 U133 ( .A(A[0]), .ZN(n137) );
  INV_X1 U134 ( .A(A[3]), .ZN(n136) );
  INV_X1 U135 ( .A(A[5]), .ZN(n135) );
  INV_X1 U136 ( .A(A[7]), .ZN(n134) );
  NOR2_X1 U137 ( .A1(n116), .A2(n114), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n113), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n92), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n114), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n113), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n91), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n115), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n95), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n95), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n116), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n115), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n94), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_125 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  INV_X1 U13 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U14 ( .A(A[5]), .Z(SUM[5]) );
  BUF_X1 U15 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U16 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U17 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U18 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U19 ( .A(A[4]), .Z(SUM[4]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_60 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_125 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_124 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_59 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_124 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_123 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_58 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_123 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_122 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_57 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_122 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_121 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_56 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_121 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_120 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_55 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_120 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_119 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_54 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_119 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_118 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_53 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_118 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_117 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_52 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_117 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_116 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_51 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_116 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_115 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_50 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_115 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_114 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_49 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_114 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_113 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_48 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_113 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_112 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_47 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_112 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_111 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_46 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_111 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_110 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_45 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_110 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_109 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_44 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_109 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_108 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_43 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_108 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_107 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_42 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_107 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_106 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_41 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_106 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_105 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_40 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_105 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_104 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_39 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_104 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_103 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_38 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_103 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_102 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_37 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_102 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_101 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_36 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_101 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_100 ( A, 
        SUM, B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_35 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_100 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_99 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_34 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_99 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_98 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_33 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_98 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_97 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_32 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_97 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_96 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_31 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_96 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_95 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_30 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_95 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_94 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_29 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_94 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_93 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_28 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_93 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_92 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_27 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_92 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_91 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_26 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_91 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_90 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_25 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_90 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_89 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_24 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_89 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_88 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_23 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_88 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_87 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_22 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_87 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_86 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_21 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_86 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_85 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_20 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_85 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_84 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_19 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_84 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_83 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_18 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_83 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_82 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_17 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_82 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_81 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_16 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_81 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_80 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_15 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_80 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_79 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_14 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_79 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_78 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_13 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_78 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_77 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_12 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_77 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_76 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_11 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_76 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_75 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_10 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_75 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_74 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_9 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_74 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_73 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_8 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_73 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_72 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_7 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_72 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_71 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_6 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_71 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_70 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_5 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_70 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_69 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_4 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_69 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_68 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_3 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_68 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_67 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_2 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_67 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_66 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_1 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_66 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_65 ( A, SUM, 
        B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_ );
  input [13:0] A;
  output [13:0] SUM;
  input B_13_, B_12_, B_11_, B_10_, B_9_, B_8_, B_7_, B_6_;
  wire   n1, n2, n3, n4, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42;

  BUF_X1 U2 ( .A(A[7]), .Z(n1) );
  OR2_X1 U3 ( .A1(n18), .A2(n17), .ZN(n2) );
  INV_X1 U4 ( .A(n2), .ZN(n3) );
  INV_X1 U5 ( .A(n2), .ZN(n4) );
  INV_X1 U6 ( .A(A[6]), .ZN(n17) );
  INV_X1 U7 ( .A(n30), .ZN(n11) );
  INV_X1 U8 ( .A(n26), .ZN(n15) );
  INV_X1 U9 ( .A(n38), .ZN(n13) );
  INV_X1 U10 ( .A(n22), .ZN(n14) );
  INV_X1 U11 ( .A(n36), .ZN(n12) );
  INV_X1 U12 ( .A(n42), .ZN(n16) );
  BUF_X1 U13 ( .A(A[0]), .Z(SUM[0]) );
  BUF_X1 U14 ( .A(A[1]), .Z(SUM[1]) );
  BUF_X1 U15 ( .A(A[2]), .Z(SUM[2]) );
  BUF_X1 U16 ( .A(A[3]), .Z(SUM[3]) );
  BUF_X1 U17 ( .A(A[4]), .Z(SUM[4]) );
  INV_X1 U18 ( .A(B_6_), .ZN(n18) );
  BUF_X1 U19 ( .A(A[5]), .Z(SUM[5]) );
  XOR2_X1 U20 ( .A(n19), .B(n20), .Z(SUM[9]) );
  NOR2_X1 U21 ( .A1(n21), .A2(n22), .ZN(n20) );
  XOR2_X1 U22 ( .A(n23), .B(n24), .Z(SUM[8]) );
  NAND2_X1 U23 ( .A1(n15), .A2(n25), .ZN(n23) );
  XOR2_X1 U24 ( .A(n3), .B(n27), .Z(SUM[7]) );
  XOR2_X1 U25 ( .A(B_7_), .B(A[7]), .Z(n27) );
  AOI21_X1 U26 ( .B1(n18), .B2(n17), .A(n3), .ZN(SUM[6]) );
  XOR2_X1 U27 ( .A(n28), .B(n29), .Z(SUM[13]) );
  XOR2_X1 U28 ( .A(B_13_), .B(A[13]), .Z(n29) );
  OAI21_X1 U29 ( .B1(n30), .B2(n31), .A(n32), .ZN(n28) );
  XOR2_X1 U30 ( .A(n33), .B(n31), .Z(SUM[12]) );
  AOI21_X1 U31 ( .B1(n12), .B2(n34), .A(n35), .ZN(n31) );
  NAND2_X1 U32 ( .A1(n11), .A2(n32), .ZN(n33) );
  NAND2_X1 U33 ( .A1(B_12_), .A2(A[12]), .ZN(n32) );
  NOR2_X1 U34 ( .A1(B_12_), .A2(A[12]), .ZN(n30) );
  XOR2_X1 U35 ( .A(n34), .B(n37), .Z(SUM[11]) );
  NOR2_X1 U36 ( .A1(n35), .A2(n36), .ZN(n37) );
  NOR2_X1 U37 ( .A1(B_11_), .A2(A[11]), .ZN(n36) );
  AND2_X1 U38 ( .A1(B_11_), .A2(A[11]), .ZN(n35) );
  OAI21_X1 U39 ( .B1(n38), .B2(n39), .A(n40), .ZN(n34) );
  XOR2_X1 U40 ( .A(n41), .B(n39), .Z(SUM[10]) );
  AOI21_X1 U41 ( .B1(n19), .B2(n14), .A(n21), .ZN(n39) );
  AND2_X1 U42 ( .A1(B_9_), .A2(A[9]), .ZN(n21) );
  NOR2_X1 U43 ( .A1(B_9_), .A2(A[9]), .ZN(n22) );
  OAI21_X1 U44 ( .B1(n24), .B2(n26), .A(n25), .ZN(n19) );
  NAND2_X1 U45 ( .A1(B_8_), .A2(A[8]), .ZN(n25) );
  NOR2_X1 U46 ( .A1(B_8_), .A2(A[8]), .ZN(n26) );
  AOI21_X1 U47 ( .B1(n4), .B2(n1), .A(n16), .ZN(n24) );
  OAI21_X1 U48 ( .B1(n4), .B2(n1), .A(B_7_), .ZN(n42) );
  NAND2_X1 U49 ( .A1(n13), .A2(n40), .ZN(n41) );
  NAND2_X1 U50 ( .A1(B_10_), .A2(A[10]), .ZN(n40) );
  NOR2_X1 U51 ( .A1(B_10_), .A2(A[10]), .ZN(n38) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_0 ( A, B, 
        PRODUCT );
  input [7:0] A;
  input [7:0] B;
  output [15:0] PRODUCT;
  wire   ab_7__7_, ab_7__6_, ab_7__5_, ab_7__4_, ab_7__3_, ab_7__2_, ab_7__1_,
         ab_7__0_, ab_6__7_, ab_6__6_, ab_6__5_, ab_6__4_, ab_6__3_, ab_6__2_,
         ab_6__1_, ab_6__0_, ab_5__7_, ab_5__6_, ab_5__5_, ab_5__4_, ab_5__3_,
         ab_5__2_, ab_5__1_, ab_5__0_, ab_4__7_, ab_4__6_, ab_4__5_, ab_4__4_,
         ab_4__3_, ab_4__2_, ab_4__1_, ab_4__0_, ab_3__7_, ab_3__6_, ab_3__5_,
         ab_3__4_, ab_3__3_, ab_3__2_, ab_3__1_, ab_3__0_, ab_2__7_, ab_2__6_,
         ab_2__5_, ab_2__4_, ab_2__3_, ab_2__2_, ab_2__1_, ab_2__0_, ab_1__7_,
         ab_1__6_, ab_1__5_, ab_1__4_, ab_1__3_, ab_1__2_, ab_1__1_, ab_1__0_,
         ab_0__7_, ab_0__6_, ab_0__5_, ab_0__4_, ab_0__3_, ab_0__2_, ab_0__1_,
         CARRYB_7__7_, CARRYB_7__6_, CARRYB_7__5_, CARRYB_7__4_, CARRYB_7__3_,
         CARRYB_7__2_, CARRYB_7__1_, CARRYB_7__0_, CARRYB_6__6_, CARRYB_6__5_,
         CARRYB_6__4_, CARRYB_6__3_, CARRYB_6__2_, CARRYB_6__1_, CARRYB_6__0_,
         CARRYB_5__6_, CARRYB_5__5_, CARRYB_5__4_, CARRYB_5__3_, CARRYB_5__2_,
         CARRYB_5__1_, CARRYB_5__0_, CARRYB_4__6_, CARRYB_4__5_, CARRYB_4__4_,
         CARRYB_4__3_, CARRYB_4__2_, CARRYB_4__1_, CARRYB_4__0_, CARRYB_3__6_,
         CARRYB_3__5_, CARRYB_3__4_, CARRYB_3__3_, CARRYB_3__2_, CARRYB_3__1_,
         CARRYB_3__0_, CARRYB_2__6_, CARRYB_2__5_, CARRYB_2__4_, CARRYB_2__3_,
         CARRYB_2__2_, CARRYB_2__1_, CARRYB_2__0_, SUMB_7__7_, SUMB_7__6_,
         SUMB_7__5_, SUMB_7__4_, SUMB_7__3_, SUMB_7__2_, SUMB_7__1_,
         SUMB_7__0_, SUMB_6__6_, SUMB_6__5_, SUMB_6__4_, SUMB_6__3_,
         SUMB_6__2_, SUMB_6__1_, SUMB_5__6_, SUMB_5__5_, SUMB_5__4_,
         SUMB_5__3_, SUMB_5__2_, SUMB_5__1_, SUMB_4__6_, SUMB_4__5_,
         SUMB_4__4_, SUMB_4__3_, SUMB_4__2_, SUMB_4__1_, SUMB_3__6_,
         SUMB_3__5_, SUMB_3__4_, SUMB_3__3_, SUMB_3__2_, SUMB_3__1_,
         SUMB_2__6_, SUMB_2__5_, SUMB_2__4_, SUMB_2__3_, SUMB_2__2_,
         SUMB_2__1_, A1_13_, A1_5_, A1_4_, A1_3_, A1_2_, A1_1_, A1_0_, A2_6_,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87,
         n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137;

  FA_X1 S14_7_0 ( .A(A[7]), .B(B[7]), .CI(SUMB_7__0_), .CO(A2_6_), .S(A1_5_)
         );
  FA_X1 S4_0 ( .A(ab_7__0_), .B(CARRYB_6__0_), .CI(SUMB_6__1_), .CO(
        CARRYB_7__0_), .S(SUMB_7__0_) );
  FA_X1 S4_1 ( .A(ab_7__1_), .B(CARRYB_6__1_), .CI(SUMB_6__2_), .CO(
        CARRYB_7__1_), .S(SUMB_7__1_) );
  FA_X1 S4_2 ( .A(ab_7__2_), .B(CARRYB_6__2_), .CI(SUMB_6__3_), .CO(
        CARRYB_7__2_), .S(SUMB_7__2_) );
  FA_X1 S4_3 ( .A(ab_7__3_), .B(CARRYB_6__3_), .CI(SUMB_6__4_), .CO(
        CARRYB_7__3_), .S(SUMB_7__3_) );
  FA_X1 S4_4 ( .A(ab_7__4_), .B(CARRYB_6__4_), .CI(SUMB_6__5_), .CO(
        CARRYB_7__4_), .S(SUMB_7__4_) );
  FA_X1 S4_5 ( .A(ab_7__5_), .B(CARRYB_6__5_), .CI(SUMB_6__6_), .CO(
        CARRYB_7__5_), .S(SUMB_7__5_) );
  FA_X1 S5_6 ( .A(ab_7__6_), .B(CARRYB_6__6_), .CI(ab_6__7_), .CO(CARRYB_7__6_), .S(SUMB_7__6_) );
  FA_X1 S14_7 ( .A(n94), .B(n91), .CI(ab_7__7_), .CO(CARRYB_7__7_), .S(
        SUMB_7__7_) );
  FA_X1 S1_6_0 ( .A(ab_6__0_), .B(CARRYB_5__0_), .CI(SUMB_5__1_), .CO(
        CARRYB_6__0_), .S(A1_4_) );
  FA_X1 S2_6_1 ( .A(ab_6__1_), .B(CARRYB_5__1_), .CI(SUMB_5__2_), .CO(
        CARRYB_6__1_), .S(SUMB_6__1_) );
  FA_X1 S2_6_2 ( .A(ab_6__2_), .B(CARRYB_5__2_), .CI(SUMB_5__3_), .CO(
        CARRYB_6__2_), .S(SUMB_6__2_) );
  FA_X1 S2_6_3 ( .A(ab_6__3_), .B(CARRYB_5__3_), .CI(SUMB_5__4_), .CO(
        CARRYB_6__3_), .S(SUMB_6__3_) );
  FA_X1 S2_6_4 ( .A(ab_6__4_), .B(CARRYB_5__4_), .CI(SUMB_5__5_), .CO(
        CARRYB_6__4_), .S(SUMB_6__4_) );
  FA_X1 S2_6_5 ( .A(ab_6__5_), .B(CARRYB_5__5_), .CI(SUMB_5__6_), .CO(
        CARRYB_6__5_), .S(SUMB_6__5_) );
  FA_X1 S3_6_6 ( .A(ab_6__6_), .B(CARRYB_5__6_), .CI(ab_5__7_), .CO(
        CARRYB_6__6_), .S(SUMB_6__6_) );
  FA_X1 S1_5_0 ( .A(ab_5__0_), .B(CARRYB_4__0_), .CI(SUMB_4__1_), .CO(
        CARRYB_5__0_), .S(A1_3_) );
  FA_X1 S2_5_1 ( .A(ab_5__1_), .B(CARRYB_4__1_), .CI(SUMB_4__2_), .CO(
        CARRYB_5__1_), .S(SUMB_5__1_) );
  FA_X1 S2_5_2 ( .A(ab_5__2_), .B(CARRYB_4__2_), .CI(SUMB_4__3_), .CO(
        CARRYB_5__2_), .S(SUMB_5__2_) );
  FA_X1 S2_5_3 ( .A(ab_5__3_), .B(CARRYB_4__3_), .CI(SUMB_4__4_), .CO(
        CARRYB_5__3_), .S(SUMB_5__3_) );
  FA_X1 S2_5_4 ( .A(ab_5__4_), .B(CARRYB_4__4_), .CI(SUMB_4__5_), .CO(
        CARRYB_5__4_), .S(SUMB_5__4_) );
  FA_X1 S2_5_5 ( .A(ab_5__5_), .B(CARRYB_4__5_), .CI(SUMB_4__6_), .CO(
        CARRYB_5__5_), .S(SUMB_5__5_) );
  FA_X1 S3_5_6 ( .A(ab_5__6_), .B(CARRYB_4__6_), .CI(ab_4__7_), .CO(
        CARRYB_5__6_), .S(SUMB_5__6_) );
  FA_X1 S1_4_0 ( .A(ab_4__0_), .B(CARRYB_3__0_), .CI(SUMB_3__1_), .CO(
        CARRYB_4__0_), .S(A1_2_) );
  FA_X1 S2_4_1 ( .A(ab_4__1_), .B(CARRYB_3__1_), .CI(SUMB_3__2_), .CO(
        CARRYB_4__1_), .S(SUMB_4__1_) );
  FA_X1 S2_4_2 ( .A(ab_4__2_), .B(CARRYB_3__2_), .CI(SUMB_3__3_), .CO(
        CARRYB_4__2_), .S(SUMB_4__2_) );
  FA_X1 S2_4_3 ( .A(ab_4__3_), .B(CARRYB_3__3_), .CI(SUMB_3__4_), .CO(
        CARRYB_4__3_), .S(SUMB_4__3_) );
  FA_X1 S2_4_4 ( .A(ab_4__4_), .B(CARRYB_3__4_), .CI(SUMB_3__5_), .CO(
        CARRYB_4__4_), .S(SUMB_4__4_) );
  FA_X1 S2_4_5 ( .A(ab_4__5_), .B(CARRYB_3__5_), .CI(SUMB_3__6_), .CO(
        CARRYB_4__5_), .S(SUMB_4__5_) );
  FA_X1 S3_4_6 ( .A(ab_4__6_), .B(CARRYB_3__6_), .CI(ab_3__7_), .CO(
        CARRYB_4__6_), .S(SUMB_4__6_) );
  FA_X1 S1_3_0 ( .A(ab_3__0_), .B(CARRYB_2__0_), .CI(SUMB_2__1_), .CO(
        CARRYB_3__0_), .S(A1_1_) );
  FA_X1 S2_3_1 ( .A(ab_3__1_), .B(CARRYB_2__1_), .CI(SUMB_2__2_), .CO(
        CARRYB_3__1_), .S(SUMB_3__1_) );
  FA_X1 S2_3_2 ( .A(ab_3__2_), .B(CARRYB_2__2_), .CI(SUMB_2__3_), .CO(
        CARRYB_3__2_), .S(SUMB_3__2_) );
  FA_X1 S2_3_3 ( .A(ab_3__3_), .B(CARRYB_2__3_), .CI(SUMB_2__4_), .CO(
        CARRYB_3__3_), .S(SUMB_3__3_) );
  FA_X1 S2_3_4 ( .A(ab_3__4_), .B(CARRYB_2__4_), .CI(SUMB_2__5_), .CO(
        CARRYB_3__4_), .S(SUMB_3__4_) );
  FA_X1 S2_3_5 ( .A(ab_3__5_), .B(CARRYB_2__5_), .CI(SUMB_2__6_), .CO(
        CARRYB_3__5_), .S(SUMB_3__5_) );
  FA_X1 S3_3_6 ( .A(ab_3__6_), .B(CARRYB_2__6_), .CI(ab_2__7_), .CO(
        CARRYB_3__6_), .S(SUMB_3__6_) );
  FA_X1 S1_2_0 ( .A(ab_2__0_), .B(n8), .CI(n15), .CO(CARRYB_2__0_), .S(A1_0_)
         );
  FA_X1 S2_2_1 ( .A(ab_2__1_), .B(n7), .CI(n14), .CO(CARRYB_2__1_), .S(
        SUMB_2__1_) );
  FA_X1 S2_2_2 ( .A(ab_2__2_), .B(n6), .CI(n13), .CO(CARRYB_2__2_), .S(
        SUMB_2__2_) );
  FA_X1 S2_2_3 ( .A(ab_2__3_), .B(n5), .CI(n12), .CO(CARRYB_2__3_), .S(
        SUMB_2__3_) );
  FA_X1 S2_2_4 ( .A(ab_2__4_), .B(n4), .CI(n11), .CO(CARRYB_2__4_), .S(
        SUMB_2__4_) );
  FA_X1 S2_2_5 ( .A(ab_2__5_), .B(n3), .CI(n10), .CO(CARRYB_2__5_), .S(
        SUMB_2__5_) );
  FA_X1 S3_2_6 ( .A(ab_2__6_), .B(n9), .CI(ab_1__7_), .CO(CARRYB_2__6_), .S(
        SUMB_2__6_) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_65 FS_1 ( .A({
        A1_13_, n123, n118, n122, n127, n121, n119, n128, A1_5_, A1_4_, A1_3_, 
        A1_2_, A1_1_, A1_0_}), .SUM(PRODUCT[15:2]), .B_13_(n131), .B_12_(n126), 
        .B_11_(n130), .B_10_(n125), .B_9_(n129), .B_8_(n124), .B_7_(n120), 
        .B_6_(A2_6_) );
  AND2_X1 U2 ( .A1(ab_0__6_), .A2(ab_1__5_), .ZN(n3) );
  AND2_X1 U3 ( .A1(ab_0__5_), .A2(ab_1__4_), .ZN(n4) );
  AND2_X1 U4 ( .A1(ab_0__4_), .A2(ab_1__3_), .ZN(n5) );
  AND2_X1 U5 ( .A1(ab_0__3_), .A2(ab_1__2_), .ZN(n6) );
  AND2_X1 U6 ( .A1(ab_0__2_), .A2(ab_1__1_), .ZN(n7) );
  AND2_X1 U7 ( .A1(ab_0__1_), .A2(ab_1__0_), .ZN(n8) );
  AND2_X1 U8 ( .A1(ab_0__7_), .A2(ab_1__6_), .ZN(n9) );
  XOR2_X1 U9 ( .A(ab_1__6_), .B(ab_0__7_), .Z(n10) );
  XOR2_X1 U10 ( .A(ab_1__5_), .B(ab_0__6_), .Z(n11) );
  XOR2_X1 U11 ( .A(ab_1__4_), .B(ab_0__5_), .Z(n12) );
  XOR2_X1 U12 ( .A(ab_1__3_), .B(ab_0__4_), .Z(n13) );
  XOR2_X1 U13 ( .A(ab_1__2_), .B(ab_0__3_), .Z(n14) );
  XOR2_X1 U14 ( .A(ab_1__1_), .B(ab_0__2_), .Z(n15) );
  CLKBUF_X1 U15 ( .A(n95), .Z(n16) );
  CLKBUF_X1 U16 ( .A(A[4]), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n44), .Z(n18) );
  CLKBUF_X1 U18 ( .A(A[2]), .Z(n19) );
  CLKBUF_X1 U19 ( .A(n51), .Z(n20) );
  CLKBUF_X1 U20 ( .A(A[1]), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n58), .Z(n22) );
  CLKBUF_X1 U22 ( .A(B[6]), .Z(n23) );
  CLKBUF_X1 U23 ( .A(B[5]), .Z(n24) );
  CLKBUF_X1 U24 ( .A(B[4]), .Z(n25) );
  CLKBUF_X1 U25 ( .A(B[3]), .Z(n26) );
  CLKBUF_X1 U26 ( .A(n133), .Z(n27) );
  CLKBUF_X1 U27 ( .A(B[1]), .Z(n28) );
  CLKBUF_X1 U28 ( .A(A[6]), .Z(n29) );
  CLKBUF_X1 U29 ( .A(B[2]), .Z(n30) );
  CLKBUF_X1 U30 ( .A(n132), .Z(n31) );
  CLKBUF_X1 U31 ( .A(n40), .Z(n32) );
  CLKBUF_X1 U32 ( .A(n135), .Z(n33) );
  CLKBUF_X1 U33 ( .A(n47), .Z(n34) );
  CLKBUF_X1 U34 ( .A(n136), .Z(n35) );
  CLKBUF_X1 U35 ( .A(n54), .Z(n36) );
  CLKBUF_X1 U36 ( .A(n137), .Z(n37) );
  CLKBUF_X1 U37 ( .A(n27), .Z(n38) );
  CLKBUF_X1 U38 ( .A(n82), .Z(n39) );
  INV_X1 U39 ( .A(n17), .ZN(n40) );
  INV_X1 U40 ( .A(n40), .ZN(n41) );
  INV_X1 U41 ( .A(n17), .ZN(n42) );
  INV_X1 U42 ( .A(n41), .ZN(n43) );
  INV_X1 U43 ( .A(n135), .ZN(n44) );
  INV_X1 U44 ( .A(n18), .ZN(n45) );
  INV_X1 U45 ( .A(n18), .ZN(n46) );
  INV_X1 U46 ( .A(n19), .ZN(n47) );
  INV_X1 U47 ( .A(n47), .ZN(n48) );
  INV_X1 U48 ( .A(n19), .ZN(n49) );
  INV_X1 U49 ( .A(n48), .ZN(n50) );
  INV_X1 U50 ( .A(n136), .ZN(n51) );
  INV_X1 U51 ( .A(n20), .ZN(n52) );
  INV_X1 U52 ( .A(n20), .ZN(n53) );
  INV_X1 U53 ( .A(n21), .ZN(n54) );
  INV_X1 U54 ( .A(n54), .ZN(n55) );
  INV_X1 U55 ( .A(n21), .ZN(n56) );
  INV_X1 U56 ( .A(n55), .ZN(n57) );
  INV_X1 U57 ( .A(n137), .ZN(n58) );
  INV_X1 U58 ( .A(n22), .ZN(n59) );
  INV_X1 U59 ( .A(n22), .ZN(n60) );
  INV_X1 U60 ( .A(n23), .ZN(n61) );
  INV_X1 U61 ( .A(n61), .ZN(n62) );
  INV_X1 U62 ( .A(n23), .ZN(n63) );
  INV_X1 U63 ( .A(n62), .ZN(n64) );
  INV_X1 U64 ( .A(n24), .ZN(n65) );
  INV_X1 U65 ( .A(n65), .ZN(n66) );
  INV_X1 U66 ( .A(n24), .ZN(n67) );
  INV_X1 U67 ( .A(n66), .ZN(n68) );
  INV_X1 U68 ( .A(n25), .ZN(n69) );
  INV_X1 U69 ( .A(n69), .ZN(n70) );
  INV_X1 U70 ( .A(n25), .ZN(n71) );
  INV_X1 U71 ( .A(n70), .ZN(n72) );
  INV_X1 U72 ( .A(n26), .ZN(n73) );
  INV_X1 U73 ( .A(n73), .ZN(n74) );
  INV_X1 U74 ( .A(n26), .ZN(n75) );
  INV_X1 U75 ( .A(n74), .ZN(n76) );
  INV_X1 U76 ( .A(n27), .ZN(n77) );
  INV_X1 U77 ( .A(n28), .ZN(n78) );
  INV_X1 U78 ( .A(n78), .ZN(n79) );
  INV_X1 U79 ( .A(n28), .ZN(n80) );
  INV_X1 U80 ( .A(n79), .ZN(n81) );
  INV_X1 U81 ( .A(n29), .ZN(n82) );
  INV_X1 U82 ( .A(n82), .ZN(n83) );
  INV_X1 U83 ( .A(n29), .ZN(n84) );
  INV_X1 U84 ( .A(n83), .ZN(n85) );
  INV_X1 U85 ( .A(n30), .ZN(n86) );
  INV_X1 U86 ( .A(n86), .ZN(n87) );
  INV_X1 U87 ( .A(n30), .ZN(n88) );
  INV_X1 U88 ( .A(n87), .ZN(n89) );
  INV_X1 U89 ( .A(n132), .ZN(n90) );
  INV_X1 U90 ( .A(n90), .ZN(n91) );
  INV_X1 U91 ( .A(n90), .ZN(n92) );
  INV_X1 U92 ( .A(n134), .ZN(n93) );
  INV_X1 U93 ( .A(n93), .ZN(n94) );
  INV_X1 U94 ( .A(n93), .ZN(n95) );
  INV_X1 U95 ( .A(n31), .ZN(n96) );
  INV_X1 U96 ( .A(n134), .ZN(n97) );
  INV_X1 U97 ( .A(n41), .ZN(n98) );
  INV_X1 U98 ( .A(n44), .ZN(n99) );
  INV_X1 U99 ( .A(n48), .ZN(n100) );
  INV_X1 U100 ( .A(n51), .ZN(n101) );
  INV_X1 U101 ( .A(n55), .ZN(n102) );
  INV_X1 U102 ( .A(n58), .ZN(n103) );
  INV_X1 U103 ( .A(n62), .ZN(n104) );
  INV_X1 U104 ( .A(n66), .ZN(n105) );
  INV_X1 U105 ( .A(n70), .ZN(n106) );
  INV_X1 U106 ( .A(n74), .ZN(n107) );
  INV_X1 U107 ( .A(n77), .ZN(n108) );
  INV_X1 U108 ( .A(n77), .ZN(n109) );
  INV_X1 U109 ( .A(n79), .ZN(n110) );
  INV_X1 U110 ( .A(n83), .ZN(n111) );
  INV_X1 U111 ( .A(n87), .ZN(n112) );
  INV_X1 U112 ( .A(n96), .ZN(n113) );
  INV_X1 U113 ( .A(n96), .ZN(n114) );
  INV_X1 U114 ( .A(n97), .ZN(n115) );
  INV_X1 U115 ( .A(n97), .ZN(n116) );
  XOR2_X1 U116 ( .A(ab_1__0_), .B(ab_0__1_), .Z(PRODUCT[1]) );
  XOR2_X1 U117 ( .A(CARRYB_7__5_), .B(SUMB_7__6_), .Z(n118) );
  XOR2_X1 U118 ( .A(CARRYB_7__1_), .B(SUMB_7__2_), .Z(n119) );
  AND2_X1 U119 ( .A1(CARRYB_7__0_), .A2(SUMB_7__1_), .ZN(n120) );
  XOR2_X1 U120 ( .A(CARRYB_7__2_), .B(SUMB_7__3_), .Z(n121) );
  XOR2_X1 U121 ( .A(CARRYB_7__4_), .B(SUMB_7__5_), .Z(n122) );
  XOR2_X1 U122 ( .A(CARRYB_7__6_), .B(SUMB_7__7_), .Z(n123) );
  AND2_X1 U123 ( .A1(CARRYB_7__1_), .A2(SUMB_7__2_), .ZN(n124) );
  AND2_X1 U124 ( .A1(CARRYB_7__3_), .A2(SUMB_7__4_), .ZN(n125) );
  AND2_X1 U125 ( .A1(CARRYB_7__5_), .A2(SUMB_7__6_), .ZN(n126) );
  XOR2_X1 U126 ( .A(CARRYB_7__3_), .B(SUMB_7__4_), .Z(n127) );
  XOR2_X1 U127 ( .A(CARRYB_7__0_), .B(SUMB_7__1_), .Z(n128) );
  AND2_X1 U128 ( .A1(CARRYB_7__2_), .A2(SUMB_7__3_), .ZN(n129) );
  AND2_X1 U129 ( .A1(CARRYB_7__4_), .A2(SUMB_7__5_), .ZN(n130) );
  AND2_X1 U130 ( .A1(CARRYB_7__6_), .A2(SUMB_7__7_), .ZN(n131) );
  INV_X1 U131 ( .A(A[7]), .ZN(n134) );
  INV_X1 U132 ( .A(B[7]), .ZN(n132) );
  INV_X1 U133 ( .A(B[0]), .ZN(n133) );
  INV_X1 U134 ( .A(A[0]), .ZN(n137) );
  INV_X1 U135 ( .A(A[3]), .ZN(n136) );
  INV_X1 U136 ( .A(A[5]), .ZN(n135) );
  NOR2_X1 U137 ( .A1(n114), .A2(n116), .ZN(ab_7__7_) );
  NOR2_X1 U138 ( .A1(B[6]), .A2(n16), .ZN(ab_7__6_) );
  NOR2_X1 U139 ( .A1(B[5]), .A2(n115), .ZN(ab_7__5_) );
  NOR2_X1 U140 ( .A1(B[4]), .A2(n95), .ZN(ab_7__4_) );
  NOR2_X1 U141 ( .A1(B[3]), .A2(n116), .ZN(ab_7__3_) );
  NOR2_X1 U142 ( .A1(B[2]), .A2(n16), .ZN(ab_7__2_) );
  NOR2_X1 U143 ( .A1(B[1]), .A2(n115), .ZN(ab_7__1_) );
  NOR2_X1 U144 ( .A1(B[0]), .A2(n94), .ZN(ab_7__0_) );
  NOR2_X1 U145 ( .A1(A[6]), .A2(n113), .ZN(ab_6__7_) );
  NOR2_X1 U146 ( .A1(n84), .A2(n63), .ZN(ab_6__6_) );
  NOR2_X1 U147 ( .A1(n111), .A2(n67), .ZN(ab_6__5_) );
  NOR2_X1 U148 ( .A1(n39), .A2(n71), .ZN(ab_6__4_) );
  NOR2_X1 U149 ( .A1(n85), .A2(n75), .ZN(ab_6__3_) );
  NOR2_X1 U150 ( .A1(n39), .A2(n88), .ZN(ab_6__2_) );
  NOR2_X1 U151 ( .A1(n84), .A2(n80), .ZN(ab_6__1_) );
  NOR2_X1 U152 ( .A1(n111), .A2(n108), .ZN(ab_6__0_) );
  NOR2_X1 U153 ( .A1(A[5]), .A2(n92), .ZN(ab_5__7_) );
  NOR2_X1 U154 ( .A1(n104), .A2(n45), .ZN(ab_5__6_) );
  NOR2_X1 U155 ( .A1(n105), .A2(n33), .ZN(ab_5__5_) );
  NOR2_X1 U156 ( .A1(n106), .A2(n99), .ZN(ab_5__4_) );
  NOR2_X1 U157 ( .A1(n107), .A2(n33), .ZN(ab_5__3_) );
  NOR2_X1 U158 ( .A1(n112), .A2(n45), .ZN(ab_5__2_) );
  NOR2_X1 U159 ( .A1(n110), .A2(n99), .ZN(ab_5__1_) );
  NOR2_X1 U160 ( .A1(n109), .A2(n46), .ZN(ab_5__0_) );
  NOR2_X1 U161 ( .A1(A[4]), .A2(n92), .ZN(ab_4__7_) );
  NOR2_X1 U162 ( .A1(n64), .A2(n42), .ZN(ab_4__6_) );
  NOR2_X1 U163 ( .A1(n68), .A2(n98), .ZN(ab_4__5_) );
  NOR2_X1 U164 ( .A1(n72), .A2(n32), .ZN(ab_4__4_) );
  NOR2_X1 U165 ( .A1(n76), .A2(n42), .ZN(ab_4__3_) );
  NOR2_X1 U166 ( .A1(n89), .A2(n98), .ZN(ab_4__2_) );
  NOR2_X1 U167 ( .A1(n81), .A2(n43), .ZN(ab_4__1_) );
  NOR2_X1 U168 ( .A1(n108), .A2(n32), .ZN(ab_4__0_) );
  NOR2_X1 U169 ( .A1(A[3]), .A2(n114), .ZN(ab_3__7_) );
  NOR2_X1 U170 ( .A1(n64), .A2(n52), .ZN(ab_3__6_) );
  NOR2_X1 U171 ( .A1(n68), .A2(n35), .ZN(ab_3__5_) );
  NOR2_X1 U172 ( .A1(n72), .A2(n52), .ZN(ab_3__4_) );
  NOR2_X1 U173 ( .A1(n76), .A2(n101), .ZN(ab_3__3_) );
  NOR2_X1 U174 ( .A1(n89), .A2(n53), .ZN(ab_3__2_) );
  NOR2_X1 U175 ( .A1(n81), .A2(n101), .ZN(ab_3__1_) );
  NOR2_X1 U176 ( .A1(n109), .A2(n35), .ZN(ab_3__0_) );
  NOR2_X1 U177 ( .A1(A[2]), .A2(n113), .ZN(ab_2__7_) );
  NOR2_X1 U178 ( .A1(n104), .A2(n34), .ZN(ab_2__6_) );
  NOR2_X1 U179 ( .A1(n105), .A2(n49), .ZN(ab_2__5_) );
  NOR2_X1 U180 ( .A1(n106), .A2(n100), .ZN(ab_2__4_) );
  NOR2_X1 U181 ( .A1(n107), .A2(n50), .ZN(ab_2__3_) );
  NOR2_X1 U182 ( .A1(n112), .A2(n34), .ZN(ab_2__2_) );
  NOR2_X1 U183 ( .A1(n110), .A2(n100), .ZN(ab_2__1_) );
  NOR2_X1 U184 ( .A1(n38), .A2(n49), .ZN(ab_2__0_) );
  NOR2_X1 U185 ( .A1(A[1]), .A2(n31), .ZN(ab_1__7_) );
  NOR2_X1 U186 ( .A1(n61), .A2(n36), .ZN(ab_1__6_) );
  NOR2_X1 U187 ( .A1(n67), .A2(n56), .ZN(ab_1__5_) );
  NOR2_X1 U188 ( .A1(n69), .A2(n102), .ZN(ab_1__4_) );
  NOR2_X1 U189 ( .A1(n75), .A2(n57), .ZN(ab_1__3_) );
  NOR2_X1 U190 ( .A1(n86), .A2(n36), .ZN(ab_1__2_) );
  NOR2_X1 U191 ( .A1(n80), .A2(n102), .ZN(ab_1__1_) );
  NOR2_X1 U192 ( .A1(n133), .A2(n56), .ZN(ab_1__0_) );
  NOR2_X1 U193 ( .A1(A[0]), .A2(n91), .ZN(ab_0__7_) );
  NOR2_X1 U194 ( .A1(n63), .A2(n59), .ZN(ab_0__6_) );
  NOR2_X1 U195 ( .A1(n65), .A2(n37), .ZN(ab_0__5_) );
  NOR2_X1 U196 ( .A1(n71), .A2(n103), .ZN(ab_0__4_) );
  NOR2_X1 U197 ( .A1(n73), .A2(n60), .ZN(ab_0__3_) );
  NOR2_X1 U198 ( .A1(n88), .A2(n37), .ZN(ab_0__2_) );
  NOR2_X1 U199 ( .A1(n78), .A2(n103), .ZN(ab_0__1_) );
  NOR2_X1 U200 ( .A1(n38), .A2(n59), .ZN(PRODUCT[0]) );
  INV_X1 U202 ( .A(CARRYB_7__7_), .ZN(A1_13_) );
endmodule


module systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8 ( clk, srstn, 
        alu_start, cycle_num, sram_rdata_w0, sram_rdata_w1, sram_rdata_d0, 
        sram_rdata_d1, matrix_index, mul_outcome );
  input [8:0] cycle_num;
  input [31:0] sram_rdata_w0;
  input [31:0] sram_rdata_w1;
  input [31:0] sram_rdata_d0;
  input [31:0] sram_rdata_d1;
  input [5:0] matrix_index;
  output [167:0] mul_outcome;
  input clk, srstn, alu_start;
  wire   weight_queue_0__0__7_, weight_queue_0__0__6_, weight_queue_0__0__5_,
         weight_queue_0__0__4_, weight_queue_0__0__3_, weight_queue_0__0__2_,
         weight_queue_0__0__1_, weight_queue_0__0__0_, weight_queue_0__1__7_,
         weight_queue_0__1__6_, weight_queue_0__1__5_, weight_queue_0__1__4_,
         weight_queue_0__1__3_, weight_queue_0__1__2_, weight_queue_0__1__1_,
         weight_queue_0__1__0_, weight_queue_0__2__7_, weight_queue_0__2__6_,
         weight_queue_0__2__5_, weight_queue_0__2__4_, weight_queue_0__2__3_,
         weight_queue_0__2__2_, weight_queue_0__2__1_, weight_queue_0__2__0_,
         weight_queue_0__3__7_, weight_queue_0__3__6_, weight_queue_0__3__5_,
         weight_queue_0__3__4_, weight_queue_0__3__3_, weight_queue_0__3__2_,
         weight_queue_0__3__1_, weight_queue_0__3__0_, weight_queue_0__4__7_,
         weight_queue_0__4__6_, weight_queue_0__4__5_, weight_queue_0__4__4_,
         weight_queue_0__4__3_, weight_queue_0__4__2_, weight_queue_0__4__1_,
         weight_queue_0__4__0_, weight_queue_0__5__7_, weight_queue_0__5__6_,
         weight_queue_0__5__5_, weight_queue_0__5__4_, weight_queue_0__5__3_,
         weight_queue_0__5__2_, weight_queue_0__5__1_, weight_queue_0__5__0_,
         weight_queue_0__6__7_, weight_queue_0__6__6_, weight_queue_0__6__5_,
         weight_queue_0__6__4_, weight_queue_0__6__3_, weight_queue_0__6__2_,
         weight_queue_0__6__1_, weight_queue_0__6__0_, weight_queue_0__7__7_,
         weight_queue_0__7__6_, weight_queue_0__7__5_, weight_queue_0__7__4_,
         weight_queue_0__7__3_, weight_queue_0__7__2_, weight_queue_0__7__1_,
         weight_queue_0__7__0_, weight_queue_1__0__7_, weight_queue_1__0__6_,
         weight_queue_1__0__5_, weight_queue_1__0__4_, weight_queue_1__0__3_,
         weight_queue_1__0__2_, weight_queue_1__0__1_, weight_queue_1__0__0_,
         weight_queue_1__1__7_, weight_queue_1__1__6_, weight_queue_1__1__5_,
         weight_queue_1__1__4_, weight_queue_1__1__3_, weight_queue_1__1__2_,
         weight_queue_1__1__1_, weight_queue_1__1__0_, weight_queue_1__2__7_,
         weight_queue_1__2__6_, weight_queue_1__2__5_, weight_queue_1__2__4_,
         weight_queue_1__2__3_, weight_queue_1__2__2_, weight_queue_1__2__1_,
         weight_queue_1__2__0_, weight_queue_1__3__7_, weight_queue_1__3__6_,
         weight_queue_1__3__5_, weight_queue_1__3__4_, weight_queue_1__3__3_,
         weight_queue_1__3__2_, weight_queue_1__3__1_, weight_queue_1__3__0_,
         weight_queue_1__4__7_, weight_queue_1__4__6_, weight_queue_1__4__5_,
         weight_queue_1__4__4_, weight_queue_1__4__3_, weight_queue_1__4__2_,
         weight_queue_1__4__1_, weight_queue_1__4__0_, weight_queue_1__5__7_,
         weight_queue_1__5__6_, weight_queue_1__5__5_, weight_queue_1__5__4_,
         weight_queue_1__5__3_, weight_queue_1__5__2_, weight_queue_1__5__1_,
         weight_queue_1__5__0_, weight_queue_1__6__7_, weight_queue_1__6__6_,
         weight_queue_1__6__5_, weight_queue_1__6__4_, weight_queue_1__6__3_,
         weight_queue_1__6__2_, weight_queue_1__6__1_, weight_queue_1__6__0_,
         weight_queue_1__7__7_, weight_queue_1__7__6_, weight_queue_1__7__5_,
         weight_queue_1__7__4_, weight_queue_1__7__3_, weight_queue_1__7__2_,
         weight_queue_1__7__1_, weight_queue_1__7__0_, weight_queue_2__0__7_,
         weight_queue_2__0__6_, weight_queue_2__0__5_, weight_queue_2__0__4_,
         weight_queue_2__0__3_, weight_queue_2__0__2_, weight_queue_2__0__1_,
         weight_queue_2__0__0_, weight_queue_2__1__7_, weight_queue_2__1__6_,
         weight_queue_2__1__5_, weight_queue_2__1__4_, weight_queue_2__1__3_,
         weight_queue_2__1__2_, weight_queue_2__1__1_, weight_queue_2__1__0_,
         weight_queue_2__2__7_, weight_queue_2__2__6_, weight_queue_2__2__5_,
         weight_queue_2__2__4_, weight_queue_2__2__3_, weight_queue_2__2__2_,
         weight_queue_2__2__1_, weight_queue_2__2__0_, weight_queue_2__3__7_,
         weight_queue_2__3__6_, weight_queue_2__3__5_, weight_queue_2__3__4_,
         weight_queue_2__3__3_, weight_queue_2__3__2_, weight_queue_2__3__1_,
         weight_queue_2__3__0_, weight_queue_2__4__7_, weight_queue_2__4__6_,
         weight_queue_2__4__5_, weight_queue_2__4__4_, weight_queue_2__4__3_,
         weight_queue_2__4__2_, weight_queue_2__4__1_, weight_queue_2__4__0_,
         weight_queue_2__5__7_, weight_queue_2__5__6_, weight_queue_2__5__5_,
         weight_queue_2__5__4_, weight_queue_2__5__3_, weight_queue_2__5__2_,
         weight_queue_2__5__1_, weight_queue_2__5__0_, weight_queue_2__6__7_,
         weight_queue_2__6__6_, weight_queue_2__6__5_, weight_queue_2__6__4_,
         weight_queue_2__6__3_, weight_queue_2__6__2_, weight_queue_2__6__1_,
         weight_queue_2__6__0_, weight_queue_2__7__7_, weight_queue_2__7__6_,
         weight_queue_2__7__5_, weight_queue_2__7__4_, weight_queue_2__7__3_,
         weight_queue_2__7__2_, weight_queue_2__7__1_, weight_queue_2__7__0_,
         weight_queue_3__0__7_, weight_queue_3__0__6_, weight_queue_3__0__5_,
         weight_queue_3__0__4_, weight_queue_3__0__3_, weight_queue_3__0__2_,
         weight_queue_3__0__1_, weight_queue_3__0__0_, weight_queue_3__1__7_,
         weight_queue_3__1__6_, weight_queue_3__1__5_, weight_queue_3__1__4_,
         weight_queue_3__1__3_, weight_queue_3__1__2_, weight_queue_3__1__1_,
         weight_queue_3__1__0_, weight_queue_3__2__7_, weight_queue_3__2__6_,
         weight_queue_3__2__5_, weight_queue_3__2__4_, weight_queue_3__2__3_,
         weight_queue_3__2__2_, weight_queue_3__2__1_, weight_queue_3__2__0_,
         weight_queue_3__3__7_, weight_queue_3__3__6_, weight_queue_3__3__5_,
         weight_queue_3__3__4_, weight_queue_3__3__3_, weight_queue_3__3__2_,
         weight_queue_3__3__1_, weight_queue_3__3__0_, weight_queue_3__4__7_,
         weight_queue_3__4__6_, weight_queue_3__4__5_, weight_queue_3__4__4_,
         weight_queue_3__4__3_, weight_queue_3__4__2_, weight_queue_3__4__1_,
         weight_queue_3__4__0_, weight_queue_3__5__7_, weight_queue_3__5__6_,
         weight_queue_3__5__5_, weight_queue_3__5__4_, weight_queue_3__5__3_,
         weight_queue_3__5__2_, weight_queue_3__5__1_, weight_queue_3__5__0_,
         weight_queue_3__6__7_, weight_queue_3__6__6_, weight_queue_3__6__5_,
         weight_queue_3__6__4_, weight_queue_3__6__3_, weight_queue_3__6__2_,
         weight_queue_3__6__1_, weight_queue_3__6__0_, weight_queue_3__7__7_,
         weight_queue_3__7__6_, weight_queue_3__7__5_, weight_queue_3__7__4_,
         weight_queue_3__7__3_, weight_queue_3__7__2_, weight_queue_3__7__1_,
         weight_queue_3__7__0_, weight_queue_4__0__7_, weight_queue_4__0__6_,
         weight_queue_4__0__5_, weight_queue_4__0__4_, weight_queue_4__0__3_,
         weight_queue_4__0__2_, weight_queue_4__0__1_, weight_queue_4__0__0_,
         weight_queue_4__1__7_, weight_queue_4__1__6_, weight_queue_4__1__5_,
         weight_queue_4__1__4_, weight_queue_4__1__3_, weight_queue_4__1__2_,
         weight_queue_4__1__1_, weight_queue_4__1__0_, weight_queue_4__2__7_,
         weight_queue_4__2__6_, weight_queue_4__2__5_, weight_queue_4__2__4_,
         weight_queue_4__2__3_, weight_queue_4__2__2_, weight_queue_4__2__1_,
         weight_queue_4__2__0_, weight_queue_4__3__7_, weight_queue_4__3__6_,
         weight_queue_4__3__5_, weight_queue_4__3__4_, weight_queue_4__3__3_,
         weight_queue_4__3__2_, weight_queue_4__3__1_, weight_queue_4__3__0_,
         weight_queue_4__4__7_, weight_queue_4__4__6_, weight_queue_4__4__5_,
         weight_queue_4__4__4_, weight_queue_4__4__3_, weight_queue_4__4__2_,
         weight_queue_4__4__1_, weight_queue_4__4__0_, weight_queue_4__5__7_,
         weight_queue_4__5__6_, weight_queue_4__5__5_, weight_queue_4__5__4_,
         weight_queue_4__5__3_, weight_queue_4__5__2_, weight_queue_4__5__1_,
         weight_queue_4__5__0_, weight_queue_4__6__7_, weight_queue_4__6__6_,
         weight_queue_4__6__5_, weight_queue_4__6__4_, weight_queue_4__6__3_,
         weight_queue_4__6__2_, weight_queue_4__6__1_, weight_queue_4__6__0_,
         weight_queue_4__7__7_, weight_queue_4__7__6_, weight_queue_4__7__5_,
         weight_queue_4__7__4_, weight_queue_4__7__3_, weight_queue_4__7__2_,
         weight_queue_4__7__1_, weight_queue_4__7__0_, weight_queue_5__0__7_,
         weight_queue_5__0__6_, weight_queue_5__0__5_, weight_queue_5__0__4_,
         weight_queue_5__0__3_, weight_queue_5__0__2_, weight_queue_5__0__1_,
         weight_queue_5__0__0_, weight_queue_5__1__7_, weight_queue_5__1__6_,
         weight_queue_5__1__5_, weight_queue_5__1__4_, weight_queue_5__1__3_,
         weight_queue_5__1__2_, weight_queue_5__1__1_, weight_queue_5__1__0_,
         weight_queue_5__2__7_, weight_queue_5__2__6_, weight_queue_5__2__5_,
         weight_queue_5__2__4_, weight_queue_5__2__3_, weight_queue_5__2__2_,
         weight_queue_5__2__1_, weight_queue_5__2__0_, weight_queue_5__3__7_,
         weight_queue_5__3__6_, weight_queue_5__3__5_, weight_queue_5__3__4_,
         weight_queue_5__3__3_, weight_queue_5__3__2_, weight_queue_5__3__1_,
         weight_queue_5__3__0_, weight_queue_5__4__7_, weight_queue_5__4__6_,
         weight_queue_5__4__5_, weight_queue_5__4__4_, weight_queue_5__4__3_,
         weight_queue_5__4__2_, weight_queue_5__4__1_, weight_queue_5__4__0_,
         weight_queue_5__5__7_, weight_queue_5__5__6_, weight_queue_5__5__5_,
         weight_queue_5__5__4_, weight_queue_5__5__3_, weight_queue_5__5__2_,
         weight_queue_5__5__1_, weight_queue_5__5__0_, weight_queue_5__6__7_,
         weight_queue_5__6__6_, weight_queue_5__6__5_, weight_queue_5__6__4_,
         weight_queue_5__6__3_, weight_queue_5__6__2_, weight_queue_5__6__1_,
         weight_queue_5__6__0_, weight_queue_5__7__7_, weight_queue_5__7__6_,
         weight_queue_5__7__5_, weight_queue_5__7__4_, weight_queue_5__7__3_,
         weight_queue_5__7__2_, weight_queue_5__7__1_, weight_queue_5__7__0_,
         weight_queue_6__0__7_, weight_queue_6__0__6_, weight_queue_6__0__5_,
         weight_queue_6__0__4_, weight_queue_6__0__3_, weight_queue_6__0__2_,
         weight_queue_6__0__1_, weight_queue_6__0__0_, weight_queue_6__1__7_,
         weight_queue_6__1__6_, weight_queue_6__1__5_, weight_queue_6__1__4_,
         weight_queue_6__1__3_, weight_queue_6__1__2_, weight_queue_6__1__1_,
         weight_queue_6__1__0_, weight_queue_6__2__7_, weight_queue_6__2__6_,
         weight_queue_6__2__5_, weight_queue_6__2__4_, weight_queue_6__2__3_,
         weight_queue_6__2__2_, weight_queue_6__2__1_, weight_queue_6__2__0_,
         weight_queue_6__3__7_, weight_queue_6__3__6_, weight_queue_6__3__5_,
         weight_queue_6__3__4_, weight_queue_6__3__3_, weight_queue_6__3__2_,
         weight_queue_6__3__1_, weight_queue_6__3__0_, weight_queue_6__4__7_,
         weight_queue_6__4__6_, weight_queue_6__4__5_, weight_queue_6__4__4_,
         weight_queue_6__4__3_, weight_queue_6__4__2_, weight_queue_6__4__1_,
         weight_queue_6__4__0_, weight_queue_6__5__7_, weight_queue_6__5__6_,
         weight_queue_6__5__5_, weight_queue_6__5__4_, weight_queue_6__5__3_,
         weight_queue_6__5__2_, weight_queue_6__5__1_, weight_queue_6__5__0_,
         weight_queue_6__6__7_, weight_queue_6__6__6_, weight_queue_6__6__5_,
         weight_queue_6__6__4_, weight_queue_6__6__3_, weight_queue_6__6__2_,
         weight_queue_6__6__1_, weight_queue_6__6__0_, weight_queue_6__7__7_,
         weight_queue_6__7__6_, weight_queue_6__7__5_, weight_queue_6__7__4_,
         weight_queue_6__7__3_, weight_queue_6__7__2_, weight_queue_6__7__1_,
         weight_queue_6__7__0_, weight_queue_7__0__7_, weight_queue_7__0__6_,
         weight_queue_7__0__5_, weight_queue_7__0__4_, weight_queue_7__0__3_,
         weight_queue_7__0__2_, weight_queue_7__0__1_, weight_queue_7__0__0_,
         weight_queue_7__1__7_, weight_queue_7__1__6_, weight_queue_7__1__5_,
         weight_queue_7__1__4_, weight_queue_7__1__3_, weight_queue_7__1__2_,
         weight_queue_7__1__1_, weight_queue_7__1__0_, weight_queue_7__2__7_,
         weight_queue_7__2__6_, weight_queue_7__2__5_, weight_queue_7__2__4_,
         weight_queue_7__2__3_, weight_queue_7__2__2_, weight_queue_7__2__1_,
         weight_queue_7__2__0_, weight_queue_7__3__7_, weight_queue_7__3__6_,
         weight_queue_7__3__5_, weight_queue_7__3__4_, weight_queue_7__3__3_,
         weight_queue_7__3__2_, weight_queue_7__3__1_, weight_queue_7__3__0_,
         weight_queue_7__4__7_, weight_queue_7__4__6_, weight_queue_7__4__5_,
         weight_queue_7__4__4_, weight_queue_7__4__3_, weight_queue_7__4__2_,
         weight_queue_7__4__1_, weight_queue_7__4__0_, weight_queue_7__5__7_,
         weight_queue_7__5__6_, weight_queue_7__5__5_, weight_queue_7__5__4_,
         weight_queue_7__5__3_, weight_queue_7__5__2_, weight_queue_7__5__1_,
         weight_queue_7__5__0_, weight_queue_7__6__7_, weight_queue_7__6__6_,
         weight_queue_7__6__5_, weight_queue_7__6__4_, weight_queue_7__6__3_,
         weight_queue_7__6__2_, weight_queue_7__6__1_, weight_queue_7__6__0_,
         weight_queue_7__7__7_, weight_queue_7__7__6_, weight_queue_7__7__5_,
         weight_queue_7__7__4_, weight_queue_7__7__3_, weight_queue_7__7__2_,
         weight_queue_7__7__1_, weight_queue_7__7__0_, data_queue_0__0__7_,
         data_queue_0__0__6_, data_queue_0__0__5_, data_queue_0__0__4_,
         data_queue_0__0__3_, data_queue_0__0__2_, data_queue_0__0__1_,
         data_queue_0__0__0_, data_queue_0__1__7_, data_queue_0__1__6_,
         data_queue_0__1__5_, data_queue_0__1__4_, data_queue_0__1__3_,
         data_queue_0__1__2_, data_queue_0__1__1_, data_queue_0__1__0_,
         data_queue_0__2__7_, data_queue_0__2__6_, data_queue_0__2__5_,
         data_queue_0__2__4_, data_queue_0__2__3_, data_queue_0__2__2_,
         data_queue_0__2__1_, data_queue_0__2__0_, data_queue_0__3__7_,
         data_queue_0__3__6_, data_queue_0__3__5_, data_queue_0__3__4_,
         data_queue_0__3__3_, data_queue_0__3__2_, data_queue_0__3__1_,
         data_queue_0__3__0_, data_queue_0__4__7_, data_queue_0__4__6_,
         data_queue_0__4__5_, data_queue_0__4__4_, data_queue_0__4__3_,
         data_queue_0__4__2_, data_queue_0__4__1_, data_queue_0__4__0_,
         data_queue_0__5__7_, data_queue_0__5__6_, data_queue_0__5__5_,
         data_queue_0__5__4_, data_queue_0__5__3_, data_queue_0__5__2_,
         data_queue_0__5__1_, data_queue_0__5__0_, data_queue_0__6__7_,
         data_queue_0__6__6_, data_queue_0__6__5_, data_queue_0__6__4_,
         data_queue_0__6__3_, data_queue_0__6__2_, data_queue_0__6__1_,
         data_queue_0__6__0_, data_queue_0__7__7_, data_queue_0__7__6_,
         data_queue_0__7__5_, data_queue_0__7__4_, data_queue_0__7__3_,
         data_queue_0__7__2_, data_queue_0__7__1_, data_queue_0__7__0_,
         data_queue_1__0__7_, data_queue_1__0__6_, data_queue_1__0__5_,
         data_queue_1__0__4_, data_queue_1__0__3_, data_queue_1__0__2_,
         data_queue_1__0__1_, data_queue_1__0__0_, data_queue_1__1__7_,
         data_queue_1__1__6_, data_queue_1__1__5_, data_queue_1__1__4_,
         data_queue_1__1__3_, data_queue_1__1__2_, data_queue_1__1__1_,
         data_queue_1__1__0_, data_queue_1__2__7_, data_queue_1__2__6_,
         data_queue_1__2__5_, data_queue_1__2__4_, data_queue_1__2__3_,
         data_queue_1__2__2_, data_queue_1__2__1_, data_queue_1__2__0_,
         data_queue_1__3__7_, data_queue_1__3__6_, data_queue_1__3__5_,
         data_queue_1__3__4_, data_queue_1__3__3_, data_queue_1__3__2_,
         data_queue_1__3__1_, data_queue_1__3__0_, data_queue_1__4__7_,
         data_queue_1__4__6_, data_queue_1__4__5_, data_queue_1__4__4_,
         data_queue_1__4__3_, data_queue_1__4__2_, data_queue_1__4__1_,
         data_queue_1__4__0_, data_queue_1__5__7_, data_queue_1__5__6_,
         data_queue_1__5__5_, data_queue_1__5__4_, data_queue_1__5__3_,
         data_queue_1__5__2_, data_queue_1__5__1_, data_queue_1__5__0_,
         data_queue_1__6__7_, data_queue_1__6__6_, data_queue_1__6__5_,
         data_queue_1__6__4_, data_queue_1__6__3_, data_queue_1__6__2_,
         data_queue_1__6__1_, data_queue_1__6__0_, data_queue_1__7__7_,
         data_queue_1__7__6_, data_queue_1__7__5_, data_queue_1__7__4_,
         data_queue_1__7__3_, data_queue_1__7__2_, data_queue_1__7__1_,
         data_queue_1__7__0_, data_queue_2__0__7_, data_queue_2__0__6_,
         data_queue_2__0__5_, data_queue_2__0__4_, data_queue_2__0__3_,
         data_queue_2__0__2_, data_queue_2__0__1_, data_queue_2__0__0_,
         data_queue_2__1__7_, data_queue_2__1__6_, data_queue_2__1__5_,
         data_queue_2__1__4_, data_queue_2__1__3_, data_queue_2__1__2_,
         data_queue_2__1__1_, data_queue_2__1__0_, data_queue_2__2__7_,
         data_queue_2__2__6_, data_queue_2__2__5_, data_queue_2__2__4_,
         data_queue_2__2__3_, data_queue_2__2__2_, data_queue_2__2__1_,
         data_queue_2__2__0_, data_queue_2__3__7_, data_queue_2__3__6_,
         data_queue_2__3__5_, data_queue_2__3__4_, data_queue_2__3__3_,
         data_queue_2__3__2_, data_queue_2__3__1_, data_queue_2__3__0_,
         data_queue_2__4__7_, data_queue_2__4__6_, data_queue_2__4__5_,
         data_queue_2__4__4_, data_queue_2__4__3_, data_queue_2__4__2_,
         data_queue_2__4__1_, data_queue_2__4__0_, data_queue_2__5__7_,
         data_queue_2__5__6_, data_queue_2__5__5_, data_queue_2__5__4_,
         data_queue_2__5__3_, data_queue_2__5__2_, data_queue_2__5__1_,
         data_queue_2__5__0_, data_queue_2__6__7_, data_queue_2__6__6_,
         data_queue_2__6__5_, data_queue_2__6__4_, data_queue_2__6__3_,
         data_queue_2__6__2_, data_queue_2__6__1_, data_queue_2__6__0_,
         data_queue_2__7__7_, data_queue_2__7__6_, data_queue_2__7__5_,
         data_queue_2__7__4_, data_queue_2__7__3_, data_queue_2__7__2_,
         data_queue_2__7__1_, data_queue_2__7__0_, data_queue_3__0__7_,
         data_queue_3__0__6_, data_queue_3__0__5_, data_queue_3__0__4_,
         data_queue_3__0__3_, data_queue_3__0__2_, data_queue_3__0__1_,
         data_queue_3__0__0_, data_queue_3__1__7_, data_queue_3__1__6_,
         data_queue_3__1__5_, data_queue_3__1__4_, data_queue_3__1__3_,
         data_queue_3__1__2_, data_queue_3__1__1_, data_queue_3__1__0_,
         data_queue_3__2__7_, data_queue_3__2__6_, data_queue_3__2__5_,
         data_queue_3__2__4_, data_queue_3__2__3_, data_queue_3__2__2_,
         data_queue_3__2__1_, data_queue_3__2__0_, data_queue_3__3__7_,
         data_queue_3__3__6_, data_queue_3__3__5_, data_queue_3__3__4_,
         data_queue_3__3__3_, data_queue_3__3__2_, data_queue_3__3__1_,
         data_queue_3__3__0_, data_queue_3__4__7_, data_queue_3__4__6_,
         data_queue_3__4__5_, data_queue_3__4__4_, data_queue_3__4__3_,
         data_queue_3__4__2_, data_queue_3__4__1_, data_queue_3__4__0_,
         data_queue_3__5__7_, data_queue_3__5__6_, data_queue_3__5__5_,
         data_queue_3__5__4_, data_queue_3__5__3_, data_queue_3__5__2_,
         data_queue_3__5__1_, data_queue_3__5__0_, data_queue_3__6__7_,
         data_queue_3__6__6_, data_queue_3__6__5_, data_queue_3__6__4_,
         data_queue_3__6__3_, data_queue_3__6__2_, data_queue_3__6__1_,
         data_queue_3__6__0_, data_queue_3__7__7_, data_queue_3__7__6_,
         data_queue_3__7__5_, data_queue_3__7__4_, data_queue_3__7__3_,
         data_queue_3__7__2_, data_queue_3__7__1_, data_queue_3__7__0_,
         data_queue_4__0__7_, data_queue_4__0__6_, data_queue_4__0__5_,
         data_queue_4__0__4_, data_queue_4__0__3_, data_queue_4__0__2_,
         data_queue_4__0__1_, data_queue_4__0__0_, data_queue_4__1__7_,
         data_queue_4__1__6_, data_queue_4__1__5_, data_queue_4__1__4_,
         data_queue_4__1__3_, data_queue_4__1__2_, data_queue_4__1__1_,
         data_queue_4__1__0_, data_queue_4__2__7_, data_queue_4__2__6_,
         data_queue_4__2__5_, data_queue_4__2__4_, data_queue_4__2__3_,
         data_queue_4__2__2_, data_queue_4__2__1_, data_queue_4__2__0_,
         data_queue_4__3__7_, data_queue_4__3__6_, data_queue_4__3__5_,
         data_queue_4__3__4_, data_queue_4__3__3_, data_queue_4__3__2_,
         data_queue_4__3__1_, data_queue_4__3__0_, data_queue_4__4__7_,
         data_queue_4__4__6_, data_queue_4__4__5_, data_queue_4__4__4_,
         data_queue_4__4__3_, data_queue_4__4__2_, data_queue_4__4__1_,
         data_queue_4__4__0_, data_queue_4__5__7_, data_queue_4__5__6_,
         data_queue_4__5__5_, data_queue_4__5__4_, data_queue_4__5__3_,
         data_queue_4__5__2_, data_queue_4__5__1_, data_queue_4__5__0_,
         data_queue_4__6__7_, data_queue_4__6__6_, data_queue_4__6__5_,
         data_queue_4__6__4_, data_queue_4__6__3_, data_queue_4__6__2_,
         data_queue_4__6__1_, data_queue_4__6__0_, data_queue_4__7__7_,
         data_queue_4__7__6_, data_queue_4__7__5_, data_queue_4__7__4_,
         data_queue_4__7__3_, data_queue_4__7__2_, data_queue_4__7__1_,
         data_queue_4__7__0_, data_queue_5__0__7_, data_queue_5__0__6_,
         data_queue_5__0__5_, data_queue_5__0__4_, data_queue_5__0__3_,
         data_queue_5__0__2_, data_queue_5__0__1_, data_queue_5__0__0_,
         data_queue_5__1__7_, data_queue_5__1__6_, data_queue_5__1__5_,
         data_queue_5__1__4_, data_queue_5__1__3_, data_queue_5__1__2_,
         data_queue_5__1__1_, data_queue_5__1__0_, data_queue_5__2__7_,
         data_queue_5__2__6_, data_queue_5__2__5_, data_queue_5__2__4_,
         data_queue_5__2__3_, data_queue_5__2__2_, data_queue_5__2__1_,
         data_queue_5__2__0_, data_queue_5__3__7_, data_queue_5__3__6_,
         data_queue_5__3__5_, data_queue_5__3__4_, data_queue_5__3__3_,
         data_queue_5__3__2_, data_queue_5__3__1_, data_queue_5__3__0_,
         data_queue_5__4__7_, data_queue_5__4__6_, data_queue_5__4__5_,
         data_queue_5__4__4_, data_queue_5__4__3_, data_queue_5__4__2_,
         data_queue_5__4__1_, data_queue_5__4__0_, data_queue_5__5__7_,
         data_queue_5__5__6_, data_queue_5__5__5_, data_queue_5__5__4_,
         data_queue_5__5__3_, data_queue_5__5__2_, data_queue_5__5__1_,
         data_queue_5__5__0_, data_queue_5__6__7_, data_queue_5__6__6_,
         data_queue_5__6__5_, data_queue_5__6__4_, data_queue_5__6__3_,
         data_queue_5__6__2_, data_queue_5__6__1_, data_queue_5__6__0_,
         data_queue_5__7__7_, data_queue_5__7__6_, data_queue_5__7__5_,
         data_queue_5__7__4_, data_queue_5__7__3_, data_queue_5__7__2_,
         data_queue_5__7__1_, data_queue_5__7__0_, data_queue_6__0__7_,
         data_queue_6__0__6_, data_queue_6__0__5_, data_queue_6__0__4_,
         data_queue_6__0__3_, data_queue_6__0__2_, data_queue_6__0__1_,
         data_queue_6__0__0_, data_queue_6__1__7_, data_queue_6__1__6_,
         data_queue_6__1__5_, data_queue_6__1__4_, data_queue_6__1__3_,
         data_queue_6__1__2_, data_queue_6__1__1_, data_queue_6__1__0_,
         data_queue_6__2__7_, data_queue_6__2__6_, data_queue_6__2__5_,
         data_queue_6__2__4_, data_queue_6__2__3_, data_queue_6__2__2_,
         data_queue_6__2__1_, data_queue_6__2__0_, data_queue_6__3__7_,
         data_queue_6__3__6_, data_queue_6__3__5_, data_queue_6__3__4_,
         data_queue_6__3__3_, data_queue_6__3__2_, data_queue_6__3__1_,
         data_queue_6__3__0_, data_queue_6__4__7_, data_queue_6__4__6_,
         data_queue_6__4__5_, data_queue_6__4__4_, data_queue_6__4__3_,
         data_queue_6__4__2_, data_queue_6__4__1_, data_queue_6__4__0_,
         data_queue_6__5__7_, data_queue_6__5__6_, data_queue_6__5__5_,
         data_queue_6__5__4_, data_queue_6__5__3_, data_queue_6__5__2_,
         data_queue_6__5__1_, data_queue_6__5__0_, data_queue_6__6__7_,
         data_queue_6__6__6_, data_queue_6__6__5_, data_queue_6__6__4_,
         data_queue_6__6__3_, data_queue_6__6__2_, data_queue_6__6__1_,
         data_queue_6__6__0_, data_queue_6__7__7_, data_queue_6__7__6_,
         data_queue_6__7__5_, data_queue_6__7__4_, data_queue_6__7__3_,
         data_queue_6__7__2_, data_queue_6__7__1_, data_queue_6__7__0_,
         data_queue_7__0__7_, data_queue_7__0__6_, data_queue_7__0__5_,
         data_queue_7__0__4_, data_queue_7__0__3_, data_queue_7__0__2_,
         data_queue_7__0__1_, data_queue_7__0__0_, data_queue_7__1__7_,
         data_queue_7__1__6_, data_queue_7__1__5_, data_queue_7__1__4_,
         data_queue_7__1__3_, data_queue_7__1__2_, data_queue_7__1__1_,
         data_queue_7__1__0_, data_queue_7__2__7_, data_queue_7__2__6_,
         data_queue_7__2__5_, data_queue_7__2__4_, data_queue_7__2__3_,
         data_queue_7__2__2_, data_queue_7__2__1_, data_queue_7__2__0_,
         data_queue_7__3__7_, data_queue_7__3__6_, data_queue_7__3__5_,
         data_queue_7__3__4_, data_queue_7__3__3_, data_queue_7__3__2_,
         data_queue_7__3__1_, data_queue_7__3__0_, data_queue_7__4__7_,
         data_queue_7__4__6_, data_queue_7__4__5_, data_queue_7__4__4_,
         data_queue_7__4__3_, data_queue_7__4__2_, data_queue_7__4__1_,
         data_queue_7__4__0_, data_queue_7__5__7_, data_queue_7__5__6_,
         data_queue_7__5__5_, data_queue_7__5__4_, data_queue_7__5__3_,
         data_queue_7__5__2_, data_queue_7__5__1_, data_queue_7__5__0_,
         data_queue_7__6__7_, data_queue_7__6__6_, data_queue_7__6__5_,
         data_queue_7__6__4_, data_queue_7__6__3_, data_queue_7__6__2_,
         data_queue_7__6__1_, data_queue_7__6__0_, data_queue_7__7__7_,
         data_queue_7__7__6_, data_queue_7__7__5_, data_queue_7__7__4_,
         data_queue_7__7__3_, data_queue_7__7__2_, data_queue_7__7__1_,
         data_queue_7__7__0_, matrix_mul_2D_0__0__20_, matrix_mul_2D_0__0__19_,
         matrix_mul_2D_0__0__18_, matrix_mul_2D_0__0__17_,
         matrix_mul_2D_0__0__16_, matrix_mul_2D_0__0__15_,
         matrix_mul_2D_0__0__14_, matrix_mul_2D_0__0__13_,
         matrix_mul_2D_0__0__12_, matrix_mul_2D_0__0__11_,
         matrix_mul_2D_0__0__10_, matrix_mul_2D_0__0__9_,
         matrix_mul_2D_0__0__8_, matrix_mul_2D_0__0__7_,
         matrix_mul_2D_0__0__6_, matrix_mul_2D_0__0__5_,
         matrix_mul_2D_0__0__4_, matrix_mul_2D_0__0__3_,
         matrix_mul_2D_0__0__2_, matrix_mul_2D_0__0__1_,
         matrix_mul_2D_0__0__0_, matrix_mul_2D_0__1__20_,
         matrix_mul_2D_0__1__19_, matrix_mul_2D_0__1__18_,
         matrix_mul_2D_0__1__17_, matrix_mul_2D_0__1__16_,
         matrix_mul_2D_0__1__15_, matrix_mul_2D_0__1__14_,
         matrix_mul_2D_0__1__13_, matrix_mul_2D_0__1__12_,
         matrix_mul_2D_0__1__11_, matrix_mul_2D_0__1__10_,
         matrix_mul_2D_0__1__9_, matrix_mul_2D_0__1__8_,
         matrix_mul_2D_0__1__7_, matrix_mul_2D_0__1__6_,
         matrix_mul_2D_0__1__5_, matrix_mul_2D_0__1__4_,
         matrix_mul_2D_0__1__3_, matrix_mul_2D_0__1__2_,
         matrix_mul_2D_0__1__1_, matrix_mul_2D_0__1__0_,
         matrix_mul_2D_0__2__20_, matrix_mul_2D_0__2__19_,
         matrix_mul_2D_0__2__18_, matrix_mul_2D_0__2__17_,
         matrix_mul_2D_0__2__16_, matrix_mul_2D_0__2__15_,
         matrix_mul_2D_0__2__14_, matrix_mul_2D_0__2__13_,
         matrix_mul_2D_0__2__12_, matrix_mul_2D_0__2__11_,
         matrix_mul_2D_0__2__10_, matrix_mul_2D_0__2__9_,
         matrix_mul_2D_0__2__8_, matrix_mul_2D_0__2__7_,
         matrix_mul_2D_0__2__6_, matrix_mul_2D_0__2__5_,
         matrix_mul_2D_0__2__4_, matrix_mul_2D_0__2__3_,
         matrix_mul_2D_0__2__2_, matrix_mul_2D_0__2__1_,
         matrix_mul_2D_0__2__0_, matrix_mul_2D_0__3__20_,
         matrix_mul_2D_0__3__19_, matrix_mul_2D_0__3__18_,
         matrix_mul_2D_0__3__17_, matrix_mul_2D_0__3__16_,
         matrix_mul_2D_0__3__15_, matrix_mul_2D_0__3__14_,
         matrix_mul_2D_0__3__13_, matrix_mul_2D_0__3__12_,
         matrix_mul_2D_0__3__11_, matrix_mul_2D_0__3__10_,
         matrix_mul_2D_0__3__9_, matrix_mul_2D_0__3__8_,
         matrix_mul_2D_0__3__7_, matrix_mul_2D_0__3__6_,
         matrix_mul_2D_0__3__5_, matrix_mul_2D_0__3__4_,
         matrix_mul_2D_0__3__3_, matrix_mul_2D_0__3__2_,
         matrix_mul_2D_0__3__1_, matrix_mul_2D_0__3__0_,
         matrix_mul_2D_0__4__20_, matrix_mul_2D_0__4__19_,
         matrix_mul_2D_0__4__18_, matrix_mul_2D_0__4__17_,
         matrix_mul_2D_0__4__16_, matrix_mul_2D_0__4__15_,
         matrix_mul_2D_0__4__14_, matrix_mul_2D_0__4__13_,
         matrix_mul_2D_0__4__12_, matrix_mul_2D_0__4__11_,
         matrix_mul_2D_0__4__10_, matrix_mul_2D_0__4__9_,
         matrix_mul_2D_0__4__8_, matrix_mul_2D_0__4__7_,
         matrix_mul_2D_0__4__6_, matrix_mul_2D_0__4__5_,
         matrix_mul_2D_0__4__4_, matrix_mul_2D_0__4__3_,
         matrix_mul_2D_0__4__2_, matrix_mul_2D_0__4__1_,
         matrix_mul_2D_0__4__0_, matrix_mul_2D_0__5__20_,
         matrix_mul_2D_0__5__19_, matrix_mul_2D_0__5__18_,
         matrix_mul_2D_0__5__17_, matrix_mul_2D_0__5__16_,
         matrix_mul_2D_0__5__15_, matrix_mul_2D_0__5__14_,
         matrix_mul_2D_0__5__13_, matrix_mul_2D_0__5__12_,
         matrix_mul_2D_0__5__11_, matrix_mul_2D_0__5__10_,
         matrix_mul_2D_0__5__9_, matrix_mul_2D_0__5__8_,
         matrix_mul_2D_0__5__7_, matrix_mul_2D_0__5__6_,
         matrix_mul_2D_0__5__5_, matrix_mul_2D_0__5__4_,
         matrix_mul_2D_0__5__3_, matrix_mul_2D_0__5__2_,
         matrix_mul_2D_0__5__1_, matrix_mul_2D_0__5__0_,
         matrix_mul_2D_0__6__20_, matrix_mul_2D_0__6__19_,
         matrix_mul_2D_0__6__18_, matrix_mul_2D_0__6__17_,
         matrix_mul_2D_0__6__16_, matrix_mul_2D_0__6__15_,
         matrix_mul_2D_0__6__14_, matrix_mul_2D_0__6__13_,
         matrix_mul_2D_0__6__12_, matrix_mul_2D_0__6__11_,
         matrix_mul_2D_0__6__10_, matrix_mul_2D_0__6__9_,
         matrix_mul_2D_0__6__8_, matrix_mul_2D_0__6__7_,
         matrix_mul_2D_0__6__6_, matrix_mul_2D_0__6__5_,
         matrix_mul_2D_0__6__4_, matrix_mul_2D_0__6__3_,
         matrix_mul_2D_0__6__2_, matrix_mul_2D_0__6__1_,
         matrix_mul_2D_0__6__0_, matrix_mul_2D_0__7__20_,
         matrix_mul_2D_0__7__19_, matrix_mul_2D_0__7__18_,
         matrix_mul_2D_0__7__17_, matrix_mul_2D_0__7__16_,
         matrix_mul_2D_0__7__15_, matrix_mul_2D_0__7__14_,
         matrix_mul_2D_0__7__13_, matrix_mul_2D_0__7__12_,
         matrix_mul_2D_0__7__11_, matrix_mul_2D_0__7__10_,
         matrix_mul_2D_0__7__9_, matrix_mul_2D_0__7__8_,
         matrix_mul_2D_0__7__7_, matrix_mul_2D_0__7__6_,
         matrix_mul_2D_0__7__5_, matrix_mul_2D_0__7__4_,
         matrix_mul_2D_0__7__3_, matrix_mul_2D_0__7__2_,
         matrix_mul_2D_0__7__1_, matrix_mul_2D_0__7__0_,
         matrix_mul_2D_1__0__20_, matrix_mul_2D_1__0__19_,
         matrix_mul_2D_1__0__18_, matrix_mul_2D_1__0__17_,
         matrix_mul_2D_1__0__16_, matrix_mul_2D_1__0__15_,
         matrix_mul_2D_1__0__14_, matrix_mul_2D_1__0__13_,
         matrix_mul_2D_1__0__12_, matrix_mul_2D_1__0__11_,
         matrix_mul_2D_1__0__10_, matrix_mul_2D_1__0__9_,
         matrix_mul_2D_1__0__8_, matrix_mul_2D_1__0__7_,
         matrix_mul_2D_1__0__6_, matrix_mul_2D_1__0__5_,
         matrix_mul_2D_1__0__4_, matrix_mul_2D_1__0__3_,
         matrix_mul_2D_1__0__2_, matrix_mul_2D_1__0__1_,
         matrix_mul_2D_1__0__0_, matrix_mul_2D_1__1__20_,
         matrix_mul_2D_1__1__19_, matrix_mul_2D_1__1__18_,
         matrix_mul_2D_1__1__17_, matrix_mul_2D_1__1__16_,
         matrix_mul_2D_1__1__15_, matrix_mul_2D_1__1__14_,
         matrix_mul_2D_1__1__13_, matrix_mul_2D_1__1__12_,
         matrix_mul_2D_1__1__11_, matrix_mul_2D_1__1__10_,
         matrix_mul_2D_1__1__9_, matrix_mul_2D_1__1__8_,
         matrix_mul_2D_1__1__7_, matrix_mul_2D_1__1__6_,
         matrix_mul_2D_1__1__5_, matrix_mul_2D_1__1__4_,
         matrix_mul_2D_1__1__3_, matrix_mul_2D_1__1__2_,
         matrix_mul_2D_1__1__1_, matrix_mul_2D_1__1__0_,
         matrix_mul_2D_1__2__20_, matrix_mul_2D_1__2__19_,
         matrix_mul_2D_1__2__18_, matrix_mul_2D_1__2__17_,
         matrix_mul_2D_1__2__16_, matrix_mul_2D_1__2__15_,
         matrix_mul_2D_1__2__14_, matrix_mul_2D_1__2__13_,
         matrix_mul_2D_1__2__12_, matrix_mul_2D_1__2__11_,
         matrix_mul_2D_1__2__10_, matrix_mul_2D_1__2__9_,
         matrix_mul_2D_1__2__8_, matrix_mul_2D_1__2__7_,
         matrix_mul_2D_1__2__6_, matrix_mul_2D_1__2__5_,
         matrix_mul_2D_1__2__4_, matrix_mul_2D_1__2__3_,
         matrix_mul_2D_1__2__2_, matrix_mul_2D_1__2__1_,
         matrix_mul_2D_1__2__0_, matrix_mul_2D_1__3__20_,
         matrix_mul_2D_1__3__19_, matrix_mul_2D_1__3__18_,
         matrix_mul_2D_1__3__17_, matrix_mul_2D_1__3__16_,
         matrix_mul_2D_1__3__15_, matrix_mul_2D_1__3__14_,
         matrix_mul_2D_1__3__13_, matrix_mul_2D_1__3__12_,
         matrix_mul_2D_1__3__11_, matrix_mul_2D_1__3__10_,
         matrix_mul_2D_1__3__9_, matrix_mul_2D_1__3__8_,
         matrix_mul_2D_1__3__7_, matrix_mul_2D_1__3__6_,
         matrix_mul_2D_1__3__5_, matrix_mul_2D_1__3__4_,
         matrix_mul_2D_1__3__3_, matrix_mul_2D_1__3__2_,
         matrix_mul_2D_1__3__1_, matrix_mul_2D_1__3__0_,
         matrix_mul_2D_1__4__20_, matrix_mul_2D_1__4__19_,
         matrix_mul_2D_1__4__18_, matrix_mul_2D_1__4__17_,
         matrix_mul_2D_1__4__16_, matrix_mul_2D_1__4__15_,
         matrix_mul_2D_1__4__14_, matrix_mul_2D_1__4__13_,
         matrix_mul_2D_1__4__12_, matrix_mul_2D_1__4__11_,
         matrix_mul_2D_1__4__10_, matrix_mul_2D_1__4__9_,
         matrix_mul_2D_1__4__8_, matrix_mul_2D_1__4__7_,
         matrix_mul_2D_1__4__6_, matrix_mul_2D_1__4__5_,
         matrix_mul_2D_1__4__4_, matrix_mul_2D_1__4__3_,
         matrix_mul_2D_1__4__2_, matrix_mul_2D_1__4__1_,
         matrix_mul_2D_1__4__0_, matrix_mul_2D_1__5__20_,
         matrix_mul_2D_1__5__19_, matrix_mul_2D_1__5__18_,
         matrix_mul_2D_1__5__17_, matrix_mul_2D_1__5__16_,
         matrix_mul_2D_1__5__15_, matrix_mul_2D_1__5__14_,
         matrix_mul_2D_1__5__13_, matrix_mul_2D_1__5__12_,
         matrix_mul_2D_1__5__11_, matrix_mul_2D_1__5__10_,
         matrix_mul_2D_1__5__9_, matrix_mul_2D_1__5__8_,
         matrix_mul_2D_1__5__7_, matrix_mul_2D_1__5__6_,
         matrix_mul_2D_1__5__5_, matrix_mul_2D_1__5__4_,
         matrix_mul_2D_1__5__3_, matrix_mul_2D_1__5__2_,
         matrix_mul_2D_1__5__1_, matrix_mul_2D_1__5__0_,
         matrix_mul_2D_1__6__20_, matrix_mul_2D_1__6__19_,
         matrix_mul_2D_1__6__18_, matrix_mul_2D_1__6__17_,
         matrix_mul_2D_1__6__16_, matrix_mul_2D_1__6__15_,
         matrix_mul_2D_1__6__14_, matrix_mul_2D_1__6__13_,
         matrix_mul_2D_1__6__12_, matrix_mul_2D_1__6__11_,
         matrix_mul_2D_1__6__10_, matrix_mul_2D_1__6__9_,
         matrix_mul_2D_1__6__8_, matrix_mul_2D_1__6__7_,
         matrix_mul_2D_1__6__6_, matrix_mul_2D_1__6__5_,
         matrix_mul_2D_1__6__4_, matrix_mul_2D_1__6__3_,
         matrix_mul_2D_1__6__2_, matrix_mul_2D_1__6__1_,
         matrix_mul_2D_1__6__0_, matrix_mul_2D_1__7__20_,
         matrix_mul_2D_1__7__19_, matrix_mul_2D_1__7__18_,
         matrix_mul_2D_1__7__17_, matrix_mul_2D_1__7__16_,
         matrix_mul_2D_1__7__15_, matrix_mul_2D_1__7__14_,
         matrix_mul_2D_1__7__13_, matrix_mul_2D_1__7__12_,
         matrix_mul_2D_1__7__11_, matrix_mul_2D_1__7__10_,
         matrix_mul_2D_1__7__9_, matrix_mul_2D_1__7__8_,
         matrix_mul_2D_1__7__7_, matrix_mul_2D_1__7__6_,
         matrix_mul_2D_1__7__5_, matrix_mul_2D_1__7__4_,
         matrix_mul_2D_1__7__3_, matrix_mul_2D_1__7__2_,
         matrix_mul_2D_1__7__1_, matrix_mul_2D_1__7__0_,
         matrix_mul_2D_2__0__20_, matrix_mul_2D_2__0__19_,
         matrix_mul_2D_2__0__18_, matrix_mul_2D_2__0__17_,
         matrix_mul_2D_2__0__16_, matrix_mul_2D_2__0__15_,
         matrix_mul_2D_2__0__14_, matrix_mul_2D_2__0__13_,
         matrix_mul_2D_2__0__12_, matrix_mul_2D_2__0__11_,
         matrix_mul_2D_2__0__10_, matrix_mul_2D_2__0__9_,
         matrix_mul_2D_2__0__8_, matrix_mul_2D_2__0__7_,
         matrix_mul_2D_2__0__6_, matrix_mul_2D_2__0__5_,
         matrix_mul_2D_2__0__4_, matrix_mul_2D_2__0__3_,
         matrix_mul_2D_2__0__2_, matrix_mul_2D_2__0__1_,
         matrix_mul_2D_2__0__0_, matrix_mul_2D_2__1__20_,
         matrix_mul_2D_2__1__19_, matrix_mul_2D_2__1__18_,
         matrix_mul_2D_2__1__17_, matrix_mul_2D_2__1__16_,
         matrix_mul_2D_2__1__15_, matrix_mul_2D_2__1__14_,
         matrix_mul_2D_2__1__13_, matrix_mul_2D_2__1__12_,
         matrix_mul_2D_2__1__11_, matrix_mul_2D_2__1__10_,
         matrix_mul_2D_2__1__9_, matrix_mul_2D_2__1__8_,
         matrix_mul_2D_2__1__7_, matrix_mul_2D_2__1__6_,
         matrix_mul_2D_2__1__5_, matrix_mul_2D_2__1__4_,
         matrix_mul_2D_2__1__3_, matrix_mul_2D_2__1__2_,
         matrix_mul_2D_2__1__1_, matrix_mul_2D_2__1__0_,
         matrix_mul_2D_2__2__20_, matrix_mul_2D_2__2__19_,
         matrix_mul_2D_2__2__18_, matrix_mul_2D_2__2__17_,
         matrix_mul_2D_2__2__16_, matrix_mul_2D_2__2__15_,
         matrix_mul_2D_2__2__14_, matrix_mul_2D_2__2__13_,
         matrix_mul_2D_2__2__12_, matrix_mul_2D_2__2__11_,
         matrix_mul_2D_2__2__10_, matrix_mul_2D_2__2__9_,
         matrix_mul_2D_2__2__8_, matrix_mul_2D_2__2__7_,
         matrix_mul_2D_2__2__6_, matrix_mul_2D_2__2__5_,
         matrix_mul_2D_2__2__4_, matrix_mul_2D_2__2__3_,
         matrix_mul_2D_2__2__2_, matrix_mul_2D_2__2__1_,
         matrix_mul_2D_2__2__0_, matrix_mul_2D_2__3__20_,
         matrix_mul_2D_2__3__19_, matrix_mul_2D_2__3__18_,
         matrix_mul_2D_2__3__17_, matrix_mul_2D_2__3__16_,
         matrix_mul_2D_2__3__15_, matrix_mul_2D_2__3__14_,
         matrix_mul_2D_2__3__13_, matrix_mul_2D_2__3__12_,
         matrix_mul_2D_2__3__11_, matrix_mul_2D_2__3__10_,
         matrix_mul_2D_2__3__9_, matrix_mul_2D_2__3__8_,
         matrix_mul_2D_2__3__7_, matrix_mul_2D_2__3__6_,
         matrix_mul_2D_2__3__5_, matrix_mul_2D_2__3__4_,
         matrix_mul_2D_2__3__3_, matrix_mul_2D_2__3__2_,
         matrix_mul_2D_2__3__1_, matrix_mul_2D_2__3__0_,
         matrix_mul_2D_2__4__20_, matrix_mul_2D_2__4__19_,
         matrix_mul_2D_2__4__18_, matrix_mul_2D_2__4__17_,
         matrix_mul_2D_2__4__16_, matrix_mul_2D_2__4__15_,
         matrix_mul_2D_2__4__14_, matrix_mul_2D_2__4__13_,
         matrix_mul_2D_2__4__12_, matrix_mul_2D_2__4__11_,
         matrix_mul_2D_2__4__10_, matrix_mul_2D_2__4__9_,
         matrix_mul_2D_2__4__8_, matrix_mul_2D_2__4__7_,
         matrix_mul_2D_2__4__6_, matrix_mul_2D_2__4__5_,
         matrix_mul_2D_2__4__4_, matrix_mul_2D_2__4__3_,
         matrix_mul_2D_2__4__2_, matrix_mul_2D_2__4__1_,
         matrix_mul_2D_2__4__0_, matrix_mul_2D_2__5__20_,
         matrix_mul_2D_2__5__19_, matrix_mul_2D_2__5__18_,
         matrix_mul_2D_2__5__17_, matrix_mul_2D_2__5__16_,
         matrix_mul_2D_2__5__15_, matrix_mul_2D_2__5__14_,
         matrix_mul_2D_2__5__13_, matrix_mul_2D_2__5__12_,
         matrix_mul_2D_2__5__11_, matrix_mul_2D_2__5__10_,
         matrix_mul_2D_2__5__9_, matrix_mul_2D_2__5__8_,
         matrix_mul_2D_2__5__7_, matrix_mul_2D_2__5__6_,
         matrix_mul_2D_2__5__5_, matrix_mul_2D_2__5__4_,
         matrix_mul_2D_2__5__3_, matrix_mul_2D_2__5__2_,
         matrix_mul_2D_2__5__1_, matrix_mul_2D_2__5__0_,
         matrix_mul_2D_2__6__20_, matrix_mul_2D_2__6__19_,
         matrix_mul_2D_2__6__18_, matrix_mul_2D_2__6__17_,
         matrix_mul_2D_2__6__16_, matrix_mul_2D_2__6__15_,
         matrix_mul_2D_2__6__14_, matrix_mul_2D_2__6__13_,
         matrix_mul_2D_2__6__12_, matrix_mul_2D_2__6__11_,
         matrix_mul_2D_2__6__10_, matrix_mul_2D_2__6__9_,
         matrix_mul_2D_2__6__8_, matrix_mul_2D_2__6__7_,
         matrix_mul_2D_2__6__6_, matrix_mul_2D_2__6__5_,
         matrix_mul_2D_2__6__4_, matrix_mul_2D_2__6__3_,
         matrix_mul_2D_2__6__2_, matrix_mul_2D_2__6__1_,
         matrix_mul_2D_2__6__0_, matrix_mul_2D_2__7__20_,
         matrix_mul_2D_2__7__19_, matrix_mul_2D_2__7__18_,
         matrix_mul_2D_2__7__17_, matrix_mul_2D_2__7__16_,
         matrix_mul_2D_2__7__15_, matrix_mul_2D_2__7__14_,
         matrix_mul_2D_2__7__13_, matrix_mul_2D_2__7__12_,
         matrix_mul_2D_2__7__11_, matrix_mul_2D_2__7__10_,
         matrix_mul_2D_2__7__9_, matrix_mul_2D_2__7__8_,
         matrix_mul_2D_2__7__7_, matrix_mul_2D_2__7__6_,
         matrix_mul_2D_2__7__5_, matrix_mul_2D_2__7__4_,
         matrix_mul_2D_2__7__3_, matrix_mul_2D_2__7__2_,
         matrix_mul_2D_2__7__1_, matrix_mul_2D_2__7__0_,
         matrix_mul_2D_3__0__20_, matrix_mul_2D_3__0__19_,
         matrix_mul_2D_3__0__18_, matrix_mul_2D_3__0__17_,
         matrix_mul_2D_3__0__16_, matrix_mul_2D_3__0__15_,
         matrix_mul_2D_3__0__14_, matrix_mul_2D_3__0__13_,
         matrix_mul_2D_3__0__12_, matrix_mul_2D_3__0__11_,
         matrix_mul_2D_3__0__10_, matrix_mul_2D_3__0__9_,
         matrix_mul_2D_3__0__8_, matrix_mul_2D_3__0__7_,
         matrix_mul_2D_3__0__6_, matrix_mul_2D_3__0__5_,
         matrix_mul_2D_3__0__4_, matrix_mul_2D_3__0__3_,
         matrix_mul_2D_3__0__2_, matrix_mul_2D_3__0__1_,
         matrix_mul_2D_3__0__0_, matrix_mul_2D_3__1__20_,
         matrix_mul_2D_3__1__19_, matrix_mul_2D_3__1__18_,
         matrix_mul_2D_3__1__17_, matrix_mul_2D_3__1__16_,
         matrix_mul_2D_3__1__15_, matrix_mul_2D_3__1__14_,
         matrix_mul_2D_3__1__13_, matrix_mul_2D_3__1__12_,
         matrix_mul_2D_3__1__11_, matrix_mul_2D_3__1__10_,
         matrix_mul_2D_3__1__9_, matrix_mul_2D_3__1__8_,
         matrix_mul_2D_3__1__7_, matrix_mul_2D_3__1__6_,
         matrix_mul_2D_3__1__5_, matrix_mul_2D_3__1__4_,
         matrix_mul_2D_3__1__3_, matrix_mul_2D_3__1__2_,
         matrix_mul_2D_3__1__1_, matrix_mul_2D_3__1__0_,
         matrix_mul_2D_3__2__20_, matrix_mul_2D_3__2__19_,
         matrix_mul_2D_3__2__18_, matrix_mul_2D_3__2__17_,
         matrix_mul_2D_3__2__16_, matrix_mul_2D_3__2__15_,
         matrix_mul_2D_3__2__14_, matrix_mul_2D_3__2__13_,
         matrix_mul_2D_3__2__12_, matrix_mul_2D_3__2__11_,
         matrix_mul_2D_3__2__10_, matrix_mul_2D_3__2__9_,
         matrix_mul_2D_3__2__8_, matrix_mul_2D_3__2__7_,
         matrix_mul_2D_3__2__6_, matrix_mul_2D_3__2__5_,
         matrix_mul_2D_3__2__4_, matrix_mul_2D_3__2__3_,
         matrix_mul_2D_3__2__2_, matrix_mul_2D_3__2__1_,
         matrix_mul_2D_3__2__0_, matrix_mul_2D_3__3__20_,
         matrix_mul_2D_3__3__19_, matrix_mul_2D_3__3__18_,
         matrix_mul_2D_3__3__17_, matrix_mul_2D_3__3__16_,
         matrix_mul_2D_3__3__15_, matrix_mul_2D_3__3__14_,
         matrix_mul_2D_3__3__13_, matrix_mul_2D_3__3__12_,
         matrix_mul_2D_3__3__11_, matrix_mul_2D_3__3__10_,
         matrix_mul_2D_3__3__9_, matrix_mul_2D_3__3__8_,
         matrix_mul_2D_3__3__7_, matrix_mul_2D_3__3__6_,
         matrix_mul_2D_3__3__5_, matrix_mul_2D_3__3__4_,
         matrix_mul_2D_3__3__3_, matrix_mul_2D_3__3__2_,
         matrix_mul_2D_3__3__1_, matrix_mul_2D_3__3__0_,
         matrix_mul_2D_3__4__20_, matrix_mul_2D_3__4__19_,
         matrix_mul_2D_3__4__18_, matrix_mul_2D_3__4__17_,
         matrix_mul_2D_3__4__16_, matrix_mul_2D_3__4__15_,
         matrix_mul_2D_3__4__14_, matrix_mul_2D_3__4__13_,
         matrix_mul_2D_3__4__12_, matrix_mul_2D_3__4__11_,
         matrix_mul_2D_3__4__10_, matrix_mul_2D_3__4__9_,
         matrix_mul_2D_3__4__8_, matrix_mul_2D_3__4__7_,
         matrix_mul_2D_3__4__6_, matrix_mul_2D_3__4__5_,
         matrix_mul_2D_3__4__4_, matrix_mul_2D_3__4__3_,
         matrix_mul_2D_3__4__2_, matrix_mul_2D_3__4__1_,
         matrix_mul_2D_3__4__0_, matrix_mul_2D_3__5__20_,
         matrix_mul_2D_3__5__19_, matrix_mul_2D_3__5__18_,
         matrix_mul_2D_3__5__17_, matrix_mul_2D_3__5__16_,
         matrix_mul_2D_3__5__15_, matrix_mul_2D_3__5__14_,
         matrix_mul_2D_3__5__13_, matrix_mul_2D_3__5__12_,
         matrix_mul_2D_3__5__11_, matrix_mul_2D_3__5__10_,
         matrix_mul_2D_3__5__9_, matrix_mul_2D_3__5__8_,
         matrix_mul_2D_3__5__7_, matrix_mul_2D_3__5__6_,
         matrix_mul_2D_3__5__5_, matrix_mul_2D_3__5__4_,
         matrix_mul_2D_3__5__3_, matrix_mul_2D_3__5__2_,
         matrix_mul_2D_3__5__1_, matrix_mul_2D_3__5__0_,
         matrix_mul_2D_3__6__20_, matrix_mul_2D_3__6__19_,
         matrix_mul_2D_3__6__18_, matrix_mul_2D_3__6__17_,
         matrix_mul_2D_3__6__16_, matrix_mul_2D_3__6__15_,
         matrix_mul_2D_3__6__14_, matrix_mul_2D_3__6__13_,
         matrix_mul_2D_3__6__12_, matrix_mul_2D_3__6__11_,
         matrix_mul_2D_3__6__10_, matrix_mul_2D_3__6__9_,
         matrix_mul_2D_3__6__8_, matrix_mul_2D_3__6__7_,
         matrix_mul_2D_3__6__6_, matrix_mul_2D_3__6__5_,
         matrix_mul_2D_3__6__4_, matrix_mul_2D_3__6__3_,
         matrix_mul_2D_3__6__2_, matrix_mul_2D_3__6__1_,
         matrix_mul_2D_3__6__0_, matrix_mul_2D_3__7__20_,
         matrix_mul_2D_3__7__19_, matrix_mul_2D_3__7__18_,
         matrix_mul_2D_3__7__17_, matrix_mul_2D_3__7__16_,
         matrix_mul_2D_3__7__15_, matrix_mul_2D_3__7__14_,
         matrix_mul_2D_3__7__13_, matrix_mul_2D_3__7__12_,
         matrix_mul_2D_3__7__11_, matrix_mul_2D_3__7__10_,
         matrix_mul_2D_3__7__9_, matrix_mul_2D_3__7__8_,
         matrix_mul_2D_3__7__7_, matrix_mul_2D_3__7__6_,
         matrix_mul_2D_3__7__5_, matrix_mul_2D_3__7__4_,
         matrix_mul_2D_3__7__3_, matrix_mul_2D_3__7__2_,
         matrix_mul_2D_3__7__1_, matrix_mul_2D_3__7__0_,
         matrix_mul_2D_4__0__20_, matrix_mul_2D_4__0__19_,
         matrix_mul_2D_4__0__18_, matrix_mul_2D_4__0__17_,
         matrix_mul_2D_4__0__16_, matrix_mul_2D_4__0__15_,
         matrix_mul_2D_4__0__14_, matrix_mul_2D_4__0__13_,
         matrix_mul_2D_4__0__12_, matrix_mul_2D_4__0__11_,
         matrix_mul_2D_4__0__10_, matrix_mul_2D_4__0__9_,
         matrix_mul_2D_4__0__8_, matrix_mul_2D_4__0__7_,
         matrix_mul_2D_4__0__6_, matrix_mul_2D_4__0__5_,
         matrix_mul_2D_4__0__4_, matrix_mul_2D_4__0__3_,
         matrix_mul_2D_4__0__2_, matrix_mul_2D_4__0__1_,
         matrix_mul_2D_4__0__0_, matrix_mul_2D_4__1__20_,
         matrix_mul_2D_4__1__19_, matrix_mul_2D_4__1__18_,
         matrix_mul_2D_4__1__17_, matrix_mul_2D_4__1__16_,
         matrix_mul_2D_4__1__15_, matrix_mul_2D_4__1__14_,
         matrix_mul_2D_4__1__13_, matrix_mul_2D_4__1__12_,
         matrix_mul_2D_4__1__11_, matrix_mul_2D_4__1__10_,
         matrix_mul_2D_4__1__9_, matrix_mul_2D_4__1__8_,
         matrix_mul_2D_4__1__7_, matrix_mul_2D_4__1__6_,
         matrix_mul_2D_4__1__5_, matrix_mul_2D_4__1__4_,
         matrix_mul_2D_4__1__3_, matrix_mul_2D_4__1__2_,
         matrix_mul_2D_4__1__1_, matrix_mul_2D_4__1__0_,
         matrix_mul_2D_4__2__20_, matrix_mul_2D_4__2__19_,
         matrix_mul_2D_4__2__18_, matrix_mul_2D_4__2__17_,
         matrix_mul_2D_4__2__16_, matrix_mul_2D_4__2__15_,
         matrix_mul_2D_4__2__14_, matrix_mul_2D_4__2__13_,
         matrix_mul_2D_4__2__12_, matrix_mul_2D_4__2__11_,
         matrix_mul_2D_4__2__10_, matrix_mul_2D_4__2__9_,
         matrix_mul_2D_4__2__8_, matrix_mul_2D_4__2__7_,
         matrix_mul_2D_4__2__6_, matrix_mul_2D_4__2__5_,
         matrix_mul_2D_4__2__4_, matrix_mul_2D_4__2__3_,
         matrix_mul_2D_4__2__2_, matrix_mul_2D_4__2__1_,
         matrix_mul_2D_4__2__0_, matrix_mul_2D_4__3__20_,
         matrix_mul_2D_4__3__19_, matrix_mul_2D_4__3__18_,
         matrix_mul_2D_4__3__17_, matrix_mul_2D_4__3__16_,
         matrix_mul_2D_4__3__15_, matrix_mul_2D_4__3__14_,
         matrix_mul_2D_4__3__13_, matrix_mul_2D_4__3__12_,
         matrix_mul_2D_4__3__11_, matrix_mul_2D_4__3__10_,
         matrix_mul_2D_4__3__9_, matrix_mul_2D_4__3__8_,
         matrix_mul_2D_4__3__7_, matrix_mul_2D_4__3__6_,
         matrix_mul_2D_4__3__5_, matrix_mul_2D_4__3__4_,
         matrix_mul_2D_4__3__3_, matrix_mul_2D_4__3__2_,
         matrix_mul_2D_4__3__1_, matrix_mul_2D_4__3__0_,
         matrix_mul_2D_4__4__20_, matrix_mul_2D_4__4__19_,
         matrix_mul_2D_4__4__18_, matrix_mul_2D_4__4__17_,
         matrix_mul_2D_4__4__16_, matrix_mul_2D_4__4__15_,
         matrix_mul_2D_4__4__14_, matrix_mul_2D_4__4__13_,
         matrix_mul_2D_4__4__12_, matrix_mul_2D_4__4__11_,
         matrix_mul_2D_4__4__10_, matrix_mul_2D_4__4__9_,
         matrix_mul_2D_4__4__8_, matrix_mul_2D_4__4__7_,
         matrix_mul_2D_4__4__6_, matrix_mul_2D_4__4__5_,
         matrix_mul_2D_4__4__4_, matrix_mul_2D_4__4__3_,
         matrix_mul_2D_4__4__2_, matrix_mul_2D_4__4__1_,
         matrix_mul_2D_4__4__0_, matrix_mul_2D_4__5__20_,
         matrix_mul_2D_4__5__19_, matrix_mul_2D_4__5__18_,
         matrix_mul_2D_4__5__17_, matrix_mul_2D_4__5__16_,
         matrix_mul_2D_4__5__15_, matrix_mul_2D_4__5__14_,
         matrix_mul_2D_4__5__13_, matrix_mul_2D_4__5__12_,
         matrix_mul_2D_4__5__11_, matrix_mul_2D_4__5__10_,
         matrix_mul_2D_4__5__9_, matrix_mul_2D_4__5__8_,
         matrix_mul_2D_4__5__7_, matrix_mul_2D_4__5__6_,
         matrix_mul_2D_4__5__5_, matrix_mul_2D_4__5__4_,
         matrix_mul_2D_4__5__3_, matrix_mul_2D_4__5__2_,
         matrix_mul_2D_4__5__1_, matrix_mul_2D_4__5__0_,
         matrix_mul_2D_4__6__20_, matrix_mul_2D_4__6__19_,
         matrix_mul_2D_4__6__18_, matrix_mul_2D_4__6__17_,
         matrix_mul_2D_4__6__16_, matrix_mul_2D_4__6__15_,
         matrix_mul_2D_4__6__14_, matrix_mul_2D_4__6__13_,
         matrix_mul_2D_4__6__12_, matrix_mul_2D_4__6__11_,
         matrix_mul_2D_4__6__10_, matrix_mul_2D_4__6__9_,
         matrix_mul_2D_4__6__8_, matrix_mul_2D_4__6__7_,
         matrix_mul_2D_4__6__6_, matrix_mul_2D_4__6__5_,
         matrix_mul_2D_4__6__4_, matrix_mul_2D_4__6__3_,
         matrix_mul_2D_4__6__2_, matrix_mul_2D_4__6__1_,
         matrix_mul_2D_4__6__0_, matrix_mul_2D_4__7__20_,
         matrix_mul_2D_4__7__19_, matrix_mul_2D_4__7__18_,
         matrix_mul_2D_4__7__17_, matrix_mul_2D_4__7__16_,
         matrix_mul_2D_4__7__15_, matrix_mul_2D_4__7__14_,
         matrix_mul_2D_4__7__13_, matrix_mul_2D_4__7__12_,
         matrix_mul_2D_4__7__11_, matrix_mul_2D_4__7__10_,
         matrix_mul_2D_4__7__9_, matrix_mul_2D_4__7__8_,
         matrix_mul_2D_4__7__7_, matrix_mul_2D_4__7__6_,
         matrix_mul_2D_4__7__5_, matrix_mul_2D_4__7__4_,
         matrix_mul_2D_4__7__3_, matrix_mul_2D_4__7__2_,
         matrix_mul_2D_4__7__1_, matrix_mul_2D_4__7__0_,
         matrix_mul_2D_5__0__20_, matrix_mul_2D_5__0__19_,
         matrix_mul_2D_5__0__18_, matrix_mul_2D_5__0__17_,
         matrix_mul_2D_5__0__16_, matrix_mul_2D_5__0__15_,
         matrix_mul_2D_5__0__14_, matrix_mul_2D_5__0__13_,
         matrix_mul_2D_5__0__12_, matrix_mul_2D_5__0__11_,
         matrix_mul_2D_5__0__10_, matrix_mul_2D_5__0__9_,
         matrix_mul_2D_5__0__8_, matrix_mul_2D_5__0__7_,
         matrix_mul_2D_5__0__6_, matrix_mul_2D_5__0__5_,
         matrix_mul_2D_5__0__4_, matrix_mul_2D_5__0__3_,
         matrix_mul_2D_5__0__2_, matrix_mul_2D_5__0__1_,
         matrix_mul_2D_5__0__0_, matrix_mul_2D_5__1__20_,
         matrix_mul_2D_5__1__19_, matrix_mul_2D_5__1__18_,
         matrix_mul_2D_5__1__17_, matrix_mul_2D_5__1__16_,
         matrix_mul_2D_5__1__15_, matrix_mul_2D_5__1__14_,
         matrix_mul_2D_5__1__13_, matrix_mul_2D_5__1__12_,
         matrix_mul_2D_5__1__11_, matrix_mul_2D_5__1__10_,
         matrix_mul_2D_5__1__9_, matrix_mul_2D_5__1__8_,
         matrix_mul_2D_5__1__7_, matrix_mul_2D_5__1__6_,
         matrix_mul_2D_5__1__5_, matrix_mul_2D_5__1__4_,
         matrix_mul_2D_5__1__3_, matrix_mul_2D_5__1__2_,
         matrix_mul_2D_5__1__1_, matrix_mul_2D_5__1__0_,
         matrix_mul_2D_5__2__20_, matrix_mul_2D_5__2__19_,
         matrix_mul_2D_5__2__18_, matrix_mul_2D_5__2__17_,
         matrix_mul_2D_5__2__16_, matrix_mul_2D_5__2__15_,
         matrix_mul_2D_5__2__14_, matrix_mul_2D_5__2__13_,
         matrix_mul_2D_5__2__12_, matrix_mul_2D_5__2__11_,
         matrix_mul_2D_5__2__10_, matrix_mul_2D_5__2__9_,
         matrix_mul_2D_5__2__8_, matrix_mul_2D_5__2__7_,
         matrix_mul_2D_5__2__6_, matrix_mul_2D_5__2__5_,
         matrix_mul_2D_5__2__4_, matrix_mul_2D_5__2__3_,
         matrix_mul_2D_5__2__2_, matrix_mul_2D_5__2__1_,
         matrix_mul_2D_5__2__0_, matrix_mul_2D_5__3__20_,
         matrix_mul_2D_5__3__19_, matrix_mul_2D_5__3__18_,
         matrix_mul_2D_5__3__17_, matrix_mul_2D_5__3__16_,
         matrix_mul_2D_5__3__15_, matrix_mul_2D_5__3__14_,
         matrix_mul_2D_5__3__13_, matrix_mul_2D_5__3__12_,
         matrix_mul_2D_5__3__11_, matrix_mul_2D_5__3__10_,
         matrix_mul_2D_5__3__9_, matrix_mul_2D_5__3__8_,
         matrix_mul_2D_5__3__7_, matrix_mul_2D_5__3__6_,
         matrix_mul_2D_5__3__5_, matrix_mul_2D_5__3__4_,
         matrix_mul_2D_5__3__3_, matrix_mul_2D_5__3__2_,
         matrix_mul_2D_5__3__1_, matrix_mul_2D_5__3__0_,
         matrix_mul_2D_5__4__20_, matrix_mul_2D_5__4__19_,
         matrix_mul_2D_5__4__18_, matrix_mul_2D_5__4__17_,
         matrix_mul_2D_5__4__16_, matrix_mul_2D_5__4__15_,
         matrix_mul_2D_5__4__14_, matrix_mul_2D_5__4__13_,
         matrix_mul_2D_5__4__12_, matrix_mul_2D_5__4__11_,
         matrix_mul_2D_5__4__10_, matrix_mul_2D_5__4__9_,
         matrix_mul_2D_5__4__8_, matrix_mul_2D_5__4__7_,
         matrix_mul_2D_5__4__6_, matrix_mul_2D_5__4__5_,
         matrix_mul_2D_5__4__4_, matrix_mul_2D_5__4__3_,
         matrix_mul_2D_5__4__2_, matrix_mul_2D_5__4__1_,
         matrix_mul_2D_5__4__0_, matrix_mul_2D_5__5__20_,
         matrix_mul_2D_5__5__19_, matrix_mul_2D_5__5__18_,
         matrix_mul_2D_5__5__17_, matrix_mul_2D_5__5__16_,
         matrix_mul_2D_5__5__15_, matrix_mul_2D_5__5__14_,
         matrix_mul_2D_5__5__13_, matrix_mul_2D_5__5__12_,
         matrix_mul_2D_5__5__11_, matrix_mul_2D_5__5__10_,
         matrix_mul_2D_5__5__9_, matrix_mul_2D_5__5__8_,
         matrix_mul_2D_5__5__7_, matrix_mul_2D_5__5__6_,
         matrix_mul_2D_5__5__5_, matrix_mul_2D_5__5__4_,
         matrix_mul_2D_5__5__3_, matrix_mul_2D_5__5__2_,
         matrix_mul_2D_5__5__1_, matrix_mul_2D_5__5__0_,
         matrix_mul_2D_5__6__20_, matrix_mul_2D_5__6__19_,
         matrix_mul_2D_5__6__18_, matrix_mul_2D_5__6__17_,
         matrix_mul_2D_5__6__16_, matrix_mul_2D_5__6__15_,
         matrix_mul_2D_5__6__14_, matrix_mul_2D_5__6__13_,
         matrix_mul_2D_5__6__12_, matrix_mul_2D_5__6__11_,
         matrix_mul_2D_5__6__10_, matrix_mul_2D_5__6__9_,
         matrix_mul_2D_5__6__8_, matrix_mul_2D_5__6__7_,
         matrix_mul_2D_5__6__6_, matrix_mul_2D_5__6__5_,
         matrix_mul_2D_5__6__4_, matrix_mul_2D_5__6__3_,
         matrix_mul_2D_5__6__2_, matrix_mul_2D_5__6__1_,
         matrix_mul_2D_5__6__0_, matrix_mul_2D_5__7__20_,
         matrix_mul_2D_5__7__19_, matrix_mul_2D_5__7__18_,
         matrix_mul_2D_5__7__17_, matrix_mul_2D_5__7__16_,
         matrix_mul_2D_5__7__15_, matrix_mul_2D_5__7__14_,
         matrix_mul_2D_5__7__13_, matrix_mul_2D_5__7__12_,
         matrix_mul_2D_5__7__11_, matrix_mul_2D_5__7__10_,
         matrix_mul_2D_5__7__9_, matrix_mul_2D_5__7__8_,
         matrix_mul_2D_5__7__7_, matrix_mul_2D_5__7__6_,
         matrix_mul_2D_5__7__5_, matrix_mul_2D_5__7__4_,
         matrix_mul_2D_5__7__3_, matrix_mul_2D_5__7__2_,
         matrix_mul_2D_5__7__1_, matrix_mul_2D_5__7__0_,
         matrix_mul_2D_6__0__20_, matrix_mul_2D_6__0__19_,
         matrix_mul_2D_6__0__18_, matrix_mul_2D_6__0__17_,
         matrix_mul_2D_6__0__16_, matrix_mul_2D_6__0__15_,
         matrix_mul_2D_6__0__14_, matrix_mul_2D_6__0__13_,
         matrix_mul_2D_6__0__12_, matrix_mul_2D_6__0__11_,
         matrix_mul_2D_6__0__10_, matrix_mul_2D_6__0__9_,
         matrix_mul_2D_6__0__8_, matrix_mul_2D_6__0__7_,
         matrix_mul_2D_6__0__6_, matrix_mul_2D_6__0__5_,
         matrix_mul_2D_6__0__4_, matrix_mul_2D_6__0__3_,
         matrix_mul_2D_6__0__2_, matrix_mul_2D_6__0__1_,
         matrix_mul_2D_6__0__0_, matrix_mul_2D_6__1__20_,
         matrix_mul_2D_6__1__19_, matrix_mul_2D_6__1__18_,
         matrix_mul_2D_6__1__17_, matrix_mul_2D_6__1__16_,
         matrix_mul_2D_6__1__15_, matrix_mul_2D_6__1__14_,
         matrix_mul_2D_6__1__13_, matrix_mul_2D_6__1__12_,
         matrix_mul_2D_6__1__11_, matrix_mul_2D_6__1__10_,
         matrix_mul_2D_6__1__9_, matrix_mul_2D_6__1__8_,
         matrix_mul_2D_6__1__7_, matrix_mul_2D_6__1__6_,
         matrix_mul_2D_6__1__5_, matrix_mul_2D_6__1__4_,
         matrix_mul_2D_6__1__3_, matrix_mul_2D_6__1__2_,
         matrix_mul_2D_6__1__1_, matrix_mul_2D_6__1__0_,
         matrix_mul_2D_6__2__20_, matrix_mul_2D_6__2__19_,
         matrix_mul_2D_6__2__18_, matrix_mul_2D_6__2__17_,
         matrix_mul_2D_6__2__16_, matrix_mul_2D_6__2__15_,
         matrix_mul_2D_6__2__14_, matrix_mul_2D_6__2__13_,
         matrix_mul_2D_6__2__12_, matrix_mul_2D_6__2__11_,
         matrix_mul_2D_6__2__10_, matrix_mul_2D_6__2__9_,
         matrix_mul_2D_6__2__8_, matrix_mul_2D_6__2__7_,
         matrix_mul_2D_6__2__6_, matrix_mul_2D_6__2__5_,
         matrix_mul_2D_6__2__4_, matrix_mul_2D_6__2__3_,
         matrix_mul_2D_6__2__2_, matrix_mul_2D_6__2__1_,
         matrix_mul_2D_6__2__0_, matrix_mul_2D_6__3__20_,
         matrix_mul_2D_6__3__19_, matrix_mul_2D_6__3__18_,
         matrix_mul_2D_6__3__17_, matrix_mul_2D_6__3__16_,
         matrix_mul_2D_6__3__15_, matrix_mul_2D_6__3__14_,
         matrix_mul_2D_6__3__13_, matrix_mul_2D_6__3__12_,
         matrix_mul_2D_6__3__11_, matrix_mul_2D_6__3__10_,
         matrix_mul_2D_6__3__9_, matrix_mul_2D_6__3__8_,
         matrix_mul_2D_6__3__7_, matrix_mul_2D_6__3__6_,
         matrix_mul_2D_6__3__5_, matrix_mul_2D_6__3__4_,
         matrix_mul_2D_6__3__3_, matrix_mul_2D_6__3__2_,
         matrix_mul_2D_6__3__1_, matrix_mul_2D_6__3__0_,
         matrix_mul_2D_6__4__20_, matrix_mul_2D_6__4__19_,
         matrix_mul_2D_6__4__18_, matrix_mul_2D_6__4__17_,
         matrix_mul_2D_6__4__16_, matrix_mul_2D_6__4__15_,
         matrix_mul_2D_6__4__14_, matrix_mul_2D_6__4__13_,
         matrix_mul_2D_6__4__12_, matrix_mul_2D_6__4__11_,
         matrix_mul_2D_6__4__10_, matrix_mul_2D_6__4__9_,
         matrix_mul_2D_6__4__8_, matrix_mul_2D_6__4__7_,
         matrix_mul_2D_6__4__6_, matrix_mul_2D_6__4__5_,
         matrix_mul_2D_6__4__4_, matrix_mul_2D_6__4__3_,
         matrix_mul_2D_6__4__2_, matrix_mul_2D_6__4__1_,
         matrix_mul_2D_6__4__0_, matrix_mul_2D_6__5__20_,
         matrix_mul_2D_6__5__19_, matrix_mul_2D_6__5__18_,
         matrix_mul_2D_6__5__17_, matrix_mul_2D_6__5__16_,
         matrix_mul_2D_6__5__15_, matrix_mul_2D_6__5__14_,
         matrix_mul_2D_6__5__13_, matrix_mul_2D_6__5__12_,
         matrix_mul_2D_6__5__11_, matrix_mul_2D_6__5__10_,
         matrix_mul_2D_6__5__9_, matrix_mul_2D_6__5__8_,
         matrix_mul_2D_6__5__7_, matrix_mul_2D_6__5__6_,
         matrix_mul_2D_6__5__5_, matrix_mul_2D_6__5__4_,
         matrix_mul_2D_6__5__3_, matrix_mul_2D_6__5__2_,
         matrix_mul_2D_6__5__1_, matrix_mul_2D_6__5__0_,
         matrix_mul_2D_6__6__20_, matrix_mul_2D_6__6__19_,
         matrix_mul_2D_6__6__18_, matrix_mul_2D_6__6__17_,
         matrix_mul_2D_6__6__16_, matrix_mul_2D_6__6__15_,
         matrix_mul_2D_6__6__14_, matrix_mul_2D_6__6__13_,
         matrix_mul_2D_6__6__12_, matrix_mul_2D_6__6__11_,
         matrix_mul_2D_6__6__10_, matrix_mul_2D_6__6__9_,
         matrix_mul_2D_6__6__8_, matrix_mul_2D_6__6__7_,
         matrix_mul_2D_6__6__6_, matrix_mul_2D_6__6__5_,
         matrix_mul_2D_6__6__4_, matrix_mul_2D_6__6__3_,
         matrix_mul_2D_6__6__2_, matrix_mul_2D_6__6__1_,
         matrix_mul_2D_6__6__0_, matrix_mul_2D_6__7__20_,
         matrix_mul_2D_6__7__19_, matrix_mul_2D_6__7__18_,
         matrix_mul_2D_6__7__17_, matrix_mul_2D_6__7__16_,
         matrix_mul_2D_6__7__15_, matrix_mul_2D_6__7__14_,
         matrix_mul_2D_6__7__13_, matrix_mul_2D_6__7__12_,
         matrix_mul_2D_6__7__11_, matrix_mul_2D_6__7__10_,
         matrix_mul_2D_6__7__9_, matrix_mul_2D_6__7__8_,
         matrix_mul_2D_6__7__7_, matrix_mul_2D_6__7__6_,
         matrix_mul_2D_6__7__5_, matrix_mul_2D_6__7__4_,
         matrix_mul_2D_6__7__3_, matrix_mul_2D_6__7__2_,
         matrix_mul_2D_6__7__1_, matrix_mul_2D_6__7__0_,
         matrix_mul_2D_7__0__20_, matrix_mul_2D_7__0__19_,
         matrix_mul_2D_7__0__18_, matrix_mul_2D_7__0__17_,
         matrix_mul_2D_7__0__16_, matrix_mul_2D_7__0__15_,
         matrix_mul_2D_7__0__14_, matrix_mul_2D_7__0__13_,
         matrix_mul_2D_7__0__12_, matrix_mul_2D_7__0__11_,
         matrix_mul_2D_7__0__10_, matrix_mul_2D_7__0__9_,
         matrix_mul_2D_7__0__8_, matrix_mul_2D_7__0__7_,
         matrix_mul_2D_7__0__6_, matrix_mul_2D_7__0__5_,
         matrix_mul_2D_7__0__4_, matrix_mul_2D_7__0__3_,
         matrix_mul_2D_7__0__2_, matrix_mul_2D_7__0__1_,
         matrix_mul_2D_7__0__0_, matrix_mul_2D_7__1__20_,
         matrix_mul_2D_7__1__19_, matrix_mul_2D_7__1__18_,
         matrix_mul_2D_7__1__17_, matrix_mul_2D_7__1__16_,
         matrix_mul_2D_7__1__15_, matrix_mul_2D_7__1__14_,
         matrix_mul_2D_7__1__13_, matrix_mul_2D_7__1__12_,
         matrix_mul_2D_7__1__11_, matrix_mul_2D_7__1__10_,
         matrix_mul_2D_7__1__9_, matrix_mul_2D_7__1__8_,
         matrix_mul_2D_7__1__7_, matrix_mul_2D_7__1__6_,
         matrix_mul_2D_7__1__5_, matrix_mul_2D_7__1__4_,
         matrix_mul_2D_7__1__3_, matrix_mul_2D_7__1__2_,
         matrix_mul_2D_7__1__1_, matrix_mul_2D_7__1__0_,
         matrix_mul_2D_7__2__20_, matrix_mul_2D_7__2__19_,
         matrix_mul_2D_7__2__18_, matrix_mul_2D_7__2__17_,
         matrix_mul_2D_7__2__16_, matrix_mul_2D_7__2__15_,
         matrix_mul_2D_7__2__14_, matrix_mul_2D_7__2__13_,
         matrix_mul_2D_7__2__12_, matrix_mul_2D_7__2__11_,
         matrix_mul_2D_7__2__10_, matrix_mul_2D_7__2__9_,
         matrix_mul_2D_7__2__8_, matrix_mul_2D_7__2__7_,
         matrix_mul_2D_7__2__6_, matrix_mul_2D_7__2__5_,
         matrix_mul_2D_7__2__4_, matrix_mul_2D_7__2__3_,
         matrix_mul_2D_7__2__2_, matrix_mul_2D_7__2__1_,
         matrix_mul_2D_7__2__0_, matrix_mul_2D_7__3__20_,
         matrix_mul_2D_7__3__19_, matrix_mul_2D_7__3__18_,
         matrix_mul_2D_7__3__17_, matrix_mul_2D_7__3__16_,
         matrix_mul_2D_7__3__15_, matrix_mul_2D_7__3__14_,
         matrix_mul_2D_7__3__13_, matrix_mul_2D_7__3__12_,
         matrix_mul_2D_7__3__11_, matrix_mul_2D_7__3__10_,
         matrix_mul_2D_7__3__9_, matrix_mul_2D_7__3__8_,
         matrix_mul_2D_7__3__7_, matrix_mul_2D_7__3__6_,
         matrix_mul_2D_7__3__5_, matrix_mul_2D_7__3__4_,
         matrix_mul_2D_7__3__3_, matrix_mul_2D_7__3__2_,
         matrix_mul_2D_7__3__1_, matrix_mul_2D_7__3__0_,
         matrix_mul_2D_7__4__20_, matrix_mul_2D_7__4__19_,
         matrix_mul_2D_7__4__18_, matrix_mul_2D_7__4__17_,
         matrix_mul_2D_7__4__16_, matrix_mul_2D_7__4__15_,
         matrix_mul_2D_7__4__14_, matrix_mul_2D_7__4__13_,
         matrix_mul_2D_7__4__12_, matrix_mul_2D_7__4__11_,
         matrix_mul_2D_7__4__10_, matrix_mul_2D_7__4__9_,
         matrix_mul_2D_7__4__8_, matrix_mul_2D_7__4__7_,
         matrix_mul_2D_7__4__6_, matrix_mul_2D_7__4__5_,
         matrix_mul_2D_7__4__4_, matrix_mul_2D_7__4__3_,
         matrix_mul_2D_7__4__2_, matrix_mul_2D_7__4__1_,
         matrix_mul_2D_7__4__0_, matrix_mul_2D_7__5__20_,
         matrix_mul_2D_7__5__19_, matrix_mul_2D_7__5__18_,
         matrix_mul_2D_7__5__17_, matrix_mul_2D_7__5__16_,
         matrix_mul_2D_7__5__15_, matrix_mul_2D_7__5__14_,
         matrix_mul_2D_7__5__13_, matrix_mul_2D_7__5__12_,
         matrix_mul_2D_7__5__11_, matrix_mul_2D_7__5__10_,
         matrix_mul_2D_7__5__9_, matrix_mul_2D_7__5__8_,
         matrix_mul_2D_7__5__7_, matrix_mul_2D_7__5__6_,
         matrix_mul_2D_7__5__5_, matrix_mul_2D_7__5__4_,
         matrix_mul_2D_7__5__3_, matrix_mul_2D_7__5__2_,
         matrix_mul_2D_7__5__1_, matrix_mul_2D_7__5__0_,
         matrix_mul_2D_7__6__20_, matrix_mul_2D_7__6__19_,
         matrix_mul_2D_7__6__18_, matrix_mul_2D_7__6__17_,
         matrix_mul_2D_7__6__16_, matrix_mul_2D_7__6__15_,
         matrix_mul_2D_7__6__14_, matrix_mul_2D_7__6__13_,
         matrix_mul_2D_7__6__12_, matrix_mul_2D_7__6__11_,
         matrix_mul_2D_7__6__10_, matrix_mul_2D_7__6__9_,
         matrix_mul_2D_7__6__8_, matrix_mul_2D_7__6__7_,
         matrix_mul_2D_7__6__6_, matrix_mul_2D_7__6__5_,
         matrix_mul_2D_7__6__4_, matrix_mul_2D_7__6__3_,
         matrix_mul_2D_7__6__2_, matrix_mul_2D_7__6__1_,
         matrix_mul_2D_7__6__0_, matrix_mul_2D_7__7__20_,
         matrix_mul_2D_7__7__19_, matrix_mul_2D_7__7__18_,
         matrix_mul_2D_7__7__17_, matrix_mul_2D_7__7__16_,
         matrix_mul_2D_7__7__15_, matrix_mul_2D_7__7__14_,
         matrix_mul_2D_7__7__13_, matrix_mul_2D_7__7__12_,
         matrix_mul_2D_7__7__11_, matrix_mul_2D_7__7__10_,
         matrix_mul_2D_7__7__9_, matrix_mul_2D_7__7__8_,
         matrix_mul_2D_7__7__7_, matrix_mul_2D_7__7__6_,
         matrix_mul_2D_7__7__5_, matrix_mul_2D_7__7__4_,
         matrix_mul_2D_7__7__3_, matrix_mul_2D_7__7__2_,
         matrix_mul_2D_7__7__1_, matrix_mul_2D_7__7__0_, N2559, N2560, N2561,
         N2562, N2563, N2564, N2565, N2566, N2567, N2568, N2569, N2570, N2571,
         N2572, N2573, N2574, N2592, N2593, N2594, N2595, N2596, N2597, N2598,
         N2599, N2600, N2601, N2602, N2603, N2604, N2605, N2606, N2607, N2608,
         N2609, N2610, N2611, N2612, N2637, N2641, N2642, N2643, N2644, N2645,
         N2646, N2647, N2648, N2649, N2650, N2651, N2652, N2653, N2654, N2655,
         N2656, N2674, N2675, N2676, N2677, N2678, N2679, N2680, N2681, N2682,
         N2683, N2684, N2685, N2686, N2687, N2688, N2689, N2690, N2691, N2692,
         N2693, N2694, N2729, N2733, N2734, N2735, N2736, N2737, N2738, N2739,
         N2740, N2741, N2742, N2743, N2744, N2745, N2746, N2747, N2748, N2766,
         N2767, N2768, N2769, N2770, N2771, N2772, N2773, N2774, N2775, N2776,
         N2777, N2778, N2779, N2780, N2781, N2782, N2783, N2784, N2785, N2786,
         N2811, N2815, N2816, N2817, N2818, N2819, N2820, N2821, N2822, N2823,
         N2824, N2825, N2826, N2827, N2828, N2829, N2830, N2848, N2849, N2850,
         N2851, N2852, N2853, N2854, N2855, N2856, N2857, N2858, N2859, N2860,
         N2861, N2862, N2863, N2864, N2865, N2866, N2867, N2868, N2903, N2907,
         N2908, N2909, N2910, N2911, N2912, N2913, N2914, N2915, N2916, N2917,
         N2918, N2919, N2920, N2921, N2922, N2940, N2941, N2942, N2943, N2944,
         N2945, N2946, N2947, N2948, N2949, N2950, N2951, N2952, N2953, N2954,
         N2955, N2956, N2957, N2958, N2959, N2960, N2985, N2989, N2990, N2991,
         N2992, N2993, N2994, N2995, N2996, N2997, N2998, N2999, N3000, N3001,
         N3002, N3003, N3004, N3022, N3023, N3024, N3025, N3026, N3027, N3028,
         N3029, N3030, N3031, N3032, N3033, N3034, N3035, N3036, N3037, N3038,
         N3039, N3040, N3041, N3042, N3081, N3082, N3083, N3084, N3085, N3086,
         N3087, N3088, N3089, N3090, N3091, N3092, N3093, N3094, N3095, N3096,
         N3114, N3115, N3116, N3117, N3118, N3119, N3120, N3121, N3122, N3123,
         N3124, N3125, N3126, N3127, N3128, N3129, N3130, N3131, N3132, N3133,
         N3134, N3163, N3164, N3165, N3166, N3167, N3168, N3169, N3170, N3171,
         N3172, N3173, N3174, N3175, N3176, N3177, N3178, N3196, N3197, N3198,
         N3199, N3200, N3201, N3202, N3203, N3204, N3205, N3206, N3207, N3208,
         N3209, N3210, N3211, N3212, N3213, N3214, N3215, N3216, N3252, N3253,
         N3254, N3255, N3256, N3257, N3258, N3259, N3260, N3261, N3262, N3263,
         N3264, N3265, N3266, N3267, N3285, N3286, N3287, N3288, N3289, N3290,
         N3291, N3292, N3293, N3294, N3295, N3296, N3297, N3298, N3299, N3300,
         N3301, N3302, N3303, N3304, N3305, N3331, N3332, N3333, N3334, N3335,
         N3336, N3337, N3338, N3339, N3340, N3341, N3342, N3343, N3344, N3345,
         N3346, N3364, N3365, N3366, N3367, N3368, N3369, N3370, N3371, N3372,
         N3373, N3374, N3375, N3376, N3377, N3378, N3379, N3380, N3381, N3382,
         N3383, N3384, N3420, N3421, N3422, N3423, N3424, N3425, N3426, N3427,
         N3428, N3429, N3430, N3431, N3432, N3433, N3434, N3435, N3453, N3454,
         N3455, N3456, N3457, N3458, N3459, N3460, N3461, N3462, N3463, N3464,
         N3465, N3466, N3467, N3468, N3469, N3470, N3471, N3472, N3473, N3499,
         N3500, N3501, N3502, N3503, N3504, N3505, N3506, N3507, N3508, N3509,
         N3510, N3511, N3512, N3513, N3514, N3532, N3533, N3534, N3535, N3536,
         N3537, N3538, N3539, N3540, N3541, N3542, N3543, N3544, N3545, N3546,
         N3547, N3548, N3549, N3550, N3551, N3552, N3588, N3589, N3590, N3591,
         N3592, N3593, N3594, N3595, N3596, N3597, N3598, N3599, N3600, N3601,
         N3602, N3603, N3621, N3622, N3623, N3624, N3625, N3626, N3627, N3628,
         N3629, N3630, N3631, N3632, N3633, N3634, N3635, N3636, N3637, N3638,
         N3639, N3640, N3641, N3667, N3668, N3669, N3670, N3671, N3672, N3673,
         N3674, N3675, N3676, N3677, N3678, N3679, N3680, N3681, N3682, N3700,
         N3701, N3702, N3703, N3704, N3705, N3706, N3707, N3708, N3709, N3710,
         N3711, N3712, N3713, N3714, N3715, N3716, N3717, N3718, N3719, N3720,
         N3756, N3757, N3758, N3759, N3760, N3761, N3762, N3763, N3764, N3765,
         N3766, N3767, N3768, N3769, N3770, N3771, N3789, N3790, N3791, N3792,
         N3793, N3794, N3795, N3796, N3797, N3798, N3799, N3800, N3801, N3802,
         N3803, N3804, N3805, N3806, N3807, N3808, N3809, N3838, N3839, N3840,
         N3841, N3842, N3843, N3844, N3845, N3846, N3847, N3848, N3849, N3850,
         N3851, N3852, N3853, N3871, N3872, N3873, N3874, N3875, N3876, N3877,
         N3878, N3879, N3880, N3881, N3882, N3883, N3884, N3885, N3886, N3887,
         N3888, N3889, N3890, N3891, N3927, N3928, N3929, N3930, N3931, N3932,
         N3933, N3934, N3935, N3936, N3937, N3938, N3939, N3940, N3941, N3942,
         N3960, N3961, N3962, N3963, N3964, N3965, N3966, N3967, N3968, N3969,
         N3970, N3971, N3972, N3973, N3974, N3975, N3976, N3977, N3978, N3979,
         N3980, N4006, N4007, N4008, N4009, N4010, N4011, N4012, N4013, N4014,
         N4015, N4016, N4017, N4018, N4019, N4020, N4021, N4039, N4040, N4041,
         N4042, N4043, N4044, N4045, N4046, N4047, N4048, N4049, N4050, N4051,
         N4052, N4053, N4054, N4055, N4056, N4057, N4058, N4059, N4095, N4096,
         N4097, N4098, N4099, N4100, N4101, N4102, N4103, N4104, N4105, N4106,
         N4107, N4108, N4109, N4110, N4128, N4129, N4130, N4131, N4132, N4133,
         N4134, N4135, N4136, N4137, N4138, N4139, N4140, N4141, N4142, N4143,
         N4144, N4145, N4146, N4147, N4148, N4174, N4175, N4176, N4177, N4178,
         N4179, N4180, N4181, N4182, N4183, N4184, N4185, N4186, N4187, N4188,
         N4189, N4207, N4208, N4209, N4210, N4211, N4212, N4213, N4214, N4215,
         N4216, N4217, N4218, N4219, N4220, N4221, N4222, N4223, N4224, N4225,
         N4226, N4227, N4263, N4264, N4265, N4266, N4267, N4268, N4269, N4270,
         N4271, N4272, N4273, N4274, N4275, N4276, N4277, N4278, N4296, N4297,
         N4298, N4299, N4300, N4301, N4302, N4303, N4304, N4305, N4306, N4307,
         N4308, N4309, N4310, N4311, N4312, N4313, N4314, N4315, N4316, N4342,
         N4343, N4344, N4345, N4346, N4347, N4348, N4349, N4350, N4351, N4352,
         N4353, N4354, N4355, N4356, N4357, N4375, N4376, N4377, N4378, N4379,
         N4380, N4381, N4382, N4383, N4384, N4385, N4386, N4387, N4388, N4389,
         N4390, N4391, N4392, N4393, N4394, N4395, N4431, N4432, N4433, N4434,
         N4435, N4436, N4437, N4438, N4439, N4440, N4441, N4442, N4443, N4444,
         N4445, N4446, N4464, N4465, N4466, N4467, N4468, N4469, N4470, N4471,
         N4472, N4473, N4474, N4475, N4476, N4477, N4478, N4479, N4480, N4481,
         N4482, N4483, N4484, N4509, N4513, N4514, N4515, N4516, N4517, N4518,
         N4519, N4520, N4521, N4522, N4523, N4524, N4525, N4526, N4527, N4528,
         N4546, N4547, N4548, N4549, N4550, N4551, N4552, N4553, N4554, N4555,
         N4556, N4557, N4558, N4559, N4560, N4561, N4562, N4563, N4564, N4565,
         N4566, N4613, N4614, N4615, N4616, N4617, N4618, N4619, N4620, N4621,
         N4622, N4623, N4624, N4625, N4626, N4627, N4628, N4646, N4647, N4648,
         N4649, N4650, N4651, N4652, N4653, N4654, N4655, N4656, N4657, N4658,
         N4659, N4660, N4661, N4662, N4663, N4664, N4665, N4666, N4695, N4696,
         N4697, N4698, N4699, N4700, N4701, N4702, N4703, N4704, N4705, N4706,
         N4707, N4708, N4709, N4710, N4728, N4729, N4730, N4731, N4732, N4733,
         N4734, N4735, N4736, N4737, N4738, N4739, N4740, N4741, N4742, N4743,
         N4744, N4745, N4746, N4747, N4748, N4787, N4788, N4789, N4790, N4791,
         N4792, N4793, N4794, N4795, N4796, N4797, N4798, N4799, N4800, N4801,
         N4802, N4820, N4821, N4822, N4823, N4824, N4825, N4826, N4827, N4828,
         N4829, N4830, N4831, N4832, N4833, N4834, N4835, N4836, N4837, N4838,
         N4839, N4840, N4869, N4870, N4871, N4872, N4873, N4874, N4875, N4876,
         N4877, N4878, N4879, N4880, N4881, N4882, N4883, N4884, N4902, N4903,
         N4904, N4905, N4906, N4907, N4908, N4909, N4910, N4911, N4912, N4913,
         N4914, N4915, N4916, N4917, N4918, N4919, N4920, N4921, N4922, N4961,
         N4962, N4963, N4964, N4965, N4966, N4967, N4968, N4969, N4970, N4971,
         N4972, N4973, N4974, N4975, N4976, N4994, N4995, N4996, N4997, N4998,
         N4999, N5000, N5001, N5002, N5003, N5004, N5005, N5006, N5007, N5008,
         N5009, N5010, N5011, N5012, N5013, N5014, N5043, N5044, N5045, N5046,
         N5047, N5048, N5049, N5050, N5051, N5052, N5053, N5054, N5055, N5056,
         N5057, N5058, N5076, N5077, N5078, N5079, N5080, N5081, N5082, N5083,
         N5084, N5085, N5086, N5087, N5088, N5089, N5090, N5091, N5092, N5093,
         N5094, N5095, N5096, N5135, N5136, N5137, N5138, N5139, N5140, N5141,
         N5142, N5143, N5144, N5145, N5146, N5147, N5148, N5149, N5150, N5168,
         N5169, N5170, N5171, N5172, N5173, N5174, N5175, N5176, N5177, N5178,
         N5179, N5180, N5181, N5182, N5183, N5184, N5185, N5186, N5187, N5188,
         N5213, N5217, N5218, N5219, N5220, N5221, N5222, N5223, N5224, N5225,
         N5226, N5227, N5228, N5229, N5230, N5231, N5232, N5250, N5251, N5252,
         N5253, N5254, N5255, N5256, N5257, N5258, N5259, N5260, N5261, N5262,
         N5263, N5264, N5265, N5266, N5267, N5268, N5269, N5270, N5306, N5307,
         N5308, N5309, N5310, N5311, N5312, N5313, N5314, N5315, N5316, N5317,
         N5318, N5319, N5320, N5321, N5339, N5340, N5341, N5342, N5343, N5344,
         N5345, N5346, N5347, N5348, N5349, N5350, N5351, N5352, N5353, N5354,
         N5355, N5356, N5357, N5358, N5359, N5385, N5386, N5387, N5388, N5389,
         N5390, N5391, N5392, N5393, N5394, N5395, N5396, N5397, N5398, N5399,
         N5400, N5418, N5419, N5420, N5421, N5422, N5423, N5424, N5425, N5426,
         N5427, N5428, N5429, N5430, N5431, N5432, N5433, N5434, N5435, N5436,
         N5437, N5438, N5474, N5475, N5476, N5477, N5478, N5479, N5480, N5481,
         N5482, N5483, N5484, N5485, N5486, N5487, N5488, N5489, N5507, N5508,
         N5509, N5510, N5511, N5512, N5513, N5514, N5515, N5516, N5517, N5518,
         N5519, N5520, N5521, N5522, N5523, N5524, N5525, N5526, N5527, N5553,
         N5554, N5555, N5556, N5557, N5558, N5559, N5560, N5561, N5562, N5563,
         N5564, N5565, N5566, N5567, N5568, N5586, N5587, N5588, N5589, N5590,
         N5591, N5592, N5593, N5594, N5595, N5596, N5597, N5598, N5599, N5600,
         N5601, N5602, N5603, N5604, N5605, N5606, N5642, N5643, N5644, N5645,
         N5646, N5647, N5648, N5649, N5650, N5651, N5652, N5653, N5654, N5655,
         N5656, N5657, N5675, N5676, N5677, N5678, N5679, N5680, N5681, N5682,
         N5683, N5684, N5685, N5686, N5687, N5688, N5689, N5690, N5691, N5692,
         N5693, N5694, N5695, N5721, N5722, N5723, N5724, N5725, N5726, N5727,
         N5728, N5729, N5730, N5731, N5732, N5733, N5734, N5735, N5736, N5754,
         N5755, N5756, N5757, N5758, N5759, N5760, N5761, N5762, N5763, N5764,
         N5765, N5766, N5767, N5768, N5769, N5770, N5771, N5772, N5773, N5774,
         N5810, N5811, N5812, N5813, N5814, N5815, N5816, N5817, N5818, N5819,
         N5820, N5821, N5822, N5823, N5824, N5825, N5843, N5844, N5845, N5846,
         N5847, N5848, N5849, N5850, N5851, N5852, N5853, N5854, N5855, N5856,
         N5857, N5858, N5859, N5860, N5861, N5862, N5863, N5888, N5892, N5893,
         N5894, N5895, N5896, N5897, N5898, N5899, N5900, N5901, N5902, N5903,
         N5904, N5905, N5906, N5907, N5925, N5926, N5927, N5928, N5929, N5930,
         N5931, N5932, N5933, N5934, N5935, N5936, N5937, N5938, N5939, N5940,
         N5941, N5942, N5943, N5944, N5945, N5981, N5982, N5983, N5984, N5985,
         N5986, N5987, N5988, N5989, N5990, N5991, N5992, N5993, N5994, N5995,
         N5996, N6014, N6015, N6016, N6017, N6018, N6019, N6020, N6021, N6022,
         N6023, N6024, N6025, N6026, N6027, N6028, N6029, N6030, N6031, N6032,
         N6033, N6034, N6060, N6061, N6062, N6063, N6064, N6065, N6066, N6067,
         N6068, N6069, N6070, N6071, N6072, N6073, N6074, N6075, N6093, N6094,
         N6095, N6096, N6097, N6098, N6099, N6100, N6101, N6102, N6103, N6104,
         N6105, N6106, N6107, N6108, N6109, N6110, N6111, N6112, N6113, N6149,
         N6150, N6151, N6152, N6153, N6154, N6155, N6156, N6157, N6158, N6159,
         N6160, N6161, N6162, N6163, N6164, N6182, N6183, N6184, N6185, N6186,
         N6187, N6188, N6189, N6190, N6191, N6192, N6193, N6194, N6195, N6196,
         N6197, N6198, N6199, N6200, N6201, N6202, N6228, N6229, N6230, N6231,
         N6232, N6233, N6234, N6235, N6236, N6237, N6238, N6239, N6240, N6241,
         N6242, N6243, N6261, N6262, N6263, N6264, N6265, N6266, N6267, N6268,
         N6269, N6270, N6271, N6272, N6273, N6274, N6275, N6276, N6277, N6278,
         N6279, N6280, N6281, N6317, N6318, N6319, N6320, N6321, N6322, N6323,
         N6324, N6325, N6326, N6327, N6328, N6329, N6330, N6331, N6332, N6350,
         N6351, N6352, N6353, N6354, N6355, N6356, N6357, N6358, N6359, N6360,
         N6361, N6362, N6363, N6364, N6365, N6366, N6367, N6368, N6369, N6370,
         N6396, N6397, N6398, N6399, N6400, N6401, N6402, N6403, N6404, N6405,
         N6406, N6407, N6408, N6409, N6410, N6411, N6429, N6430, N6431, N6432,
         N6433, N6434, N6435, N6436, N6437, N6438, N6439, N6440, N6441, N6442,
         N6443, N6444, N6445, N6446, N6447, N6448, N6449, N6485, N6486, N6487,
         N6488, N6489, N6490, N6491, N6492, N6493, N6494, N6495, N6496, N6497,
         N6498, N6499, N6500, N6518, N6519, N6520, N6521, N6522, N6523, N6524,
         N6525, N6526, N6527, N6528, N6529, N6530, N6531, N6532, N6533, N6534,
         N6535, N6536, N6537, N6538, N6563, N6567, N6568, N6569, N6570, N6571,
         N6572, N6573, N6574, N6575, N6576, N6577, N6578, N6579, N6580, N6581,
         N6582, N6600, N6601, N6602, N6603, N6604, N6605, N6606, N6607, N6608,
         N6609, N6610, N6611, N6612, N6613, N6614, N6615, N6616, N6617, N6618,
         N6619, N6620, N6667, N6668, N6669, N6670, N6671, N6672, N6673, N6674,
         N6675, N6676, N6677, N6678, N6679, N6680, N6681, N6682, N6700, N6701,
         N6702, N6703, N6704, N6705, N6706, N6707, N6708, N6709, N6710, N6711,
         N6712, N6713, N6714, N6715, N6716, N6717, N6718, N6719, N6720, N6749,
         N6750, N6751, N6752, N6753, N6754, N6755, N6756, N6757, N6758, N6759,
         N6760, N6761, N6762, N6763, N6764, N6782, N6783, N6784, N6785, N6786,
         N6787, N6788, N6789, N6790, N6791, N6792, N6793, N6794, N6795, N6796,
         N6797, N6798, N6799, N6800, N6801, N6802, N6841, N6842, N6843, N6844,
         N6845, N6846, N6847, N6848, N6849, N6850, N6851, N6852, N6853, N6854,
         N6855, N6856, N6874, N6875, N6876, N6877, N6878, N6879, N6880, N6881,
         N6882, N6883, N6884, N6885, N6886, N6887, N6888, N6889, N6890, N6891,
         N6892, N6893, N6894, N6923, N6924, N6925, N6926, N6927, N6928, N6929,
         N6930, N6931, N6932, N6933, N6934, N6935, N6936, N6937, N6938, N6956,
         N6957, N6958, N6959, N6960, N6961, N6962, N6963, N6964, N6965, N6966,
         N6967, N6968, N6969, N6970, N6971, N6972, N6973, N6974, N6975, N6976,
         N7015, N7016, N7017, N7018, N7019, N7020, N7021, N7022, N7023, N7024,
         N7025, N7026, N7027, N7028, N7029, N7030, N7048, N7049, N7050, N7051,
         N7052, N7053, N7054, N7055, N7056, N7057, N7058, N7059, N7060, N7061,
         N7062, N7063, N7064, N7065, N7066, N7067, N7068, N7097, N7098, N7099,
         N7100, N7101, N7102, N7103, N7104, N7105, N7106, N7107, N7108, N7109,
         N7110, N7111, N7112, N7130, N7131, N7132, N7133, N7134, N7135, N7136,
         N7137, N7138, N7139, N7140, N7141, N7142, N7143, N7144, N7145, N7146,
         N7147, N7148, N7149, N7150, N7189, N7190, N7191, N7192, N7193, N7194,
         N7195, N7196, N7197, N7198, N7199, N7200, N7201, N7202, N7203, N7204,
         N7222, N7223, N7224, N7225, N7226, N7227, N7228, N7229, N7230, N7231,
         N7232, N7233, N7234, N7235, N7236, N7237, N7238, N7239, N7240, N7241,
         N7242, N7267, N7271, N7272, N7273, N7274, N7275, N7276, N7277, N7278,
         N7279, N7280, N7281, N7282, N7283, N7284, N7285, N7286, N7304, N7305,
         N7306, N7307, N7308, N7309, N7310, N7311, N7312, N7313, N7314, N7315,
         N7316, N7317, N7318, N7319, N7320, N7321, N7322, N7323, N7324, N7360,
         N7361, N7362, N7363, N7364, N7365, N7366, N7367, N7368, N7369, N7370,
         N7371, N7372, N7373, N7374, N7375, N7393, N7394, N7395, N7396, N7397,
         N7398, N7399, N7400, N7401, N7402, N7403, N7404, N7405, N7406, N7407,
         N7408, N7409, N7410, N7411, N7412, N7413, N7439, N7440, N7441, N7442,
         N7443, N7444, N7445, N7446, N7447, N7448, N7449, N7450, N7451, N7452,
         N7453, N7454, N7472, N7473, N7474, N7475, N7476, N7477, N7478, N7479,
         N7480, N7481, N7482, N7483, N7484, N7485, N7486, N7487, N7488, N7489,
         N7490, N7491, N7492, N7528, N7529, N7530, N7531, N7532, N7533, N7534,
         N7535, N7536, N7537, N7538, N7539, N7540, N7541, N7542, N7543, N7561,
         N7562, N7563, N7564, N7565, N7566, N7567, N7568, N7569, N7570, N7571,
         N7572, N7573, N7574, N7575, N7576, N7577, N7578, N7579, N7580, N7581,
         N7607, N7608, N7609, N7610, N7611, N7612, N7613, N7614, N7615, N7616,
         N7617, N7618, N7619, N7620, N7621, N7622, N7640, N7641, N7642, N7643,
         N7644, N7645, N7646, N7647, N7648, N7649, N7650, N7651, N7652, N7653,
         N7654, N7655, N7656, N7657, N7658, N7659, N7660, N7696, N7697, N7698,
         N7699, N7700, N7701, N7702, N7703, N7704, N7705, N7706, N7707, N7708,
         N7709, N7710, N7711, N7729, N7730, N7731, N7732, N7733, N7734, N7735,
         N7736, N7737, N7738, N7739, N7740, N7741, N7742, N7743, N7744, N7745,
         N7746, N7747, N7748, N7749, N7775, N7776, N7777, N7778, N7779, N7780,
         N7781, N7782, N7783, N7784, N7785, N7786, N7787, N7788, N7789, N7790,
         N7808, N7809, N7810, N7811, N7812, N7813, N7814, N7815, N7816, N7817,
         N7818, N7819, N7820, N7821, N7822, N7823, N7824, N7825, N7826, N7827,
         N7828, N7864, N7865, N7866, N7867, N7868, N7869, N7870, N7871, N7872,
         N7873, N7874, N7875, N7876, N7877, N7878, N7879, N7897, N7898, N7899,
         N7900, N7901, N7902, N7903, N7904, N7905, N7906, N7907, N7908, N7909,
         N7910, N7911, N7912, N7913, N7914, N7915, N7916, N7917, N7942, N7946,
         N7947, N7948, N7949, N7950, N7951, N7952, N7953, N7954, N7955, N7956,
         N7957, N7958, N7959, N7960, N7961, N7979, N7980, N7981, N7982, N7983,
         N7984, N7985, N7986, N7987, N7988, N7989, N7990, N7991, N7992, N7993,
         N7994, N7995, N7996, N7997, N7998, N7999, n949, n950, n951, n952,
         n953, n954, n955, n956, n957, n958, n959, n960, n961, n962, n963,
         n964, n965, n966, n967, n968, n969, n970, n971, n972, n973, n974,
         n975, n976, n977, n978, n979, n980, n981, n982, n983, n984, n985,
         n986, n987, n988, n989, n990, n991, n992, n993, n994, n995, n996,
         n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006,
         n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016,
         n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026,
         n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036,
         n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046,
         n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056,
         n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066,
         n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076,
         n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086,
         n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096,
         n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106,
         n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116,
         n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196,
         n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206,
         n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216,
         n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226,
         n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236,
         n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246,
         n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256,
         n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266,
         n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276,
         n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286,
         n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296,
         n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306,
         n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316,
         n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326,
         n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336,
         n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346,
         n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356,
         n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366,
         n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376,
         n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386,
         n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396,
         n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406,
         n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416,
         n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426,
         n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436,
         n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446,
         n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456,
         n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586,
         n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596,
         n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606,
         n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616,
         n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626,
         n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636,
         n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646,
         n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656,
         n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666,
         n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676,
         n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686,
         n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696,
         n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706,
         n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716,
         n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726,
         n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736,
         n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746,
         n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756,
         n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766,
         n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776,
         n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786,
         n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796,
         n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806,
         n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816,
         n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826,
         n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836,
         n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846,
         n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856,
         n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866,
         n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876,
         n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886,
         n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896,
         n1897, n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906,
         n1907, n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916,
         n1917, n1918, n1919, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440,
         n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450,
         n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460,
         n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470,
         n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480,
         n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490,
         n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500,
         n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510,
         n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520,
         n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530,
         n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540,
         n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550,
         n2551, n2552, n255900, n256000, n256100, n256200, n256300, n256400,
         n256500, n256600, n256700, n256800, n256900, n257000, n257100,
         n257200, n257300, n257400, n2575, n2576, n2577, n2578, n2579, n2580,
         n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590,
         n2591, n259200, n259300, n259400, n259500, n259600, n259700, n259800,
         n259900, n260000, n260100, n260200, n260300, n260400, n260500,
         n260600, n260700, n260800, n260900, n261000, n261100, n261200, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n263700, n2638, n2639, n2640, n264100, n264200,
         n264300, n264400, n264500, n264600, n264700, n264800, n265500,
         n265600, n2657, n2658, n2659, n2660, n2661, n2662, n2663, n2664,
         n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n267400, n267500, n267600, n267700, n267800, n267900, n268000,
         n268100, n268200, n268300, n268400, n269100, n269200, n269300,
         n269400, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n272900, n2730, n2731,
         n2732, n273300, n273400, n273500, n273600, n273700, n273800, n273900,
         n274000, n274100, n274200, n274300, n274400, n274500, n274600,
         n274700, n274800, n2749, n2750, n2751, n2752, n2753, n2754, n2755,
         n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765,
         n276600, n276700, n276800, n276900, n277000, n277100, n277200,
         n277300, n277400, n277500, n277600, n277700, n277800, n277900,
         n278000, n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794,
         n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804,
         n2805, n2806, n2807, n2808, n2809, n2810, n28110, n2812, n2813, n2814,
         n28150, n28160, n28230, n28240, n28250, n28260, n28270, n28280,
         n28290, n28300, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n28480, n28490, n28500, n28510, n28520, n28530, n28540, n28550,
         n28560, n28570, n28580, n28590, n28600, n28610, n28620, n28630,
         n28640, n28650, n28660, n28670, n28680, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n3070, n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080,
         n30810, n30820, n30830, n30840, n30850, n30860, n30870, n30880,
         n30890, n30900, n30910, n30920, n30930, n30940, n30950, n3097, n3098,
         n3099, n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3112,
         n3113, n31140, n31150, n31160, n31170, n31180, n31190, n31200, n31210,
         n31220, n31230, n31240, n31250, n31260, n31270, n31280, n31290,
         n31300, n31310, n31320, n31330, n31340, n3135, n3137, n3138, n3139,
         n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149,
         n3150, n3151, n3152, n3154, n3155, n3156, n3157, n3158, n3159, n3160,
         n3161, n3162, n31630, n31640, n31650, n31660, n31670, n31680, n31690,
         n31700, n31710, n31720, n31730, n31740, n31750, n31760, n31770,
         n31780, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n31960,
         n31970, n31980, n31990, n32000, n32010, n32020, n32040, n32050,
         n32060, n32070, n32080, n32090, n32110, n32120, n32130, n32140,
         n32150, n32160, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3229, n3230, n3231, n3232, n3233, n3234,
         n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245,
         n3246, n3247, n3248, n3249, n3250, n3251, n32520, n32540, n32550,
         n32560, n32570, n32580, n32590, n32600, n32620, n32630, n32640,
         n32650, n32660, n32670, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n32850, n32860, n32870, n32880, n32890, n32900, n32910, n32920,
         n32930, n32940, n32950, n32960, n32970, n32980, n32990, n33000,
         n33020, n33030, n33040, n33050, n3306, n3307, n3308, n3309, n3310,
         n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320,
         n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330,
         n33310, n33320, n33330, n33340, n33350, n33360, n33370, n33380,
         n33390, n33400, n33410, n33420, n33430, n33440, n33450, n33460, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n33640, n33650, n33660,
         n33670, n33680, n33690, n33700, n33710, n33720, n33730, n33740,
         n33750, n33760, n33770, n33780, n33790, n33800, n33810, n33820,
         n33830, n33840, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n34200,
         n34210, n34220, n34230, n34240, n34250, n34260, n34270, n34280,
         n34290, n34300, n34310, n34320, n34330, n34340, n3436, n3437, n3438,
         n3439, n3440, n3441, n3443, n3444, n3445, n3446, n3447, n3448, n3449,
         n3450, n3451, n3452, n34530, n34540, n34550, n34560, n34570, n34580,
         n34590, n34600, n34610, n34620, n34630, n34640, n34650, n34660,
         n34670, n34680, n34690, n34700, n34710, n34720, n34730, n3474, n3475,
         n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485,
         n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495,
         n3496, n3497, n3498, n34990, n35000, n35010, n35020, n35030, n35040,
         n35050, n35060, n35070, n35080, n35090, n35100, n35110, n35120,
         n35130, n35140, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n35320, n35330, n35340, n35350, n35360, n35370, n35380, n35390,
         n35400, n35410, n35420, n35430, n35440, n35450, n35460, n35470,
         n35480, n35490, n35500, n35510, n35520, n3553, n3554, n3555, n3556,
         n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566,
         n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576,
         n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586,
         n3587, n35880, n35890, n35900, n35910, n35920, n35930, n35940, n35950,
         n35960, n35970, n35980, n35990, n36000, n36010, n36020, n36030, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3618, n3619, n3620, n36210, n36220, n36230, n36250,
         n36260, n36270, n36280, n36290, n36300, n36310, n36320, n36330,
         n36340, n36350, n36360, n36370, n36380, n36390, n36400, n36410, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n36670, n36680, n36690, n36700, n36710,
         n36720, n36730, n36740, n36750, n36760, n36770, n36780, n36790,
         n36800, n36810, n36820, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n37000, n37010, n37020, n37030, n37040, n37050, n37060, n37070,
         n37080, n37090, n37100, n37110, n37120, n37130, n37140, n37150,
         n37160, n37170, n37180, n37190, n37200, n3721, n3722, n3723, n3724,
         n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734,
         n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744,
         n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754,
         n3755, n37560, n37570, n37580, n37590, n37600, n37610, n37620, n37630,
         n37640, n37650, n37660, n37670, n37680, n37690, n37700, n37710, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n37890, n37900, n37910,
         n37920, n37930, n37940, n37950, n37960, n37970, n37980, n37990,
         n38000, n38010, n38020, n38030, n38040, n38050, n38060, n38070,
         n38080, n38090, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n38380, n38390, n38400, n38410, n38420, n38430, n38440, n38450,
         n38470, n38480, n38490, n38500, n38510, n38520, n38530, n3854, n3855,
         n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865,
         n3866, n3867, n3868, n3869, n3870, n38710, n38720, n38730, n38740,
         n38750, n38760, n38770, n38780, n38790, n38800, n38810, n38820,
         n38830, n38840, n38850, n38860, n38870, n38880, n38890, n38900,
         n38910, n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900,
         n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910,
         n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920,
         n3921, n3922, n3923, n3924, n3925, n3926, n39270, n39280, n39290,
         n39300, n39310, n39320, n39330, n39340, n39350, n39360, n39370,
         n39380, n39390, n39400, n39410, n39420, n3943, n3944, n3945, n3946,
         n3947, n3948, n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956,
         n3957, n3958, n3959, n39600, n39610, n39620, n39630, n39640, n39650,
         n39660, n39670, n39680, n39690, n39700, n39710, n39720, n39730,
         n39740, n39750, n39760, n39770, n39780, n39790, n39800, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n40060, n40070, n40080, n40090, n40100, n40110,
         n40120, n40130, n40140, n40150, n40160, n40170, n40180, n40190,
         n40200, n40210, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n40390, n40400, n40410, n40420, n40430, n40440, n40450, n40460,
         n40470, n40480, n40490, n40500, n40510, n40520, n40530, n40540,
         n40550, n40560, n40570, n40580, n40590, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n40950, n40960, n40970, n40980, n40990, n41000, n41010, n41020,
         n41030, n41040, n41050, n41060, n41070, n41080, n41090, n41100, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n41280, n41290, n41300,
         n41310, n41320, n41330, n41340, n41350, n41360, n41370, n41380,
         n41390, n41400, n41410, n41420, n41430, n41440, n41450, n41460,
         n41470, n41480, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4172, n4173, n41740, n41750,
         n41760, n41770, n41780, n41790, n41800, n41810, n41820, n41830,
         n41840, n41850, n41860, n41870, n41880, n41890, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n42070, n42080, n42090, n42100, n42110,
         n42120, n42130, n42140, n42150, n42160, n42170, n42180, n42190,
         n42200, n42210, n42220, n42230, n42240, n42250, n42260, n42270, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n42630, n42640, n42650, n42660, n42670,
         n42680, n42690, n42700, n42710, n42720, n42730, n42740, n42750,
         n42760, n42770, n42780, n4279, n4280, n4281, n4282, n4283, n4284,
         n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294,
         n4295, n42960, n42970, n42980, n42990, n43000, n43010, n43020, n43030,
         n43040, n43050, n43060, n43070, n43080, n43090, n43100, n43110,
         n43120, n43130, n43140, n43150, n43160, n4317, n4318, n4319, n4320,
         n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330,
         n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340,
         n4341, n43420, n43430, n43440, n43450, n43460, n43470, n43480, n43490,
         n43500, n43510, n43520, n43550, n43560, n43570, n4358, n4359, n4360,
         n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370,
         n4371, n4372, n4373, n4374, n43750, n43760, n43770, n43780, n43790,
         n43800, n43810, n43820, n43830, n43840, n43850, n43860, n43870,
         n43880, n43890, n43900, n43910, n43920, n43930, n43950, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n44310, n44320, n44330, n44340, n44350, n44360,
         n44370, n44380, n44390, n44400, n44410, n44420, n44430, n44440,
         n44450, n44460, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n44640, n44650, n44660, n44670, n44680, n44690, n44700, n44710,
         n44720, n44730, n44740, n44750, n44760, n44770, n44780, n44790,
         n44800, n44810, n44820, n44830, n44840, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n45090, n4510, n4511, n4512, n45130, n45140, n45150, n45160, n45170,
         n45180, n45190, n45200, n45210, n45220, n45230, n45240, n45250,
         n45260, n45270, n45280, n4529, n4530, n4531, n4532, n4533, n4534,
         n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544,
         n4545, n45460, n45470, n45480, n45490, n45500, n45510, n45520, n45530,
         n45540, n45550, n45560, n45570, n45580, n45590, n45600, n45610,
         n45620, n45630, n45640, n45650, n45660, n4567, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n46130, n46140, n46150, n46160, n46170, n46180, n46190, n46200,
         n46210, n46220, n46230, n46240, n46250, n46260, n46270, n46280, n4629,
         n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639,
         n4640, n4641, n4642, n4643, n4644, n4645, n46460, n46470, n46480,
         n46490, n46500, n46510, n46520, n46530, n46540, n46550, n46560,
         n46570, n46580, n46590, n46600, n46610, n46620, n46630, n46640,
         n46650, n46660, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n46950, n46960, n46970, n46980, n46990, n47000, n47010, n47020,
         n47040, n47050, n47060, n47090, n47100, n4711, n4712, n4713, n4714,
         n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4723, n4724, n4725,
         n4726, n4727, n47280, n47290, n47300, n47310, n47320, n47330, n47340,
         n47350, n47360, n47370, n47380, n47390, n47400, n47410, n47420,
         n47430, n47440, n47450, n47460, n47470, n47480, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n47880, n47890, n47900, n47910,
         n47920, n47930, n47940, n47950, n47960, n47970, n47980, n47990,
         n48000, n48010, n48020, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n48200, n48210, n48220, n48230, n48240, n48250, n48260, n48270,
         n48280, n48290, n48300, n48310, n48320, n48330, n48340, n48350,
         n48360, n48370, n48380, n48390, n48400, n4841, n4842, n4843, n4844,
         n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854,
         n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864,
         n4865, n4866, n4867, n4868, n48690, n48700, n48710, n48720, n48730,
         n48740, n48750, n48760, n48770, n48780, n48790, n48810, n48820,
         n48830, n48840, n4885, n4886, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n49020,
         n49030, n49040, n49050, n49060, n49070, n49080, n49090, n49100,
         n49110, n49120, n49130, n49140, n49150, n49160, n49170, n49180,
         n49190, n49200, n49210, n49220, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n49610, n49620, n49630, n49640, n49650, n49660,
         n49670, n49680, n49690, n49700, n49710, n49720, n49730, n49740,
         n49750, n49760, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n49940, n49950, n49960, n49970, n49980, n49990, n50000, n50010,
         n50020, n50030, n50040, n50050, n50060, n50070, n50080, n50090,
         n50100, n50110, n50120, n50130, n50140, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n50430, n50440, n50450, n50460, n50470,
         n50480, n50490, n50500, n50510, n50520, n50530, n50540, n50550,
         n50560, n50570, n50580, n5059, n5060, n5061, n5062, n5063, n5064,
         n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074,
         n5075, n50760, n50770, n50780, n50800, n50810, n50820, n50830, n50840,
         n50850, n50860, n50870, n50880, n50890, n50900, n50910, n50920,
         n50930, n50940, n50950, n50960, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n51360, n51370, n51380, n51390, n51400, n51410, n51420,
         n51430, n51440, n51450, n51460, n51470, n51480, n51490, n51500, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n51680, n51690, n51700,
         n51710, n51720, n51730, n51740, n51750, n51760, n51770, n51780,
         n51790, n51800, n51810, n51820, n51830, n51840, n51850, n51860,
         n51870, n51880, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5202, n5203, n5204, n5205, n5206,
         n5207, n5208, n5209, n5210, n5211, n5212, n52130, n5214, n5215, n5216,
         n52170, n52180, n52190, n52200, n52210, n52220, n52230, n52240,
         n52250, n52260, n52270, n52280, n52290, n52300, n52310, n52320, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n52500, n52510, n52520,
         n52530, n52540, n52550, n52560, n52570, n52580, n52590, n52600,
         n52610, n52620, n52630, n52640, n52650, n52660, n52670, n52680,
         n52690, n52700, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n53060, n53070,
         n53080, n53090, n53100, n53110, n53120, n53130, n53140, n53150,
         n53160, n53170, n53180, n53190, n53200, n53210, n5322, n5323, n5324,
         n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334,
         n5335, n5336, n5337, n5338, n53390, n53400, n53410, n53420, n53430,
         n53440, n53450, n53460, n53470, n53480, n53490, n53500, n53510,
         n53520, n53530, n53540, n53550, n53560, n53570, n53580, n53590, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n53850, n53860, n53870, n53880, n53890,
         n53900, n53910, n53920, n53930, n53940, n53950, n53960, n53970,
         n53980, n53990, n54000, n5401, n5402, n5403, n5404, n5405, n5406,
         n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n54180,
         n54190, n54200, n54210, n54220, n54230, n54240, n54250, n54260,
         n54270, n54280, n54290, n54300, n54310, n54320, n54330, n54340,
         n54350, n54360, n54370, n54380, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n54740, n54750, n54760, n54770, n54780, n54790, n54800, n54810,
         n54820, n54830, n54840, n54850, n54860, n54870, n54880, n54890, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n55070, n55080, n55090,
         n55100, n55110, n55120, n55130, n55140, n55150, n55160, n55170,
         n55180, n55190, n55200, n55210, n55220, n55230, n55240, n55250,
         n55260, n55270, n5528, n5529, n5530, n5531, n5532, n5533, n5534,
         n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544,
         n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n55530,
         n55540, n55550, n55560, n55570, n55580, n55590, n55600, n55610,
         n55620, n55630, n55640, n55650, n55660, n55670, n55680, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n55860, n55870, n55880, n55890,
         n55900, n55910, n55920, n55930, n55940, n55950, n55960, n55970,
         n55980, n55990, n56000, n56010, n56020, n56030, n56040, n56050,
         n56060, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n56420, n56430, n56440,
         n56450, n56460, n56470, n56480, n56490, n56500, n56510, n56520,
         n56530, n56540, n56550, n56560, n56570, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n56750, n56760, n56770, n56780, n56790, n56800,
         n56810, n56820, n56830, n56840, n56850, n56860, n56870, n56880,
         n56890, n56900, n56910, n56920, n56930, n56940, n56950, n5696, n5697,
         n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707,
         n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717,
         n5718, n5719, n5720, n57210, n57220, n57230, n57240, n57250, n57260,
         n57270, n57280, n57290, n57300, n57310, n57320, n57330, n57340,
         n57350, n57360, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n57540, n57550, n57560, n57570, n57580, n57590, n57600, n57610,
         n57620, n57630, n57640, n57650, n57660, n57670, n57680, n57690,
         n57700, n57710, n57720, n57730, n57740, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n58100, n58110, n58120, n58130, n58140, n58150, n58160, n58170,
         n58180, n58190, n58200, n58210, n58220, n58230, n58240, n58250, n5826,
         n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836,
         n5837, n5838, n5839, n5840, n5841, n5842, n58430, n58440, n58450,
         n58460, n58470, n58480, n58490, n58500, n58510, n58520, n58530,
         n58540, n58550, n58560, n58570, n58580, n58590, n58600, n58610,
         n58620, n58630, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n58880, n5889, n5890,
         n5891, n58920, n58930, n58940, n58950, n58960, n58970, n58980, n58990,
         n59000, n59010, n59020, n59030, n59040, n59050, n59060, n59070, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n59250, n59260, n59270,
         n59280, n59290, n59300, n59310, n59320, n59330, n59340, n59350,
         n59360, n59370, n59380, n59390, n59400, n59410, n59420, n59430,
         n59440, n59450, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n59810,
         n59820, n59830, n59840, n59850, n59860, n59870, n59880, n59890,
         n59900, n59910, n59920, n59930, n59940, n59950, n59960, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n60140, n60150, n60160, n60170,
         n60180, n60190, n60200, n60210, n60220, n60230, n60240, n60250,
         n60260, n60270, n60280, n60290, n60300, n60310, n60320, n60330,
         n60340, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n60600, n60610, n60620,
         n60630, n60640, n60650, n60660, n60670, n60680, n60690, n60700,
         n60710, n60720, n60730, n60740, n60750, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n60930, n60940, n60950, n60960, n60970, n60980,
         n60990, n61000, n61010, n61020, n61030, n61040, n61050, n61060,
         n61070, n61080, n61090, n61100, n61110, n61120, n61130, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n61490, n61500, n61510, n61520, n61530, n61540,
         n61550, n61560, n61570, n61580, n61590, n61600, n61610, n61620,
         n61630, n61640, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n61820, n61830, n61840, n61850, n61860, n61870, n61880, n61890,
         n61900, n61910, n61920, n61930, n61940, n61950, n61960, n61970,
         n61980, n61990, n62000, n62010, n62020, n6203, n6204, n6205, n6206,
         n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216,
         n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226,
         n6227, n62280, n62290, n62300, n62310, n62320, n62330, n62340, n62350,
         n62360, n62370, n62380, n62390, n62400, n62410, n62420, n62430, n6244,
         n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254,
         n6255, n6256, n6257, n6258, n6259, n6260, n62610, n62620, n62630,
         n62640, n62650, n62660, n62670, n62680, n62690, n62700, n62710,
         n62720, n62730, n62740, n62750, n62760, n62770, n62780, n62790,
         n62800, n62810, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n63170,
         n63180, n63190, n63200, n63210, n63220, n63230, n63240, n63250,
         n63260, n63270, n63280, n63290, n63300, n63310, n63320, n6333, n6334,
         n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344,
         n6345, n6346, n6347, n6348, n6349, n63500, n63510, n63520, n63530,
         n63540, n63550, n63560, n63570, n63580, n63590, n63600, n63610,
         n63620, n63630, n63640, n63650, n63660, n63670, n63680, n63690,
         n63700, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n63960, n63970, n63980,
         n63990, n64000, n64010, n64020, n64030, n64040, n64050, n64060,
         n64070, n64080, n64090, n64100, n64110, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n64290, n64300, n64310, n64320, n64330, n64340,
         n64350, n64360, n64370, n64380, n64390, n64400, n64410, n64420,
         n64430, n64440, n64450, n64460, n64470, n64480, n64490, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n64850, n64860, n64870, n64880, n64890, n64900,
         n64910, n64920, n64930, n64940, n64950, n64960, n64970, n64980,
         n64990, n65000, n6501, n6502, n6503, n6504, n6505, n6506, n6507,
         n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517,
         n65180, n65190, n65200, n65210, n65220, n65230, n65240, n65250,
         n65260, n65270, n65280, n65290, n65300, n65310, n65320, n65330,
         n65340, n65350, n65360, n65370, n65380, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n65630, n6564, n6565, n6566, n65670, n65680, n65690, n65700, n65710,
         n65720, n65730, n65740, n65750, n65760, n65770, n65780, n65790,
         n65800, n65810, n65820, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n66000, n66010, n66020, n66030, n66040, n66050, n66060, n66070,
         n66080, n66090, n66100, n66110, n66120, n66130, n66140, n66150,
         n66160, n66170, n66180, n66190, n66200, n6621, n6622, n6623, n6624,
         n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634,
         n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644,
         n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654,
         n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664,
         n6665, n6666, n66670, n66680, n66690, n66700, n66710, n66720, n66730,
         n66740, n66750, n66760, n66770, n66780, n66790, n66800, n66810,
         n66820, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n67000,
         n67010, n67020, n67030, n67040, n67050, n67060, n67070, n67080,
         n67090, n67100, n67110, n67120, n67130, n67140, n67150, n67160,
         n67170, n67180, n67190, n67200, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n67490, n67500, n67510, n67520, n67530, n67540,
         n67550, n67560, n67570, n67580, n67590, n67600, n67610, n67620,
         n67630, n67640, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n67820, n67830, n67840, n67850, n67860, n67870, n67880, n67890,
         n67900, n67910, n67920, n67930, n67940, n67950, n67960, n67970,
         n67980, n67990, n68000, n68010, n68020, n6803, n6804, n6805, n6806,
         n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816,
         n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826,
         n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836,
         n6837, n6838, n6839, n6840, n68410, n68420, n68430, n68440, n68450,
         n68460, n68470, n68480, n68490, n68500, n68510, n68520, n68530,
         n68540, n68550, n68560, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n68740, n68750, n68760, n68770, n68780, n68790, n68800, n68810,
         n68820, n68830, n68840, n68850, n68860, n68870, n68880, n68890,
         n68900, n68910, n68920, n68930, n68940, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n69230, n69240, n69250, n69260, n69270,
         n69280, n69290, n69300, n69310, n69320, n69330, n69340, n69350,
         n69360, n69370, n69380, n6939, n6940, n6941, n6942, n6943, n6944,
         n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954,
         n6955, n69560, n69570, n69580, n69590, n69600, n69610, n69620, n69630,
         n69640, n69650, n69660, n69670, n69680, n69690, n69700, n69710,
         n69720, n69730, n69740, n69750, n69760, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n70150, n70160, n70170, n70180, n70190,
         n70200, n70210, n70220, n70230, n70240, n70250, n70260, n70270,
         n70280, n70290, n70300, n7031, n7032, n7033, n7034, n7035, n7036,
         n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046,
         n7047, n70480, n70490, n70500, n70510, n70520, n70530, n70540, n70550,
         n70560, n70570, n70580, n70590, n70600, n70610, n70620, n70630,
         n70640, n70650, n70660, n70670, n70680, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n70970, n70980, n70990, n71000, n71010,
         n71020, n71030, n71040, n71050, n71060, n71070, n71080, n71090,
         n71100, n71110, n71120, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n71300, n71310, n71320, n71330, n71340, n71350, n71360, n71370,
         n71380, n71390, n71400, n71410, n71420, n71430, n71440, n71450,
         n71460, n71470, n71480, n71490, n71500, n7151, n7152, n7153, n7154,
         n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164,
         n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174,
         n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184,
         n7185, n7186, n7187, n7188, n71890, n71900, n71910, n71920, n71930,
         n71940, n71950, n71960, n71970, n71980, n71990, n72000, n72010,
         n72020, n72030, n72040, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n72220, n72230, n72240, n72250, n72260, n72270, n72280, n72290,
         n72300, n72310, n72320, n72330, n72340, n72350, n72360, n72370,
         n72380, n72390, n72400, n72410, n72420, n7243, n7244, n7245, n7246,
         n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256,
         n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266,
         n72670, n7268, n7269, n7270, n72710, n72720, n72730, n72740, n72750,
         n72760, n72770, n72780, n72790, n72800, n72810, n72820, n72830,
         n72840, n72850, n72860, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n73040, n73050, n73060, n73070, n73080, n73090, n73100, n73110,
         n73120, n73130, n73140, n73150, n73160, n73170, n73180, n73190,
         n73200, n73210, n73220, n73230, n73240, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n73600, n73610, n73620, n73630, n73640, n73650, n73660, n73670,
         n73680, n73690, n73700, n73710, n73720, n73730, n73740, n73750, n7376,
         n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386,
         n7387, n7388, n7389, n7390, n7391, n7392, n73930, n73940, n73950,
         n73960, n73970, n73980, n73990, n74000, n74010, n74020, n74030,
         n74040, n74050, n74060, n74070, n74080, n74090, r899_B_1_, r899_B_2_,
         r899_B_3_, r899_B_4_, r899_B_6_, r899_B_7_, r899_B_9_, r924_LT_LE,
         r929_LT_LE, r948_LT_LE, add_124_aco_B_3_, n1, n2, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n1920, n1921, n1922, n1923, n1924, n1925, n2205, n2206,
         n2207, n2208, n2209, n2210, n2286, n2287, n2288, n2289, n2290, n2291,
         n2427, n2428, n2429, n2430, n2431, n2432, n2553, n2554, n2555, n2556,
         n2557, n2558, n264900, n265000, n265100, n265200, n265300, n265400,
         n268500, n268600, n268700, n268800, n268900, n269000, n278100,
         n278200, n278300, n278400, n278500, n278600, n28170, n28180, n28190,
         n28200, n28210, n28220, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n29030, n2904, n2905, n2906, n29070,
         n29080, n29090, n29100, n29110, n29120, n29130, n29140, n29150,
         n29160, n29170, n29180, n29190, n29200, n29210, n29220, n2923, n2924,
         n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934,
         n2935, n2936, n2937, n2938, n2939, n29400, n29410, n29420, n29430,
         n29440, n29450, n29460, n29470, n29480, n29490, n29500, n29510,
         n29520, n29530, n29540, n29550, n29560, n29570, n29580, n29590,
         n29600, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969,
         n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979,
         n2980, n2981, n2982, n2983, n2984, n29850, n2986, n2987, n2988,
         n29890, n29900, n29910, n29920, n29930, n29940, n29950, n29960,
         n29970, n29980, n29990, n30000, n30010, n30020, n30030, n30040, n3005,
         n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015,
         n3016, n3017, n3018, n3019, n3020, n3021, n30220, n30230, n30240,
         n30250, n30260, n30270, n30280, n30290, n30300, n30310, n30320,
         n30330, n30340, n30350, n30360, n30370, n30380, n30390, n30400,
         n30410, n30420, n3043, n3044, n3045, n3046, n3047, n3048, n3049,
         n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059,
         n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069,
         n3071, n30960, n3100, n3101, n3110, n3111, n3136, n3153, n32030,
         n32100, n3228, n3235, n32530, n32610, n33010, n34350, n3442, n3617,
         n36240, n38460, n4171, n43530, n43540, n43940, n4568, n47030, n47070,
         n47080, n4722, n47870, n48800, n4887, n4888, n50790, n5107, n51350,
         n5201, n5296, n5416, n5417, n74100, n74110, n74120, n74130, n7414,
         n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424,
         n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434,
         n7435, n7436, n7437, n7438, n74390, n74400, n74410, n74420, n74430,
         n74440, n74450, n74460, n74470, n74480, n74490, n74500, n74510,
         n74520, n74530, n74540, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n74720, n74730, n74740, n74750, n74760, n74770, n74780, n74790,
         n74800, n74810, n74820, n74830, n74840, n74850, n74860, n74870,
         n74880, n74890, n74900, n74910, n74920, n7493, n7494, n7495, n7496,
         n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506,
         n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516,
         n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526,
         n7527, n75280, n75290, n75300, n75310, n75320, n75330, n75340, n75350,
         n75360, n75370, n75380, n75390, n75400, n75410, n75420, n75430, n7544,
         n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554,
         n7555, n7556, n7557, n7558, n7559, n7560, n75610, n75620, n75630,
         n75640, n75650, n75660, n75670, n75680, n75690, n75700, n75710,
         n75720, n75730, n75740, n75750, n75760, n75770, n75780, n75790,
         n75800, n75810, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n76070,
         n76080, n76090, n76100, n76110, n76120, n76130, n76140, n76150,
         n76160, n76170, n76180, n76190, n76200, n76210, n76220, n7623, n7624,
         n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634,
         n7635, n7636, n7637, n7638, n7639, n76400, n76410, n76420, n76430,
         n76440, n76450, n76460, n76470, n76480, n76490, n76500, n76510,
         n76520, n76530, n76540, n76550, n76560, n76570, n76580, n76590,
         n76600, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n76960, n76970, n76980,
         n76990, n77000, n77010, n77020, n77030, n77040, n77050, n77060,
         n77070, n77080, n77090, n77100, n77110, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n77290, n77300, n77310, n77320, n77330, n77340,
         n77350, n77360, n77370, n77380, n77390, n77400, n77410, n77420,
         n77430, n77440, n77450, n77460, n77470, n77480, n77490, n7750, n7751,
         n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761,
         n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771,
         n7772, n7773, n7774, n77750, n77760, n77770, n77780, n77790, n77800,
         n77810, n77820, n77830, n77840, n77850, n77860, n77870, n77880,
         n77890, n77900, n7791, n7792, n7793, n7794, n7795, n7796, n7797,
         n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807,
         n78080, n78090, n78100, n78110, n78120, n78130, n78140, n78150,
         n78160, n78170, n78180, n78190, n78200, n78210, n78220, n78230,
         n78240, n78250, n78260, n78270, n78280, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n78640, n78650, n78660, n78670, n78680, n78690, n78700, n78710,
         n78720, n78730, n78740, n78750, n78760, n78770, n78780, n78790, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n78970, n78980, n78990,
         n79000, n79010, n79020, n79030, n79040, n79050, n79060, n79070,
         n79080, n79090, n79100, n79110, n79120, n79130, n79140, n79150,
         n79160, n79170, n7918, n7919, n7920, n7921, n7922, n7923, n7924,
         n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934,
         n7935, n7936, n7937, n7938, n7939, n7940, n7941, n79420, n7943, n7944,
         n7945, n79460, n79470, n79480, n79490, n79500, n79510, n79520, n79530,
         n79540, n79550, n79560, n79570, n79580, n79590, n79600, n79610, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n79790, n79800, n79810,
         n79820, n79830, n79840, n79850, n79860, n79870, n79880, n79890,
         n79900, n79910, n79920, n79930, n79940, n79950, n79960, n79970,
         n79980, n79990, n8000, n8001, n8002, n8003, n8004, n8005, n8006,
         n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016,
         n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026,
         n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036,
         n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046,
         n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056,
         n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066,
         n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076,
         n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086,
         n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096,
         n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106,
         n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116,
         n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126,
         n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136,
         n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146,
         n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156,
         n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166,
         n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176,
         n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186,
         n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196,
         n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206,
         n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216,
         n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226,
         n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236,
         n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246,
         n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256,
         n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266,
         n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276,
         n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286,
         n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296,
         n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306,
         n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316,
         n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326,
         n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336,
         n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346,
         n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356,
         n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366,
         n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376,
         n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386,
         n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396,
         n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406,
         n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416,
         n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426,
         n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436,
         n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446,
         n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456,
         n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466,
         n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476,
         n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486,
         n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496,
         n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506,
         n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516,
         n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526,
         n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536,
         n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546,
         n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556,
         n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566,
         n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576,
         n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586,
         n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596,
         n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606,
         n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616,
         n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626,
         n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636,
         n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646,
         n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656,
         n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666,
         n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676,
         n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686,
         n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696,
         n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706,
         n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716,
         n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726,
         n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736,
         n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746,
         n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756,
         n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766,
         n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776,
         n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786,
         n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796,
         n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806,
         n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816,
         n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826,
         n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836,
         n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846,
         n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856,
         n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866,
         n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876,
         n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886,
         n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896,
         n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906,
         n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916,
         n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926,
         n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936,
         n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946,
         n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956,
         n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966,
         n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976,
         n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986,
         n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996,
         n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006,
         n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016,
         n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026,
         n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036,
         n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046,
         n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056,
         n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066,
         n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076,
         n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086,
         n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096,
         n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106,
         n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116,
         n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126,
         n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136,
         n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146,
         n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156,
         n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166,
         n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176,
         n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186,
         n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196,
         n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206,
         n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216,
         n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226,
         n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236,
         n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246,
         n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256,
         n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266,
         n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276,
         n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286,
         n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296,
         n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306,
         n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316,
         n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326,
         n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336,
         n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346,
         n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356,
         n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366,
         n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376,
         n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386,
         n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396,
         n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406,
         n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416,
         n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426,
         n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436,
         n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446,
         n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456,
         n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466,
         n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476,
         n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486,
         n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496,
         n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506,
         n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516,
         n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526,
         n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536,
         n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546,
         n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556,
         n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566,
         n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576,
         n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586,
         n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596,
         n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606,
         n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616,
         n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626,
         n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636,
         n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646,
         n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656,
         n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666,
         n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676,
         n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686,
         n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696,
         n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706,
         n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716,
         n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726,
         n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736,
         n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746,
         n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756,
         n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766,
         n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776,
         n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786,
         n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796,
         n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806,
         n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816,
         n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826,
         n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836,
         n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846,
         n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856,
         n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866,
         n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876,
         n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886,
         n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896,
         n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906,
         n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916,
         n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926,
         n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936,
         n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946,
         n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956,
         n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966,
         n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976,
         n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986,
         n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996,
         n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004, n10005,
         n10006, n10007, n10008, n10009, n10010, n10011, n10012, n10013,
         n10014, n10015, n10016, n10017, n10018, n10019, n10020, n10021,
         n10022, n10023, n10024, n10025, n10026, n10027, n10028, n10029,
         n10030, n10031, n10032, n10033, n10034, n10035, n10036, n10037,
         n10038, n10039, n10040, n10041, n10042, n10043, n10044, n10045,
         n10046, n10047, n10048, n10049, n10050, n10051, n10052, n10053,
         n10054, n10055, n10056, n10057, n10058, n10059, n10060, n10061,
         n10062, n10063, n10064, n10065, n10066, n10067, n10068, n10069,
         n10070, n10071, n10072, n10073, n10074, n10075, n10076, n10077,
         n10078, n10079, n10080, n10081, n10082, n10083, n10084, n10085,
         n10086, n10087, n10088, n10089, n10090, n10091, n10092, n10093,
         n10094, n10095, n10096, n10097, n10098, n10099, n10100, n10101,
         n10102, n10103, n10104, n10105, n10106, n10107, n10108, n10109,
         n10110, n10111, n10112, n10113, n10114, n10115, n10116, n10117,
         n10118, n10119, n10120, n10121, n10122, n10123, n10124, n10125,
         n10126, n10127, n10128, n10129, n10130, n10131, n10132, n10133,
         n10134, n10135, n10136, n10137, n10138, n10139, n10140, n10141,
         n10142, n10143, n10144, n10145, n10146, n10147, n10148, n10149,
         n10150, n10151, n10152, n10153, n10154, n10155, n10156, n10157,
         n10158, n10159, n10160, n10161, n10162, n10163, n10164, n10165,
         n10166, n10167, n10168, n10169, n10170, n10171, n10172, n10173,
         n10174, n10175, n10176, n10177, n10178, n10179, n10180, n10181,
         n10182, n10183, n10184, n10185, n10186, n10187, n10188, n10189,
         n10190, n10191, n10192, n10193, n10194, n10195, n10196, n10197,
         n10198, n10199, n10200, n10201, n10202, n10203, n10204, n10205,
         n10206, n10207, n10208, n10209, n10210, n10211, n10212, n10213,
         n10214, n10215, n10216, n10217, n10218, n10219, n10220, n10221,
         n10222, n10223, n10224, n10225, n10226, n10227, n10228, n10229,
         n10230, n10231, n10232, n10233, n10234, n10235, n10236, n10237,
         n10238, n10239, n10240, n10241, n10242, n10243, n10244, n10245,
         n10246, n10247, n10248, n10249, n10250, n10251, n10252, n10253,
         n10254, n10255, n10256, n10257, n10258, n10259, n10260, n10261,
         n10262, n10263, n10264, n10265, n10266, n10267, n10268, n10269,
         n10270, n10271, n10272, n10273, n10274, n10275, n10276, n10277,
         n10278, n10279, n10280, n10281, n10282, n10283, n10284, n10285,
         n10286, n10287, n10288, n10289, n10290, n10291, n10292, n10293,
         n10294, n10295, n10296, n10297, n10298, n10299, n10300, n10301,
         n10302, n10303, n10304, n10305, n10306, n10307, n10308, n10309,
         n10310, n10311, n10312, n10313, n10314, n10315, n10316, n10317,
         n10318, n10319, n10320, n10321, n10322, n10323, n10324, n10325,
         n10326, n10327, n10328, n10329, n10330, n10331, n10332, n10333,
         n10334, n10335, n10336, n10337, n10338, n10339, n10340, n10341,
         n10342, n10343, n10344, n10345, n10346, n10347, n10348, n10349,
         n10350, n10351, n10352, n10353, n10354, n10355, n10356, n10357,
         n10358, n10359, n10360, n10361, n10362, n10363, n10364, n10365,
         n10366, n10367, n10368, n10369, n10370, n10371, n10372, n10373,
         n10374, n10375, n10376, n10377, n10378, n10379, n10380, n10381,
         n10382, n10383, n10384, n10385, n10386, n10387, n10388, n10389,
         n10390, n10391, n10392, n10393, n10394, n10395, n10396, n10397,
         n10398, n10399, n10400, n10401, n10402, n10403, n10404, n10405,
         n10406, n10407, n10408, n10409, n10410, n10411, n10412, n10413,
         n10414, n10415, n10416, n10417, n10418, n10419, n10420, n10421,
         n10422, n10423, n10424, n10425, n10426, n10427, n10428, n10429,
         n10430, n10431, n10432, n10433, n10434, n10435, n10436, n10437,
         n10438, n10439, n10440, n10441, n10442, n10443, n10444, n10445,
         n10446, n10447, n10448, n10449, n10450, n10451, n10452, n10453,
         n10454, n10455, n10456, n10457, n10458, n10459, n10460, n10461,
         n10462, n10463, n10464, n10465, n10466, n10467, n10468, n10469,
         n10470, n10471, n10472, n10473, n10474, n10475, n10476, n10477,
         n10478, n10479, n10480, n10481, n10482, n10483, n10484, n10485,
         n10486, n10487, n10488, n10489, n10490, n10491, n10492, n10493,
         n10494, n10495, n10496, n10497, n10498, n10499, n10500, n10501,
         n10502, n10503, n10504, n10505, n10506, n10507, n10508, n10509,
         n10510, n10511, n10512, n10513, n10514, n10515, n10516, n10517,
         n10518, n10519, n10520, n10521, n10522, n10523, n10524, n10525,
         n10526, n10527, n10528, n10529, n10530, n10531, n10532, n10533,
         n10534, n10535, n10536, n10537, n10538, n10539, n10540, n10541,
         n10542, n10543, n10544, n10545, n10546, n10547, n10548, n10549,
         n10550, n10551, n10552, n10553, n10554, n10555, n10556, n10557,
         n10558, n10559, n10560, n10561, n10562, n10563, n10564, n10565,
         n10566, n10567, n10568, n10569, n10570, n10571, n10572, n10573,
         n10574, n10575, n10576, n10577, n10578, n10579, n10580, n10581,
         n10582, n10583, n10584, n10585, n10586, n10587, n10588, n10589,
         n10590, n10591, n10592, n10593, n10594, n10595, n10596, n10597,
         n10598, n10599, n10600, n10601, n10602, n10603, n10604, n10605,
         n10606, n10607, n10608, n10609, n10610, n10611, n10612, n10613,
         n10614, n10615, n10616, n10617, n10618, n10619, n10620, n10621,
         n10622, n10623, n10624, n10625, n10626, n10627, n10628, n10629,
         n10630, n10631, n10632, n10633, n10634, n10635, n10636, n10637,
         n10638, n10639, n10640, n10641, n10642, n10643, n10644, n10645,
         n10646, n10647, n10648, n10649, n10650, n10651, n10652, n10653,
         n10654, n10655, n10656, n10657, n10658, n10659, n10660, n10661,
         n10662, n10663, n10664, n10665, n10666, n10667, n10668, n10669,
         n10670, n10671, n10672, n10673, n10674, n10675, n10676, n10677,
         n10678, n10679, n10680, n10681, n10682, n10683, n10684, n10685,
         n10686, n10687, n10688, n10689, n10690, n10691, n10692, n10693,
         n10694, n10695, n10696, n10697, n10698, n10699, n10700, n10701,
         n10702, n10703, n10704, n10705, n10706, n10707, n10708, n10709,
         n10710, n10711, n10712, n10713, n10714, n10715, n10716, n10717,
         n10718, n10719, n10720, n10721, n10722, n10723, n10724, n10725,
         n10726, n10727, n10728, n10729, n10730, n10731, n10732, n10733,
         n10734, n10735, n10736, n10737, n10738, n10739, n10740, n10741,
         n10742, n10743, n10744, n10745, n10746, n10747, n10748, n10749,
         n10750, n10751, n10752, n10753, n10754, n10755, n10756, n10757,
         n10758, n10759, n10760, n10761, n10762, n10763, n10764, n10765,
         n10766, n10767, n10768, n10769, n10770, n10771, n10772, n10773,
         n10774, n10775, n10776, n10777, n10778, n10779, n10780, n10781,
         n10782, n10783, n10784, n10785, n10786, n10787, n10788, n10789,
         n10790, n10791, n10792, n10793, n10794, n10795, n10796, n10797,
         n10798, n10799, n10800, n10801, n10802, n10803, n10804, n10805,
         n10806, n10807, n10808, n10809, n10810, n10811, n10812, n10813,
         n10814, n10815, n10816, n10817, n10818, n10819, n10820, n10821,
         n10822, n10823, n10824, n10825, n10826, n10827, n10828, n10829,
         n10830, n10831, n10832, n10833, n10834, n10835, n10836, n10837,
         n10838, n10839, n10840, n10841, n10842, n10843, n10844, n10845,
         n10846, n10847, n10848, n10849, n10850, n10851, n10852, n10853,
         n10854, n10855, n10856, n10857, n10858, n10859, n10860, n10861,
         n10862, n10863, n10864, n10865, n10866, n10867, n10868, n10869,
         n10870, n10871, n10872, n10873, n10874, n10875, n10876, n10877,
         n10878, n10879, n10880, n10881, n10882, n10883, n10884, n10885,
         n10886, n10887, n10888, n10889, n10890, n10891, n10892, n10893,
         n10894, n10895, n10896, n10897, n10898, n10899, n10900, n10901,
         n10902, n10903, n10904, n10905, n10906, n10907, n10908, n10909,
         n10910, n10911, n10912, n10913, n10914, n10915, n10916, n10917,
         n10918, n10919, n10920, n10921, n10922, n10923, n10924, n10925,
         n10926, n10927, n10928, n10929, n10930, n10931, n10932, n10933,
         n10934, n10935, n10936, n10937, n10938, n10939, n10940, n10941,
         n10942, n10943, n10944, n10945, n10946, n10947, n10948, n10949,
         n10950, n10951, n10952, n10953, n10954, n10955, n10956, n10957,
         n10958, n10959, n10960, n10961, n10962, n10963, n10964, n10965,
         n10966, n10967, n10968, n10969, n10970, n10971, n10972, n10973,
         n10974, n10975, n10976, n10977, n10978, n10979, n10980, n10981,
         n10982, n10983, n10984, n10985, n10986, n10987, n10988, n10989,
         n10990, n10991, n10992, n10993, n10994, n10995, n10996, n10997,
         n10998, n10999, n11000, n11001, n11002, n11003, n11004, n11005,
         n11006, n11007, n11008, n11009, n11010, n11011, n11012, n11013,
         n11014, n11015, n11016, n11017, n11018, n11019, n11020, n11021,
         n11022, n11023, n11024, n11025, n11026, n11027, n11028, n11029,
         n11030, n11031, n11032, n11033, n11034, n11035, n11036, n11037,
         n11038, n11039, n11040, n11041, n11042, n11043, n11044, n11045,
         n11046, n11047, n11048, n11049, n11050, n11051, n11052, n11053,
         n11054, n11055, n11056, n11057, n11058, n11059, n11060, n11061,
         n11062, n11063, n11064, n11065, n11066, n11067, n11068, n11069,
         n11070, n11071, n11072, n11073, n11074, n11075, n11076, n11077,
         n11078, n11079, n11080, n11081, n11082, n11083, n11084, n11085,
         n11086, n11087, n11088, n11089, n11090, n11091, n11092, n11093,
         n11094, n11095, n11096, n11097, n11098, n11099, n11100, n11101,
         n11102, n11103, n11104, n11105, n11106, n11107, n11108, n11109,
         n11110, n11111, n11112, n11113, n11114, n11115, n11116, n11117,
         n11118, n11119, n11120, n11121, n11122, n11123, n11124, n11125,
         n11126, n11127, n11128, n11129, n11130, n11131, n11132, n11133,
         n11134, n11135, n11136, n11137, n11138, n11139, n11140, n11141,
         n11142, n11143, n11144, n11145, n11146, n11147, n11148, n11149,
         n11150, n11151, n11152, n11153, n11154, n11155, n11156, n11157,
         n11158, n11159, n11160, n11161, n11162, n11163, n11164, n11165,
         n11166, n11167, n11168, n11169, n11170, n11171, n11172, n11173,
         n11174, n11175, n11176, n11177, n11178, n11179, n11180, n11181,
         n11182, n11183, n11184, n11185, n11186, n11187, n11188, n11189,
         n11190, n11191, n11192, n11193, n11194, n11195, n11196, n11197,
         n11198, n11199, n11200, n11201, n11202, n11203, n11204, n11205,
         n11206, n11207, n11208, n11209, n11210, n11211, n11212, n11213,
         n11214, n11215, n11216, n11217, n11218, n11219, n11220, n11221,
         n11222, n11223, n11224, n11225, n11226, n11227, n11228, n11229,
         n11230, n11231, n11232, n11233, n11234, n11235, n11236, n11237,
         n11238, n11239, n11240, n11241, n11242, n11243, n11244, n11245,
         n11246, n11247, n11248, n11249, n11250, n11251, n11252, n11253,
         n11254, n11255, n11256, n11257, n11258, n11259, n11260, n11261,
         n11262, n11263, n11264, n11265, n11266, n11267, n11268, n11269,
         n11270, n11271, n11272, n11273, n11274, n11275, n11276, n11277,
         n11278, n11279, n11280, n11281, n11282, n11283, n11284, n11285,
         n11286, n11287, n11288, n11289, n11290, n11291, n11292, n11293,
         n11294, n11295, n11296, n11297, n11298, n11299, n11300, n11301,
         n11302, n11303, n11304, n11305, n11306, n11307, n11308, n11309,
         n11310, n11311, n11312, n11313, n11314, n11315, n11316, n11317,
         n11318, n11319, n11320, n11321, n11322, n11323, n11324, n11325,
         n11326, n11327, n11328, n11329, n11330, n11331, n11332, n11333,
         n11334, n11335, n11336, n11337, n11338, n11339, n11340, n11341,
         n11342, n11343, n11344, n11345, n11346, n11347, n11348, n11349,
         n11350, n11351, n11352, n11353, n11354, n11355, n11356, n11357,
         n11358, n11359, n11360, n11361, n11362, n11363, n11364, n11365,
         n11366, n11367, n11368, n11369, n11370, n11371, n11372, n11373,
         n11374, n11375, n11376, n11377, n11378, n11379, n11380, n11381,
         n11382, n11383, n11384, n11385, n11386, n11387, n11388, n11389,
         n11390, n11391, n11392, n11393, n11394, n11395, n11396, n11397,
         n11398, n11399, n11400, n11401, n11402, n11403, n11404, n11405,
         n11406, n11407, n11408, n11409, n11410, n11411, n11412, n11413,
         n11414, n11415, n11416, n11417, n11418, n11419, n11420, n11421,
         n11422, n11423, n11424, n11425, n11426, n11427, n11428, n11429,
         n11430, n11431, n11432, n11433, n11434, n11435, n11436, n11437,
         n11438, n11439, n11440, n11441, n11442, n11443, n11444, n11445,
         n11446, n11447, n11448, n11449, n11450, n11451, n11452, n11453,
         n11454, n11455, n11456, n11457, n11458, n11459, n11460, n11461,
         n11462, n11463, n11464, n11465, n11466, n11467, n11468, n11469,
         n11470, n11471, n11472, n11473, n11474, n11475, n11476, n11477,
         n11478, n11479, n11480, n11481, n11482, n11483, n11484, n11485,
         n11486, n11487, n11488, n11489, n11490, n11491, n11492, n11493,
         n11494, n11495, n11496, n11497, n11498, n11499, n11500, n11501,
         n11502, n11503, n11504, n11505, n11506, n11507, n11508, n11509,
         n11510, n11511, n11512, n11513, n11514, n11515, n11516, n11517,
         n11518, n11519, n11520, n11521, n11522, n11523, n11524, n11525,
         n11526, n11527, n11528, n11529, n11530, n11531, n11532, n11533,
         n11534, n11535, n11536, n11537, n11538, n11539, n11540, n11541,
         n11542, n11543, n11544, n11545, n11546, n11547, n11548, n11549,
         n11550, n11551, n11552, n11553, n11554, n11555, n11556, n11557,
         n11558, n11559, n11560, n11561, n11562, n11563, n11564, n11565,
         n11566, n11567, n11568, n11569, n11570, n11571, n11572, n11573,
         n11574, n11575, n11576, n11577, n11578, n11579, n11580, n11581,
         n11582, n11583, n11584, n11585, n11586, n11587, n11588, n11589,
         n11590, n11591, n11592, n11593, n11594, n11595, n11596, n11597,
         n11598, n11599, n11600, n11601, n11602, n11603, n11604, n11605,
         n11606, n11607, n11608, n11609, n11610, n11611, n11612, n11613,
         n11614, n11615, n11616, n11617, n11618, n11619, n11620, n11621,
         n11622, n11623, n11624, n11625, n11626, n11627, n11628, n11629,
         n11630, n11631, n11632, n11633, n11634, n11635, n11636, n11637,
         n11638, n11639, n11640, n11641, n11642, n11643, n11644, n11645,
         n11646, n11647, n11648, n11649, n11650, n11651, n11652, n11653,
         n11654, n11655, n11656, n11657, n11658, n11659, n11660, n11661,
         n11662, n11663, n11664, n11665, n11666, n11667, n11668, n11669,
         n11670, n11671, n11672, n11673, n11674, n11675, n11676, n11677,
         n11678, n11679, n11680, n11681, n11682, n11683, n11684, n11685,
         n11686, n11687, n11688, n11689, n11690, n11691, n11692, n11693,
         n11694, n11695, n11696, n11697, n11698, n11699, n11700, n11701,
         n11702, n11703, n11704, n11705, n11706, n11707, n11708, n11709,
         n11710, n11711, n11712, n11713, n11714, n11715, n11716, n11717,
         n11718, n11719, n11720, n11721, n11722, n11723, n11724, n11725,
         n11726, n11727, n11728, n11729, n11730, n11731, n11732, n11733,
         n11734, n11735, n11736, n11737, n11738, n11739, n11740, n11741,
         n11742, n11743, n11744, n11745, n11746, n11747, n11748, n11749,
         n11750, n11751, n11752, n11753, n11754, n11755, n11756, n11757,
         n11758, n11759, n11760, n11761, n11762, n11763, n11764, n11765,
         n11766, n11767, n11768, n11769, n11770, n11771, n11772, n11773,
         n11774, n11775, n11776, n11777, n11778, n11779, n11780, n11781,
         n11782, n11783, n11784, n11785, n11786, n11787, n11788, n11789,
         n11790, n11791, n11792, n11793, n11794, n11795, n11796, n11797,
         n11798, n11799, n11800, n11801, n11802, n11803, n11804, n11805,
         n11806, n11807, n11808, n11809, n11810, n11811, n11812, n11813,
         n11814, n11815, n11816, n11817, n11818, n11819, n11820, n11821,
         n11822, n11823, n11824, n11825, n11826, n11827, n11828, n11829,
         n11830, n11831, n11832, n11833, n11834, n11835, n11836, n11837,
         n11838, n11839, n11840, n11841, n11842, n11843, n11844, n11845,
         n11846, n11847, n11848, n11849, n11850, n11851, n11852, n11853,
         n11854, n11855, n11856, n11857, n11858, n11859, n11860, n11861,
         n11862, n11863, n11864, n11865, n11866, n11867, n11868, n11869,
         n11870, n11871, n11872, n11873, n11874, n11875, n11876, n11877,
         n11878, n11879, n11880, n11881, n11882, n11883, n11884, n11885,
         n11886, n11887, n11888, n11889, n11890, n11891, n11892, n11893,
         n11894, n11895, n11896, n11897, n11898, n11899, n11900, n11901,
         n11902, n11903, n11904, n11905, n11906, n11907, n11908, n11909,
         n11910, n11911, n11912, n11913, n11914, n11915, n11916, n11917,
         n11918, n11919, n11920, n11921, n11922, n11923, n11924, n11925,
         n11926, n11927, n11928, n11929, n11930, n11931, n11932, n11933,
         n11934, n11935, n11936, n11937, n11938, n11939, n11940, n11941,
         n11942, n11943, n11944, n11945, n11946, n11947, n11948, n11949,
         n11950, n11951, n11952, n11953, n11954, n11955, n11956, n11957,
         n11958, n11959, n11960, n11961, n11962, n11963, n11964, n11965,
         n11966, n11967, n11968, n11969, n11970, n11971, n11972, n11973,
         n11974, n11975, n11976, n11977, n11978, n11979, n11980, n11981,
         n11982, n11983, n11984, n11985, n11986, n11987, n11988, n11989,
         n11990, n11991, n11992, n11993, n11994, n11995, n11996, n11997,
         n11998, n11999, n12000, n12001, n12002, n12003, n12004, n12005,
         n12006, n12007, n12008, n12009, n12010, n12011, n12012, n12013,
         n12014, n12015, n12016, n12017, n12018, n12019, n12020, n12021,
         n12022, n12023, n12024, n12025, n12026, n12027, n12028, n12029,
         n12030, n12031, n12032, n12033, n12034, n12035, n12036, n12037,
         n12038, n12039, n12040, n12041, n12042, n12043, n12044, n12045,
         n12046, n12047, n12048, n12049, n12050, n12051, n12052, n12053,
         n12054, n12055, n12056, n12057, n12058, n12059, n12060, n12061,
         n12062, n12063, n12064, n12065, n12066, n12067, n12068, n12069,
         n12070, n12071, n12072, n12073, n12074, n12075, n12076, n12077,
         n12078, n12079, n12080, n12081, n12082, n12083, n12084, n12085,
         n12086, n12087, n12088, n12089, n12090, n12091, n12092, n12093,
         n12094, n12095, n12096, n12097, n12098, n12099, n12100, n12101,
         n12102, n12103, n12104, n12105, n12106, n12107, n12108, n12109,
         n12110, n12111, n12112, n12113, n12114, n12115, n12116, n12117,
         n12118, n12119, n12120, n12121, n12122, n12123, n12124, n12125,
         n12126, n12127, n12128, n12129, n12130, n12131, n12132, n12133,
         n12134, n12135, n12136, n12137, n12138, n12139, n12140, n12141,
         n12142, n12143, n12144, n12145, n12146, n12147, n12148, n12149,
         n12150, n12151, n12152, n12153, n12154, n12155, n12156, n12157,
         n12158, n12159, n12160, n12161, n12162, n12163, n12164, n12165,
         n12166, n12167, n12168, n12169, n12170, n12171, n12172, n12173,
         n12174, n12175, n12176, n12177, n12178, n12179, n12180, n12181,
         n12182, n12183, n12184, n12185, n12186, n12187, n12188, n12189,
         n12190, n12191, n12192, n12193, n12194, n12195, n12196, n12197,
         n12198, n12199, n12200, n12201, n12202, n12203, n12204, n12205,
         n12206, n12207, n12208, n12209, n12210, n12211, n12212, n12213,
         n12214, n12215, n12216, n12217, n12218, n12219, n12220, n12221,
         n12222, n12223, n12224, n12225, n12226, n12227, n12228, n12229,
         n12230, n12231, n12232, n12233, n12234, n12235, n12236, n12237,
         n12238, n12239, n12240, n12241, n12242, n12243, n12244, n12245,
         n12246, n12247, n12248, n12249, n12250, n12251, n12252, n12253,
         n12254, n12255, n12256, n12257, n12258, n12259, n12260, n12261,
         n12262, n12263, n12264, n12265, n12266, n12267, n12268, n12269,
         n12270, n12271, n12272, n12273, n12274, n12275, n12276, n12277,
         n12278, n12279, n12280, n12281, n12282, n12283, n12284, n12285,
         n12286, n12287, n12288, n12289, n12290, n12291, n12292, n12293,
         n12294, n12295, n12296, n12297, n12298, n12299, n12300, n12301,
         n12302, n12303, n12304, n12305, n12306, n12307, n12308, n12309,
         n12310, n12311, n12312, n12313, n12314, n12315, n12316, n12317,
         n12318, n12319, n12320, n12321, n12322, n12323, n12324, n12325,
         n12326, n12327, n12328, n12329, n12330, n12331, n12332, n12333,
         n12334, n12335, n12336, n12337, n12338, n12339, n12340, n12341,
         n12342, n12343, n12344, n12345, n12346, n12347, n12348, n12349,
         n12350, n12351, n12352, n12353, n12354, n12355, n12356, n12357,
         n12358, n12359, n12360, n12361, n12362, n12363, n12364, n12365,
         n12366, n12367, n12368, n12369, n12370, n12371, n12372, n12373,
         n12374, n12375, n12376, n12377, n12378, n12379, n12380, n12381,
         n12382, n12383, n12384, n12385, n12386, n12387, n12388, n12389,
         n12390, n12391, n12392, n12393, n12394, n12395, n12396, n12397,
         n12398, n12399, n12400, n12401, n12402, n12403, n12404, n12405,
         n12406, n12407, n12408, n12409, n12410, n12411, n12412, n12413,
         n12414, n12415, n12416, n12417, n12418, n12419, n12420, n12421,
         n12422, n12423, n12424, n12425, n12426, n12427, n12428, n12429,
         n12430, n12431, n12432, n12433, n12434, n12435, n12436, n12437,
         n12438, n12439, n12440, n12441, n12442, n12443, n12444, n12445,
         n12446, n12447, n12448, n12449, n12450, n12451, n12452, n12453,
         n12454, n12455, n12456, n12457, n12458, n12459, n12460, n12461,
         n12462, n12463, n12464, n12465, n12466, n12467, n12468, n12469,
         n12470, n12471, n12472, n12473, n12474, n12475, n12476, n12477,
         n12478, n12479, n12480, n12481, n12482, n12483, n12484, n12485,
         n12486, n12487, n12488, n12489, n12490, n12491, n12492, n12493,
         n12494, n12495, n12496, n12497, n12498, n12499, n12500, n12501,
         n12502, n12503, n12504, n12505, n12506, n12507, n12508, n12509,
         n12510, n12511, n12512, n12513, n12514, n12515, n12516, n12517,
         n12518, n12519, n12520, n12521, n12522, n12523, n12524, n12525,
         n12526, n12527, n12528, n12529, n12530, n12531, n12532, n12533,
         n12534, n12535, n12536, n12537, n12538, n12539, n12540, n12541,
         n12542, n12543, n12544, n12545, n12546, n12547, n12548, n12549,
         n12550, n12551, n12552, n12553, n12554, n12555, n12556, n12557,
         n12558, n12559, n12560, n12561, n12562, n12563, n12564, n12565,
         n12566, n12567, n12568, n12569, n12570, n12571, n12572, n12573,
         n12574, n12575, n12576, n12577, n12578, n12579, n12580, n12581,
         n12582, n12583, n12584, n12585, n12586, n12587, n12588, n12589,
         n12590, n12591, n12592, n12593, n12594, n12595, n12596, n12597,
         n12598, n12599, n12600, n12601, n12602, n12603, n12604, n12605,
         n12606, n12607, n12608, n12609, n12610, n12611, n12612, n12613,
         n12614, n12615, n12616, n12617, n12618, n12619, n12620, n12621,
         n12622, n12623, n12624, n12625, n12626, n12627, n12628, n12629,
         n12630, n12631, n12632, n12633, n12634, n12635, n12636, n12637,
         n12638, n12639, n12640, n12641, n12642, n12643, n12644, n12645,
         n12646, n12647, n12648, n12649, n12650, n12651, n12652, n12653,
         n12654, n12655, n12656, n12657, n12658, n12659, n12660, n12661,
         n12662, n12663, n12664, n12665, n12666, n12667, n12668, n12669,
         n12670, n12671, n12672, n12673, n12674, n12675, n12676, n12677,
         n12678, n12679, n12680, n12681, n12682, n12683, n12684, n12685,
         n12686, n12687, n12688, n12689, n12690, n12691, n12692, n12693,
         n12694, n12695, n12696, n12697, n12698, n12699, n12700, n12701,
         n12702, n12703, n12704, n12705, n12706, n12707, n12708, n12709,
         n12710, n12711, n12712, n12713, n12714, n12715, n12716, n12717,
         n12718, n12719, n12720, n12721, n12722, n12723, n12724, n12725,
         n12726, n12727, n12728, n12729, n12730, n12731, n12732, n12733,
         n12734, n12735, n12736, n12737, n12738, n12739, n12740, n12741,
         n12742, n12743, n12744, n12745, n12746, n12747, n12748, n12749,
         n12750, n12751, n12752, n12753, n12754, n12755, n12756, n12757,
         n12758, n12759, n12760, n12761, n12762, n12763, n12764, n12765,
         n12766, n12767, n12768, n12769, n12770, n12771, n12772, n12773,
         n12774, n12775, n12776, n12777, n12778, n12779, n12780, n12781,
         n12782, n12783, n12784, n12785, n12786, n12787, n12788, n12789,
         n12790, n12791, n12792, n12793, n12794, n12795, n12796, n12797,
         n12798, n12799, n12800, n12801, n12802, n12803, n12804, n12805,
         n12806, n12807, n12808, n12809, n12810, n12811, n12812, n12813,
         n12814, n12815, n12816, n12817, n12818, n12819, n12820, n12821,
         n12822, n12823, n12824, n12825, n12826, n12827, n12828, n12829,
         n12830, n12831, n12832, n12833, n12834, n12835, n12836, n12837,
         n12838, n12839, n12840, n12841, n12842, n12843, n12844, n12845,
         n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         n13014, n13015, n13016, n13017, n13018, n13019, n13020, n13021,
         n13022, n13023, n13024, n13025, n13026, n13027, n13028, n13029,
         n13030, n13031, n13032, n13033, n13034, n13035, n13036, n13037,
         n13038, n13039, n13040, n13041, n13042, n13043, n13044, n13045,
         n13046, n13047, n13048, n13049, n13050, n13051, n13052, n13053,
         n13054, n13055, n13056, n13057, n13058, n13059, n13060, n13061,
         n13062, n13063, n13064, n13065, n13066, n13067, n13068, n13069,
         n13070, n13071, n13072, n13073, n13074, n13075, n13076, n13077,
         n13078, n13079, n13080, n13081, n13082, n13083, n13084, n13085,
         n13086, n13087, n13088, n13089, n13090, n13091, n13092, n13093,
         n13094, n13095, n13096, n13097, n13098, n13099, n13100, n13101,
         n13102, n13103, n13104, n13105, n13106, n13107, n13108, n13109,
         n13110, n13111, n13112, n13113, n13114, n13115, n13116, n13117,
         n13118, n13119, n13120, n13121, n13122, n13123, n13124, n13125,
         n13126, n13127, n13128, n13129, n13130, n13131, n13132, n13133,
         n13134, n13135, n13136, n13137, n13138, n13139, n13140, n13141,
         n13142, n13143, n13144, n13145, n13146, n13147, n13148, n13149,
         n13150, n13151, n13152, n13153, n13154, n13155, n13156, n13157,
         n13158, n13159, n13160, n13161, n13162, n13163, n13164, n13165,
         n13166, n13167, n13168, n13169, n13170, n13171, n13172, n13173,
         n13174, n13175, n13176, n13177, n13178, n13179, n13180, n13181,
         n13182, n13183, n13184, n13185, n13186, n13187, n13188, n13189,
         n13190, n13191, n13192, n13193, n13194, n13195, n13196, n13197,
         n13198, n13199, n13200, n13201, n13202, n13203, n13204, n13205,
         n13206, n13207, n13208, n13209, n13210, n13211, n13212, n13213,
         n13214, n13215, n13216, n13217, n13218, n13219, n13220, n13221,
         n13222, n13223, n13224, n13225, n13226, n13227, n13228, n13229,
         n13230, n13231, n13232, n13233, n13234, n13235, n13236, n13237,
         n13238, n13239, n13240, n13241, n13242, n13243, n13244, n13245,
         n13246, n13247, n13248, n13249, n13250, n13251, n13252, n13253,
         n13254, n13255, n13256, n13257, n13258, n13259, n13260, n13261,
         n13262, n13263, n13264, n13265, n13266, n13267, n13268, n13269,
         n13270, n13271, n13272, n13273, n13274, n13275, n13276, n13277,
         n13278, n13279, n13280, n13281, n13282, n13283, n13284, n13285,
         n13286, n13287, n13288, n13289, n13290, n13291, n13292, n13293,
         n13294, n13295, n13296, n13297, n13298, n13299, n13300, n13301,
         n13302, n13303, n13304, n13305, n13306, n13307, n13308, n13309,
         n13310, n13311, n13312, n13313, n13314, n13315, n13316, n13317,
         n13318, n13319, n13320, n13321, n13322, n13323, n13324, n13325,
         n13326, n13327, n13328, n13329, n13330, n13331, n13332, n13333,
         n13334, n13335, n13336, n13337, n13338, n13339, n13340, n13341,
         n13342, n13343, n13344, n13345, n13346, n13347, n13348, n13349,
         n13350, n13351, n13352, n13353, n13354, n13355, n13356, n13357,
         n13358, n13359, n13360, n13361, n13362, n13363, n13364, n13365,
         n13366, n13367, n13368, n13369, n13370, n13371, n13372, n13373,
         n13374, n13375, n13376, n13377, n13378, n13379, n13380, n13381,
         n13382, n13383, n13384, n13385, n13386, n13387, n13388, n13389,
         n13390, n13391, n13392, n13393, n13394, n13395, n13396, n13397,
         n13398, n13399, n13400, n13401, n13402, n13403, n13404, n13405,
         n13406, n13407, n13408, n13409, n13410, n13411, n13412, n13413,
         n13414, n13415, n13416, n13417, n13418, n13419, n13420, n13421,
         n13422, n13423, n13424, n13425, n13426, n13427, n13428, n13429,
         n13430, n13431, n13432, n13433, n13434, n13435, n13436, n13437,
         n13438, n13439, n13440, n13441, n13442, n13443, n13444, n13445,
         n13446, n13447, n13448, n13449, n13450, n13451, n13452, n13453,
         n13454, n13455, n13456, n13457, n13458, n13459, n13460, n13461,
         n13462, n13463, n13464, n13465, n13466, n13467, n13468, n13469,
         n13470, n13471, n13472, n13473, n13474, n13475, n13476, n13477,
         n13478, n13479, n13480, n13481, n13482, n13483, n13484, n13485,
         n13486, n13487, n13488, n13489, n13490, n13491, n13492, n13493,
         n13494, n13495, n13496, n13497, n13498, n13499, n13500, n13501,
         n13502, n13503, n13504, n13505, n13506, n13507, n13508, n13509,
         n13510, n13511, n13512, n13513, n13514, n13515, n13516, n13517,
         n13518, n13519, n13520, n13521, n13522, n13523, n13524, n13525,
         n13526, n13527, n13528, n13529, n13530, n13531, n13532, n13533,
         n13534, n13535, n13536, n13537, n13538, n13539, n13540, n13541,
         n13542, n13543, n13544, n13545, n13546, n13547, n13548, n13549,
         n13550, n13551, n13552, n13553, n13554, n13555, n13556, n13557,
         n13558, n13559, n13560, n13561, n13562, n13563, n13564, n13565,
         n13566, n13567, n13568, n13569, n13570, n13571, n13572, n13573,
         n13574, n13575, n13576, n13577, n13578, n13579, n13580, n13581,
         n13582, n13583, n13584, n13585, n13586, n13587, n13588, n13589,
         n13590, n13591, n13592, n13593, n13594, n13595, n13596, n13597,
         n13598, n13599, n13600, n13601, n13602, n13603, n13604, n13605,
         n13606, n13607, n13608, n13609, n13610, n13611, n13612, n13613,
         n13614, n13615, n13616, n13617, n13618, n13619, n13620, n13621,
         n13622, n13623, n13624, n13625, n13626, n13627, n13628, n13629,
         n13630, n13631, n13632, n13633, n13634, n13635, n13636, n13637,
         n13638, n13639, n13640, n13641, n13642, n13643, n13644, n13645,
         n13646, n13647, n13648, n13649, n13650, n13651, n13652, n13653,
         n13654, n13655, n13656, n13657, n13658, n13659, n13660, n13661,
         n13662, n13663, n13664, n13665, n13666, n13667, n13668, n13669,
         n13670, n13671, n13672, n13673, n13674, n13675, n13676, n13677,
         n13678, n13679, n13680, n13681, n13682, n13683, n13684, n13685,
         n13686, n13687, n13688, n13689, n13690, n13691, n13692, n13693,
         n13694, n13695, n13696, n13697, n13698, n13699, n13700, n13701,
         n13702, n13703, n13704, n13705, n13706, n13707, n13708, n13709,
         n13710, n13711, n13712, n13713, n13714, n13715, n13716, n13717,
         n13718, n13719, n13720, n13721, n13722, n13723, n13724, n13725,
         n13726, n13727, n13728, n13729, n13730, n13731, n13732, n13733,
         n13734, n13735, n13736, n13737, n13738, n13739, n13740, n13741,
         n13742, n13743, n13744, n13745, n13746, n13747, n13748, n13749,
         n13750, n13751, n13752, n13753, n13754, n13755, n13756, n13757,
         n13758, n13759, n13760, n13761, n13762, n13763, n13764, n13765,
         n13766, n13767, n13768, n13769, n13770, n13771, n13772, n13773,
         n13774, n13775, n13776, n13777, n13778, n13779, n13780, n13781,
         n13782, n13783, n13784, n13785, n13786, n13787, n13788, n13789,
         n13790, n13791, n13792, n13793, n13794, n13795, n13796, n13797,
         n13798, n13799, n13800, n13801, n13802, n13803, n13804, n13805,
         n13806, n13807, n13808, n13809, n13810, n13811, n13812, n13813,
         n13814, n13815, n13816, n13817, n13818, n13819, n13820, n13821,
         n13822, n13823, n13824, n13825, n13826, n13827, n13828, n13829,
         n13830, n13831, n13832, n13833, n13834, n13835, n13836, n13837,
         n13838, n13839, n13840, n13841, n13842, n13843, n13844, n13845,
         n13846, n13847, n13848, n13849, n13850, n13851, n13852, n13853,
         n13854, n13855, n13856, n13857, n13858, n13859, n13860, n13861,
         n13862, n13863, n13864, n13865, n13866, n13867, n13868, n13869,
         n13870, n13871, n13872, n13873, n13874, n13875, n13876, n13877,
         n13878, n13879, n13880, n13881, n13882, n13883, n13884, n13885,
         n13886, n13887, n13888, n13889, n13890, n13891, n13892, n13893,
         n13894, n13895, n13896, n13897, n13898, n13899, n13900, n13901,
         n13902, n13903, n13904, n13905, n13906, n13907, n13908, n13909,
         n13910, n13911, n13912, n13913, n13914, n13915, n13916, n13917,
         n13918, n13919, n13920, n13921, n13922, n13923, n13924, n13925,
         n13926, n13927, n13928, n13929, n13930, n13931, n13932, n13933,
         n13934, n13935, n13936, n13937, n13938, n13939, n13940, n13941,
         n13942, n13943, n13944, n13945, n13946, n13947, n13948, n13949,
         n13950, n13951, n13952, n13953, n13954, n13955, n13956, n13957,
         n13958, n13959, n13960, n13961, n13962, n13963, n13964, n13965,
         n13966, n13967, n13968, n13969, n13970, n13971, n13972, n13973,
         n13974, n13975, n13976, n13977, n13978, n13979, n13980, n13981,
         n13982, n13983, n13984, n13985, n13986, n13987, n13988, n13989,
         n13990, n13991, n13992, n13993, n13994, n13995, n13996, n13997,
         n13998, n13999, n14000, n14001, n14002, n14003, n14004, n14005,
         n14006, n14007, n14008, n14009, n14010, n14011, n14012, n14013,
         n14014, n14015, n14016, n14017, n14018, n14019, n14020, n14021,
         n14022, n14023, n14024, n14025, n14026, n14027, n14028, n14029,
         n14030, n14031, n14032, n14033, n14034, n14035, n14036, n14037,
         n14038, n14039, n14040, n14041, n14042, n14043, n14044, n14045,
         n14046, n14047, n14048, n14049, n14050, n14051, n14052, n14053,
         n14054, n14055, n14056, n14057, n14058, n14059, n14060, n14061,
         n14062, n14063, n14064, n14065, n14066, n14067, n14068, n14069,
         n14070, n14071, n14072, n14073, n14074, n14075, n14076, n14077,
         n14078, n14079, n14080, n14081, n14082, n14083, n14084, n14085,
         n14086, n14087, n14088, n14089, n14090, n14091, n14092, n14093,
         n14094, n14095, n14096, n14097, n14098, n14099, n14100, n14101,
         n14102, n14103, n14104, n14105, n14106, n14107, n14108, n14109,
         n14110, n14111, n14112, n14113, n14114, n14115, n14116, n14117,
         n14118, n14119, n14120, n14121, n14122, n14123, n14124, n14125,
         n14126, n14127, n14128, n14129, n14130, n14131, n14132, n14133,
         n14134, n14135, n14136, n14137, n14138, n14139, n14140, n14141,
         n14142, n14143, n14144, n14145, n14146, n14147, n14148, n14149,
         n14150, n14151, n14152, n14153, n14154, n14155, n14156, n14157,
         n14158, n14159, n14160, n14161, n14162, n14163, n14164, n14165,
         n14166, n14167, n14168, n14169, n14170, n14171, n14172, n14173,
         n14174, n14175, n14176, n14177, n14178, n14179, n14180, n14181,
         n14182, n14183, n14184, n14185, n14186, n14187, n14188, n14189,
         n14190, n14191, n14192, n14193, n14194, n14195, n14196, n14197,
         n14198, n14199, n14200, n14201, n14202, n14203, n14204, n14205,
         n14206, n14207, n14208, n14209, n14210, n14211, n14212, n14213,
         n14214, n14215, n14216, n14217, n14218, n14219, n14220, n14221,
         n14222, n14223, n14224, n14225, n14226, n14227, n14228, n14229,
         n14230, n14231, n14232, n14233, n14234, n14235, n14236, n14237,
         n14238, n14239, n14240, n14241, n14242, n14243, n14244, n14245,
         n14246, n14247, n14248, n14249, n14250, n14251, n14252, n14253,
         n14254, n14255, n14256, n14257, n14258, n14259, n14260, n14261,
         n14262, n14263, n14264, n14265, n14266, n14267, n14268, n14269,
         n14270, n14271, n14272, n14273, n14274, n14275, n14276, n14277,
         n14278, n14279, n14280, n14281, n14282, n14283, n14284, n14285,
         n14286, n14287, n14288, n14289, n14290, n14291, n14292, n14293,
         n14294, n14295, n14296, n14297, n14298, n14299, n14300, n14301,
         n14302, n14303, n14304, n14305, n14306, n14307, n14308, n14309,
         n14310, n14311, n14312, n14313, n14314, n14315, n14316, n14317,
         n14318, n14319, n14320, n14321, n14322, n14323, n14324, n14325,
         n14326, n14327, n14328, n14329, n14330, n14331, n14332, n14333,
         n14334, n14335, n14336, n14337, n14338, n14339, n14340, n14341,
         n14342, n14343, n14344, n14345, n14346, n14347, n14348, n14349,
         n14350, n14351, n14352, n14353, n14354, n14355, n14356, n14357,
         n14358, n14359, n14360, n14361, n14362, n14363, n14364, n14365,
         n14366, n14367, n14368, n14369, n14370, n14371, n14372, n14373,
         n14374, n14375, n14376, n14377, n14378, n14379, n14380, n14381,
         n14382, n14383, n14384, n14385, n14386, n14387, n14388, n14389,
         n14390, n14391, n14392, n14393, n14394, n14395, n14396, n14397,
         n14398, n14399, n14400, n14401, n14402, n14403, n14404, n14405,
         n14406, n14407, n14408, n14409, n14410, n14411, n14412, n14413,
         n14414, n14415, n14416, n14417, n14418, n14419, n14420, n14421,
         n14422, n14423, n14424, n14425, n14426, n14427, n14428, n14429,
         n14430, n14431, n14432, n14433, n14434, n14435, n14436, n14437,
         n14438, n14439, n14440, n14441, n14442, n14443, n14444, n14445,
         n14446, n14447, n14448, n14449, n14450, n14451, n14452, n14453,
         n14454, n14455, n14456, n14457, n14458, n14459, n14460, n14461,
         n14462, n14463, n14464, n14465, n14466, n14467, n14468, n14469,
         n14470, n14471, n14472, n14473, n14474, n14475, n14476, n14477,
         n14478, n14479, n14480, n14481, n14482, n14483, n14484, n14485,
         n14486, n14487, n14488, n14489, n14490, n14491, n14492, n14493,
         n14494, n14495, n14496, n14497, n14498, n14499, n14500, n14501,
         n14502, n14503, n14504, n14505, n14506, n14507, n14508, n14509,
         n14510, n14511, n14512, n14513, n14514, n14515, n14516, n14517,
         n14518, n14519, n14520, n14521, n14522, n14523, n14524, n14525,
         n14526, n14527, n14528, n14529, n14530, n14531, n14532, n14533,
         n14534, n14535, n14536, n14537, n14538, n14539, n14540, n14541,
         n14542, n14543, n14544, n14545, n14546, n14547, n14548, n14549,
         n14550, n14551, n14552, n14553, n14554, n14555, n14556, n14557,
         n14558, n14559, n14560, n14561, n14562, n14563, n14564, n14565,
         n14566, n14567, n14568, n14569, n14570, n14571, n14572, n14573,
         n14574, n14575, n14576, n14577, n14578, n14579, n14580, n14581,
         n14582, n14583, n14584, n14585, n14586, n14587, n14588, n14589,
         n14590, n14591, n14592, n14593, n14594, n14595, n14596, n14597,
         n14598, n14599, n14600, n14601, n14602, n14603, n14604, n14605,
         n14606, n14607, n14608, n14609, n14610, n14611, n14612, n14613,
         n14614, n14615, n14616, n14617, n14618, n14619, n14620, n14621,
         n14622, n14623, n14624, n14625, n14626, n14627, n14628, n14629,
         n14630, n14631, n14632, n14633, n14634, n14635, n14636, n14637,
         n14638, n14639, n14640, n14641, n14642, n14643, n14644, n14645,
         n14646, n14647, n14648, n14649, n14650, n14651, n14652, n14653,
         n14654, n14655, n14656, n14657, n14658, n14659, n14660, n14661,
         n14662, n14663, n14664, n14665, n14666, n14667, n14668, n14669,
         n14670, n14671, n14672, n14673, n14674, n14675, n14676, n14677,
         n14678, n14679, n14680, n14681, n14682, n14683, n14684, n14685,
         n14686, n14687, n14688, n14689, n14690, n14691, n14692, n14693,
         n14694, n14695, n14696, n14697, n14698, n14699, n14700, n14701,
         n14702, n14703, n14704, n14705, n14706, n14707, n14708, n14709,
         n14710, n14711, n14712, n14713, n14714, n14715, n14716, n14717,
         n14718, n14719, n14720, n14721, n14722, n14723, n14724, n14725,
         n14726, n14727, n14728, n14729, n14730, n14731, n14732, n14733,
         n14734, n14735, n14736, n14737, n14738, n14739, n14740, n14741,
         n14742, n14743, n14744, n14745, n14746, n14747, n14748, n14749,
         n14750, n14751, n14752, n14753, n14754, n14755, n14756, n14757,
         n14758, n14759, n14760, n14761, n14762, n14763, n14764, n14765,
         n14766, n14767, n14768, n14769, n14770, n14771, n14772, n14773,
         n14774, n14775, n14776, n14777, n14778, n14779, n14780, n14781,
         n14782, n14783, n14784, n14785, n14786, n14787, n14788, n14789,
         n14790, n14791, n14792, n14793, n14794, n14795, n14796, n14797,
         n14798, n14799, n14800, n14801, n14802, n14803, n14804, n14805,
         n14806, n14807, n14808, n14809, n14810, n14811, n14812, n14813,
         n14814, n14815, n14816, n14817, n14818, n14819, n14820, n14821,
         n14822, n14823, n14824, n14825, n14826, n14827, n14828, n14829,
         n14830, n14831, n14832, n14833, n14834, n14835, n14836, n14837,
         n14838, n14839, n14840, n14841, n14842, n14843, n14844, n14845,
         n14846, n14847, n14848, n14849, n14850, n14851, n14852, n14853,
         n14854, n14855, n14856, n14857, n14858, n14859, n14860, n14861,
         n14862, n14863, n14864, n14865, n14866, n14867, n14868, n14869,
         n14870, n14871, n14872, n14873, n14874, n14875, n14876, n14877,
         n14878, n14879, n14880, n14881, n14882, n14883, n14884, n14885,
         n14886, n14887, n14888, n14889, n14890, n14891, n14892, n14893,
         n14894, n14895, n14896, n14897, n14898, n14899, n14900, n14901,
         n14902, n14903, n14904, n14905, n14906, n14907, n14908, n14909,
         n14910, n14911, n14912, n14913, n14914, n14915, n14916, n14917,
         n14918, n14919, n14920, n14921, n14922, n14923, n14924, n14925,
         n14926, n14927, n14928, n14929, n14930, n14931, n14932, n14933,
         n14934, n14935, n14936, n14937, n14938, n14939, n14940, n14941,
         n14942, n14943, n14944, n14945, n14946, n14947, n14948, n14949,
         n14950, n14951, n14952, n14953, n14954, n14955, n14956, n14957,
         n14958, n14959, n14960, n14961, n14962, n14963, n14964, n14965,
         n14966, n14967, n14968, n14969, n14970, n14971, n14972, n14973,
         n14974, n14975, n14976, n14977, n14978, n14979, n14980, n14981,
         n14982, n14983, n14984, n14985, n14986, n14987, n14988, n14989,
         n14990, n14991, n14992, n14993, n14994, n14995, n14996, n14997,
         n14998, n14999, n15000, n15001, n15002, n15003, n15004, n15005,
         n15006, n15007, n15008, n15009, n15010, n15011, n15012, n15013,
         n15014, n15015, n15016, n15017, n15018, n15019, n15020, n15021,
         n15022, n15023, n15024, n15025, n15026, n15027, n15028, n15029,
         n15030, n15031, n15032, n15033, n15034, n15035, n15036, n15037,
         n15038, n15039, n15040, n15041, n15042, n15043, n15044, n15045,
         n15046, n15047, n15048, n15049, n15050, n15051, n15052, n15053,
         n15054, n15055, n15056, n15057, n15058, n15059, n15060, n15061,
         n15062, n15063, n15064, n15065, n15066, n15067, n15068, n15069,
         n15070, n15071, n15072, n15073, n15074, n15075, n15076, n15077,
         n15078, n15079, n15080, n15081, n15082, n15083, n15084, n15085,
         n15086, n15087, n15088, n15089, n15090, n15091, n15092, n15093,
         n15094, n15095, n15096, n15097, n15098, n15099, n15100, n15101,
         n15102, n15103, n15104, n15105, n15106, n15107, n15108, n15109,
         n15110, n15111, n15112, n15113, n15114, n15115, n15116, n15117,
         n15118, n15119, n15120, n15121, n15122, n15123, n15124, n15125,
         n15126, n15127, n15128, n15129, n15130, n15131, n15132, n15133,
         n15134, n15135, n15136, n15137, n15138, n15139, n15140, n15141,
         n15142, n15143, n15144, n15145, n15146, n15147, n15148, n15149,
         n15150, n15151, n15152, n15153, n15154, n15155, n15156, n15157,
         n15158, n15159, n15160, n15161, n15162, n15163, n15164, n15165,
         n15166, n15167, n15168, n15169, n15170, n15171, n15172, n15173,
         n15174, n15175, n15176, n15177, n15178, n15179, n15180, n15181,
         n15182, n15183, n15184, n15185, n15186, n15187, n15188, n15189,
         n15190, n15191, n15192, n15193, n15194, n15195, n15196, n15197,
         n15198, n15199, n15200, n15201, n15202, n15203, n15204, n15205,
         n15206, n15207, n15208, n15209, n15210, n15211, n15212, n15213,
         n15214, n15215, n15216, n15217, n15218, n15219, n15220, n15221,
         n15222, n15223, n15224, n15225, n15226, n15227, n15228, n15229,
         n15230, n15231, n15232, n15233, n15234, n15235, n15236, n15237,
         n15238, n15239, n15240, n15241, n15242, n15243, n15244, n15245,
         n15246, n15247, n15248, n15249, n15250, n15251, n15252, n15253,
         n15254, n15255, n15256, n15257, n15258, n15259, n15260, n15261,
         n15262, n15263, n15264, n15265, n15266, n15267, n15268, n15269,
         n15270, n15271, n15272, n15273, n15274, n15275, n15276, n15277,
         n15278, n15279, n15280, n15281, n15282, n15283, n15284, n15285,
         n15286, n15287, n15288, n15289, n15290, n15291, n15292, n15293,
         n15294, n15295, n15296, n15297, n15298, n15299, n15300, n15301,
         n15302, n15303, n15304, n15305, n15306, n15307, n15308, n15309,
         n15310, n15311, n15312, n15313, n15314, n15315, n15316, n15317,
         n15318, n15319, n15320, n15321, n15322, n15323, n15324, n15325,
         n15326, n15327, n15328, n15329, n15330, n15331, n15332, n15333,
         n15334, n15335, n15336, n15337, n15338, n15339, n15340, n15341,
         n15342, n15343, n15344, n15345, n15346, n15347, n15348, n15349,
         n15350, n15351, n15352, n15353, n15354, n15355, n15356, n15357,
         n15358, n15359, n15360, n15361, n15362, n15363, n15364, n15365,
         n15366, n15367, n15368, n15369, n15370, n15371, n15372, n15373,
         n15374, n15375, n15376, n15377, n15378, n15379, n15380, n15381,
         n15382, n15383, n15384, n15385, n15386, n15387, n15388, n15389,
         n15390, n15391, n15392, n15393, n15394, n15395, n15396, n15397,
         n15398, n15399, n15400, n15401, n15402, n15403, n15404, n15405,
         n15406, n15407, n15408, n15409, n15410, n15411, n15412, n15413,
         n15414, n15415, n15416, n15417, n15418, n15419, n15420, n15421,
         n15422, n15423, n15424, n15425, n15426, n15427, n15428, n15429,
         n15430, n15431, n15432, n15433, n15434, n15435, n15436, n15437,
         n15438, n15439, n15440, n15441, n15442, n15443, n15444, n15445,
         n15446, n15447, n15448, n15449, n15450, n15451, n15452, n15453,
         n15454, n15455, n15456, n15457, n15458, n15459, n15460, n15461,
         n15462, n15463, n15464, n15465, n15466, n15467, n15468, n15469,
         n15470, n15471, n15472, n15473, n15474, n15475, n15476, n15477,
         n15478, n15479, n15480, n15481, n15482, n15483, n15484, n15485,
         n15486, n15487, n15488, n15489, n15490, n15491, n15492, n15493,
         n15494, n15495, n15496, n15497, n15498, n15499, n15500, n15501,
         n15502, n15503, n15504, n15505, n15506, n15507, n15508, n15509,
         n15510, n15511, n15512, n15513, n15514, n15515, n15516, n15517,
         n15518, n15519, n15520, n15521, n15522, n15523, n15524, n15525,
         n15526, n15527, n15528, n15529, n15530, n15531, n15532, n15533,
         n15534, n15535, n15536, n15537, n15538, n15539, n15540, n15541,
         n15542, n15543, n15544, n15545, n15546, n15547, n15548, n15549,
         n15550, n15551, n15552, n15553, n15554, n15555, n15556, n15557,
         n15558, n15559, n15560, n15561, n15562, n15563, n15564, n15565,
         n15566, n15567, n15568, n15569, n15570, n15571, n15572, n15573,
         n15574, n15575, n15576, n15577, n15578, n15579, n15580, n15581,
         n15582, n15583, n15584, n15585, n15586, n15587, n15588, n15589,
         n15590, n15591, n15592, n15593, n15594, n15595, n15596, n15597,
         n15598, n15599, n15600, n15601, n15602, n15603, n15604, n15605,
         n15606, n15607, n15608, n15609, n15610, n15611, n15612, n15613,
         n15614, n15615, n15616, n15617, n15618, n15619, n15620, n15621,
         n15622, n15623, n15624, n15625, n15626, n15627, n15628, n15629,
         n15630, n15631, n15632, n15633, n15634, n15635, n15636, n15637,
         n15638, n15639, n15640, n15641, n15642, n15643, n15644, n15645,
         n15646, n15647, n15648, n15649, n15650, n15651, n15652, n15653,
         n15654, n15655, n15656, n15657, n15658, n15659, n15660, n15661,
         n15662, n15663, n15664, n15665, n15666, n15667, n15668, n15669,
         n15670, n15671, n15672, n15673, n15674, n15675, n15676, n15677,
         n15678, n15679, n15680, n15681, n15682, n15683, n15684, n15685,
         n15686, n15687, n15688, n15689, n15690, n15691, n15692, n15693,
         n15694, n15695, n15696, n15697, n15698, n15699, n15700, n15701,
         n15702, n15703, n15704, n15705, n15706, n15707, n15708, n15709,
         n15710, n15711, n15712, n15713, n15714, n15715, n15716, n15717,
         n15718, n15719, n15720, n15721, n15722, n15723, n15724, n15725,
         n15726, n15727, n15728, n15729, n15730, n15731, n15732, n15733,
         n15734, n15735, n15736, n15737, n15738, n15739, n15740, n15741,
         n15742, n15743, n15744, n15745, n15746, n15747, n15748, n15749,
         n15750, n15751, n15752, n15753, n15754, n15755, n15756, n15757,
         n15758, n15759, n15760, n15761, n15762, n15763, n15764, n15765,
         n15766, n15767, n15768, n15769, n15770, n15771, n15772, n15773,
         n15774, n15775, n15776, n15777, n15778, n15779, n15780, n15781,
         n15782, n15783, n15784, n15785, n15786, n15787, n15788, n15789,
         n15790, n15791, n15792, n15793, n15794, n15795, n15796, n15797,
         n15798, n15799, n15800, n15801, n15802, n15803, n15804, n15805,
         n15806, n15807, n15808, n15809, n15810, n15811, n15812, n15813,
         n15814, n15815, n15816, n15817, n15818, n15819, n15820, n15821,
         n15822, n15823, n15824, n15825, n15826, n15827, n15828, n15829,
         n15830, n15831, n15832, n15833, n15834, n15835, n15836, n15837,
         n15838, n15839, n15840, n15841, n15842, n15843, n15844, n15845,
         n15846, n15847, n15848, n15849, n15850, n15851, n15852, n15853,
         n15854, n15855, n15856, n15857, n15858, n15859, n15860, n15861,
         n15862, n15863, n15864, n15865, n15866, n15867, n15868, n15869,
         n15870, n15871, n15872, n15873, n15874, n15875, n15876, n15877,
         n15878, n15879, n15880, n15881, n15882, n15883, n15884, n15885,
         n15886, n15887, n15888, n15889, n15890, n15891, n15892, n15893,
         n15894, n15895, n15896, n15897, n15898, n15899, n15900, n15901,
         n15902, n15903, n15904, n15905, n15906, n15907, n15908, n15909,
         n15910, n15911, n15912, n15913, n15914, n15915, n15916, n15917,
         n15918, n15919, n15920, n15921, n15922, n15923, n15924, n15925,
         n15926, n15927, n15928, n15929, n15930, n15931, n15932, n15933,
         n15934, n15935, n15936, n15937, n15938, n15939, n15940, n15941,
         n15942, n15943, n15944, n15945, n15946, n15947, n15948, n15949,
         n15950, n15951, n15952, n15953, n15954, n15955, n15956, n15957,
         n15958, n15959, n15960, n15961, n15962, n15963, n15964, n15965,
         n15966, n15967, n15968, n15969, n15970, n15971, n15972, n15973,
         n15974, n15975, n15976, n15977, n15978, n15979, n15980, n15981,
         n15982, n15983, n15984, n15985, n15986, n15987, n15988, n15989,
         n15990, n15991, n15992, n15993, n15994, n15995, n15996, n15997,
         n15998, n15999, n16000, n16001, n16002, n16003, n16004, n16005,
         n16006, n16007, n16008, n16009, n16010, n16011, n16012, n16013,
         n16014, n16015, n16016, n16017, n16018, n16019, n16020, n16021,
         n16022, n16023, n16024, n16025, n16026, n16027, n16028, n16029,
         n16030, n16031, n16032, n16033, n16034, n16035, n16036, n16037,
         n16038, n16039, n16040, n16041, n16042, n16043, n16044, n16045,
         n16046, n16047, n16048, n16049, n16050, n16051, n16052, n16053,
         n16054, n16055, n16056, n16057, n16058, n16059, n16060, n16061,
         n16062, n16063, n16064, n16065, n16066, n16067, n16068, n16069,
         n16070, n16071, n16072, n16073, n16074, n16075, n16076, n16077,
         n16078, n16079, n16080, n16081, n16082, n16083, n16084, n16085,
         n16086, n16087, n16088, n16089, n16090, n16091, n16092, n16093,
         n16094, n16095, n16096, n16097, n16098, n16099, n16100, n16101,
         n16102, n16103, n16104, n16105, n16106, n16107, n16108, n16109,
         n16110, n16111, n16112, n16113, n16114, n16115, n16116, n16117,
         n16118, n16119, n16120, n16121, n16122, n16123, n16124, n16125,
         n16126, n16127, n16128, n16129, n16130, n16131, n16132, n16133,
         n16134, n16135, n16136, n16137, n16138, n16139, n16140, n16141,
         n16142, n16143, n16144, n16145, n16146, n16147, n16148, n16149,
         n16150, n16151, n16152, n16153, n16154, n16155, n16156, n16157,
         n16158, n16159, n16160, n16161, n16162, n16163, n16164, n16165,
         n16166, n16167, n16168, n16169, n16170, n16171, n16172, n16173,
         n16174, n16175, n16176, n16177, n16178, n16179, n16180, n16181,
         n16182, n16183, n16184, n16185, n16186, n16187, n16188, n16189,
         n16190, n16191, n16192, n16193, n16194, n16195, n16196, n16197,
         n16198, n16199, n16200, n16201, n16202, n16203, n16204, n16205,
         n16206, n16207, n16208, n16209, n16210, n16211, n16212, n16213,
         n16214, n16215, n16216, n16217, n16218, n16219, n16220, n16221,
         n16222, n16223, n16224, n16225, n16226, n16227, n16228, n16229,
         n16230, n16231, n16232, n16233, n16234, n16235, n16236, n16237,
         n16238, n16239, n16240, n16241, n16242, n16243, n16244, n16245,
         n16246, n16247, n16248, n16249, n16250, n16251, n16252, n16253,
         n16254, n16255, n16256, n16257, n16258, n16259, n16260, n16261,
         n16262, n16263, n16264, n16265, n16266, n16267, n16268, n16269,
         n16270, n16271, n16272, n16273, n16274, n16275, n16276, n16277,
         n16278, n16279, n16280, n16281, n16282, n16283, n16284, n16285,
         n16286, n16287, n16288, n16289, n16290, n16291, n16292, n16293,
         n16294, n16295, n16296, n16297, n16298, n16299, n16300, n16301,
         n16302, n16303, n16304, n16305, n16306, n16307, n16308, n16309,
         n16310, n16311, n16312, n16313, n16314, n16315, n16316, n16317,
         n16318, n16319, n16320, n16321, n16322, n16323, n16324, n16325,
         n16326, n16327, n16328, n16329, n16330, n16331, n16332, n16333,
         n16334, n16335, n16336, n16337, n16338, n16339, n16340, n16341,
         n16342, n16343, n16344, n16345, n16346, n16347, n16348, n16349,
         n16350, n16351, n16352, n16353, n16354, n16355, n16356, n16357,
         n16358, n16359, n16360, n16361, n16362, n16363, n16364, n16365,
         n16366, n16367, n16368, n16369, n16370, n16371, n16372, n16373,
         n16374, n16375, n16376, n16377, n16378, n16379, n16380, n16381,
         n16382, n16383, n16384, n16385, n16386, n16387, n16388, n16389,
         n16390, n16391, n16392, n16393, n16394, n16395, n16396, n16397,
         n16398, n16399, n16400, n16401, n16402, n16403, n16404, n16405,
         n16406, n16407, n16408, n16409, n16410, n16411, n16412, n16413,
         n16414, n16415, n16416, n16417, n16418, n16419, n16420, n16421,
         n16422, n16423, n16424, n16425, n16426, n16427, n16428, n16429,
         n16430, n16431, n16432, n16433, n16434, n16435, n16436, n16437,
         n16438, n16439, n16440, n16441, n16442, n16443, n16444, n16445,
         n16446, n16447, n16448, n16449, n16450, n16451, n16452, n16453,
         n16454, n16455, n16456, n16457, n16458, n16459, n16460, n16461,
         n16462, n16463, n16464, n16465, n16466, n16467, n16468, n16469,
         n16470, n16471, n16472, n16473, n16474, n16475, n16476, n16477,
         n16478, n16479, n16480, n16481, n16482, n16483, n16484, n16485,
         n16486, n16487, n16488, n16489, n16490, n16491, n16492, n16493,
         n16494, n16495, n16496, n16497, n16498, n16499, n16500, n16501,
         n16502, n16503, n16504, n16505, n16506, n16507, n16508, n16509,
         n16510, n16511, n16512, n16513, n16514, n16515, n16516, n16517,
         n16518, n16519, n16520, n16521, n16522, n16523, n16524, n16525,
         n16526, n16527, n16528, n16529, n16530, n16531, n16532, n16533,
         n16534, n16535, n16536, n16537, n16538, n16539, n16540, n16541,
         n16542, n16543, n16544, n16545, n16546, n16547, n16548, n16549,
         n16550, n16551, n16552, n16553, n16554, n16555, n16556, n16557,
         n16558, n16559, n16560, n16561, n16562, n16563, n16564, n16565,
         n16566, n16567, n16568, n16569, n16570, n16571, n16572, n16573,
         n16574, n16575, n16576, n16577, n16578, n16579, n16580, n16581,
         n16582, n16583, n16584, n16585, n16586, n16587, n16588, n16589,
         n16590, n16591, n16592, n16593, n16594, n16595, n16596, n16597,
         n16598, n16599, n16600, n16601, n16602, n16603, n16604, n16605,
         n16606, n16607, n16608, n16609, n16610, n16611, n16612, n16613,
         n16614, n16615, n16616, n16617, n16618, n16619, n16620, n16621,
         n16622, n16623, n16624, n16625, n16626, n16627, n16628, n16629,
         n16630, n16631, n16632, n16633, n16634, n16635, n16636, n16637,
         n16638, n16639, n16640, n16641, n16642, n16643, n16644, n16645,
         n16646, n16647, n16648, n16649, n16650, n16651, n16652, n16653,
         n16654, n16655, n16656, n16657, n16658, n16659, n16660, n16661,
         n16662, n16663, n16664, n16665, n16666, n16667, n16668, n16669,
         n16670, n16671, n16672, n16673, n16674, n16675, n16676, n16677,
         n16678, n16679, n16680, n16681, n16682, n16683, n16684, n16685,
         n16686, n16687, n16688, n16689, n16690, n16691, n16692, n16693,
         n16694, n16695, n16696, n16697, n16698, n16699, n16700, n16701,
         n16702, n16703, n16704, n16705, n16706, n16707, n16708, n16709,
         n16710, n16711, n16712, n16713, n16714, n16715, n16716, n16717,
         n16718, n16719, n16720, n16721, n16722, n16723, n16724, n16725,
         n16726, n16727, n16728, n16729, n16730, n16731, n16732, n16733,
         n16734, n16735, n16736, n16737, n16738, n16739, n16740, n16741,
         n16742, n16743, n16744, n16745, n16746, n16747, n16748, n16749,
         n16750, n16751, n16752, n16753, n16754, n16755, n16756, n16757,
         n16758, n16759, n16760, n16761, n16762, n16763, n16764, n16765,
         n16766, n16767, n16768, n16769, n16770, n16771, n16772, n16773,
         n16774, n16775, n16776, n16777, n16778, n16779, n16780, n16781,
         n16782, n16783, n16784, n16785, n16786, n16787, n16788, n16789,
         n16790, n16791, n16792, n16793, n16794, n16795, n16796, n16797,
         n16798, n16799, n16800, n16801, n16802, n16803, n16804, n16805,
         n16806, n16807, n16808, n16809, n16810, n16811, n16812, n16813,
         n16814, n16815, n16816, n16817, n16818, n16819, n16820, n16821,
         n16822, n16823, n16824, n16825, n16826, n16827, n16828, n16829,
         n16830, n16831, n16832, n16833, n16834, n16835, n16836, n16837,
         n16838, n16839, n16840, n16841, n16842, n16843, n16844, n16845,
         n16846, n16847, n16848, n16849, n16850, n16851, n16852, n16853,
         n16854, n16855, n16856, n16857, n16858, n16859, n16860, n16861,
         n16862, n16863, n16864, n16865, n16866, n16867, n16868, n16869,
         n16870, n16871, n16872, n16873, n16874, n16875, n16876, n16877,
         n16878, n16879, n16880, n16881, n16882, n16883, n16884, n16885,
         n16886, n16887, n16888, n16889, n16890, n16891, n16892, n16893,
         n16894, n16895, n16896, n16897, n16898, n16899, n16900, n16901,
         n16902, n16903, n16904, n16905, n16906, n16907, n16908, n16909,
         n16910, n16911, n16912, n16913, n16914, n16915, n16916, n16917,
         n16918, n16919, n16920, n16921, n16922, n16923, n16924, n16925,
         n16926, n16927, n16928, n16929, n16930, n16931, n16932, n16933,
         n16934, n16935, n16936, n16937, n16938, n16939, n16940, n16941,
         n16942, n16943, n16944, n16945, n16946, n16947, n16948, n16949,
         n16950, n16951, n16952, n16953, n16954, n16955, n16956, n16957,
         n16958, n16959, n16960, n16961, n16962, n16963, n16964, n16965,
         n16966, n16967, n16968, n16969, n16970, n16971, n16972, n16973,
         n16974, n16975, n16976, n16977, n16978, n16979, n16980, n16981,
         n16982, n16983, n16984, n16985, n16986, n16987, n16988, n16989,
         n16990, n16991, n16992, n16993, n16994, n16995, n16996, n16997,
         n16998, n16999, n17000, n17001, n17002, n17003, n17004, n17005,
         n17006, n17007, n17008, n17009, n17010, n17011, n17012, n17013,
         n17014, n17015, n17016, n17017, n17018, n17019, n17020, n17021,
         n17022, n17023, n17024, n17025, n17026, n17027, n17028, n17029,
         n17030, n17031, n17032, n17033, n17034, n17035, n17036, n17037,
         n17038, n17039, n17040, n17041, n17042, n17043, n17044, n17045,
         n17046, n17047, n17048, n17049, n17050, n17051, n17052, n17053,
         n17054, n17055, n17056, n17057, n17058, n17059, n17060, n17061,
         n17062, n17063, n17064, n17065, n17066, n17067, n17068, n17069,
         n17070, n17071, n17072, n17073, n17074, n17075, n17076, n17077,
         n17078, n17079, n17080, n17081, n17082, n17083, n17084, n17085,
         n17086, n17087, n17088, n17089, n17090, n17091, n17092, n17093,
         n17094, n17095, n17096, n17097, n17098, n17099, n17100, n17101,
         n17102, n17103, n17104, n17105, n17106, n17107, n17108, n17109,
         n17110, n17111, n17112, n17113, n17114, n17115, n17116, n17117,
         n17118, n17119, n17120, n17121, n17122, n17123, n17124, n17125,
         n17126, n17127, n17128, n17129, n17130, n17131, n17132, n17133,
         n17134, n17135, n17136, n17137, n17138, n17139, n17140, n17141,
         n17142, n17143, n17144, n17145, n17146, n17147, n17148, n17149,
         n17150, n17151, n17152, n17153, n17154, n17155, n17156, n17157,
         n17158, n17159, n17160, n17161, n17162, n17163, n17164, n17165,
         n17166, n17167, n17168, n17169, n17170, n17171, n17172, n17173,
         n17174, n17175, n17176, n17177, n17178, n17179, n17180, n17181,
         n17182, n17183, n17184, n17185, n17186, n17187, n17188, n17189,
         n17190, n17191, n17192, n17193, n17194, n17195, n17196, n17197,
         n17198, n17199, n17200, n17201, n17202, n17203, n17204, n17205,
         n17206, n17207, n17208, n17209, n17210, n17211, n17212, n17213,
         n17214, n17215, n17216, n17217, n17218, n17219, n17220, n17221,
         n17222, n17223, n17224, n17225, n17226, n17227, n17228, n17229,
         n17230, n17231, n17232, n17233, n17234, n17235, n17236, n17237,
         n17238, n17239, n17240, n17241, n17242, n17243, n17244, n17245,
         n17246, n17247, n17248, n17249, n17250, n17251, n17252, n17253,
         n17254, n17255, n17256, n17257, n17258, n17259, n17260, n17261,
         n17262, n17263, n17264, n17265, n17266, n17267, n17268, n17269,
         n17270, n17271, n17272, n17273, n17274, n17275, n17276, n17277,
         n17278, n17279, n17280, n17281, n17282, n17283, n17284, n17285,
         n17286, n17287, n17288, n17289, n17290, n17291, n17292, n17293,
         n17294, n17295, n17296, n17297, n17298, n17299, n17300, n17301,
         n17302, n17303, n17304, n17305, n17306, n17307, n17308, n17309,
         n17310, n17311, n17312, n17313, n17314, n17315, n17316, n17317,
         n17318, n17319, n17320, n17321, n17322, n17323, n17324, n17325,
         n17326, n17327, n17328, n17329, n17330, n17331, n17332, n17333,
         n17334, n17335, n17336, n17337, n17338, n17339, n17340, n17341,
         n17342, n17343, n17344, n17345, n17346, n17347, n17348, n17349,
         n17350, n17351, n17352, n17353, n17354, n17355, n17356, n17357,
         n17358, n17359, n17360, n17361, n17362, n17363, n17364, n17365,
         n17366, n17367, n17368, n17369, n17370, n17371, n17372, n17373,
         n17374, n17375, n17376, n17377, n17378, n17379, n17380, n17381,
         n17382, n17383, n17384, n17385, n17386, n17387, n17388, n17389,
         n17390, n17391, n17392, n17393, n17394, n17395, n17396, n17397,
         n17398, n17399, n17400, n17401, n17402, n17403, n17404, n17405,
         n17406, n17407, n17408, n17409, n17410, n17411, n17412, n17413,
         n17414, n17415, n17416, n17417, n17418, n17419, n17420, n17421,
         n17422, n17423, n17424, n17425, n17426, n17427, n17428, n17429,
         n17430, n17431, n17432, n17433, n17434, n17435, n17436, n17437,
         n17438, n17439, n17440, n17441, n17442, n17443, n17444, n17445,
         n17446, n17447, n17448, n17449, n17450, n17451, n17452, n17453,
         n17454, n17455, n17456, n17457, n17458, n17459, n17460, n17461,
         n17462, n17463, n17464, n17465, n17466, n17467, n17468, n17469,
         n17470, n17471, n17472, n17473, n17474, n17475, n17476, n17477,
         n17478, n17479, n17480, n17481, n17482, n17483, n17484, n17485,
         n17486, n17487, n17488, n17489, n17490, n17491, n17492, n17493,
         n17494, n17495, n17496, n17497, n17498, n17499, n17500, n17501,
         n17502, n17503, n17504, n17505, n17506, n17507, n17508, n17509,
         n17510, n17511, n17512, n17513, n17514, n17515, n17516, n17517,
         n17518, n17519, n17520, n17521, n17522, n17523, n17524, n17525,
         n17526, n17527, n17528, n17529, n17530, n17531, n17532, n17533,
         n17534, n17535, n17536, n17537, n17538, n17539, n17540, n17541,
         n17542, n17543, n17544, n17545, n17546, n17547, n17548, n17549,
         n17550, n17551, n17552, n17553, n17554, n17555, n17556, n17557,
         n17558, n17559, n17560, n17561, n17562, n17563, n17564, n17565,
         n17566, n17567, n17568, n17569, n17570, n17571, n17572, n17573,
         n17574, n17575, n17576, n17577, n17578, n17579, n17580, n17581,
         n17582, n17583, n17584, n17585, n17586, n17587, n17588, n17589,
         n17590, n17591, n17592, n17593, n17594, n17595, n17596, n17597,
         n17598, n17599, n17600, n17601, n17602, n17603, n17604, n17605,
         n17606, n17607, n17608, n17609, n17610, n17611, n17612, n17613,
         n17614, n17615, n17616, n17617, n17618, n17619, n17620, n17621,
         n17622, n17623, n17624, n17625, n17626, n17627, n17628, n17629,
         n17630, n17631, n17632, n17633, n17634, n17635, n17636, n17637,
         n17638, n17639, n17640, n17641, n17642, n17643, n17644, n17645,
         n17646, n17647, n17648, n17649, n17650, n17651, n17652, n17653,
         n17654, n17655, n17656, n17657, n17658, n17659, n17660, n17661,
         n17662, n17663, n17664, n17665, n17666, n17667, n17668, n17669,
         n17670, n17671, n17672, n17673, n17674, n17675, n17676, n17677,
         n17678, n17679, n17680, n17681, n17682, n17683, n17684, n17685,
         n17686, n17687, n17688, n17689, n17690, n17691, n17692, n17693,
         n17694, n17695, n17696, n17697, n17698, n17699, n17700, n17701,
         n17702, n17703, n17704, n17705, n17706, n17707, n17708, n17709,
         n17710, n17711, n17712, n17713, n17714, n17715, n17716, n17717,
         n17718, n17719, n17720, n17721, n17722, n17723, n17724, n17725,
         n17726, n17727, n17728, n17729, n17730, n17731, n17732, n17733,
         n17734, n17735, n17736, n17737, n17738, n17739, n17740, n17741,
         n17742, n17743, n17744, n17745, n17746, n17747, n17748, n17749,
         n17750, n17751, n17752, n17753, n17754, n17755, n17756, n17757,
         n17758, n17759, n17760, n17761, n17762, n17763, n17764, n17765,
         n17766, n17767, n17768, n17769, n17770, n17771, n17772, n17773,
         n17774, n17775, n17776, n17777, n17778, n17779, n17780, n17781,
         n17782, n17783, n17784, n17785, n17786, n17787, n17788, n17789,
         n17790, n17791, n17792, n17793, n17794, n17795, n17796, n17797,
         n17798, n17799, n17800, n17801, n17802, n17803, n17804, n17805,
         n17806, n17807, n17808, n17809, n17810, n17811, n17812, n17813,
         n17814, n17815, n17816, n17817, n17818, n17819, n17820, n17821,
         n17822, n17823, n17824, n17825, n17826, n17827, n17828, n17829,
         n17830, n17831, n17832, n17833, n17834, n17835, n17836, n17837,
         n17838, n17839, n17840, n17841, n17842, n17843, n17844, n17845,
         n17846, n17847, n17848, n17849, n17850, n17851, n17852, n17853,
         n17854, n17855, n17856, n17857, n17858, n17859, n17860, n17861,
         n17862, n17863, n17864, n17865, n17866, n17867, n17868, n17869,
         n17870, n17871, n17872, n17873, n17874, n17875, n17876, n17877,
         n17878, n17879, n17880, n17881, n17882, n17883, n17884, n17885,
         n17886, n17887, n17888, n17889, n17890, n17891, n17892, n17893,
         n17894, n17895, n17896, n17897, n17898, n17899, n17900, n17901,
         n17902, n17903, n17904, n17905, n17906, n17907, n17908, n17909,
         n17910, n17911, n17912, n17913, n17914, n17915, n17916, n17917,
         n17918, n17919, n17920, n17921, n17922, n17923, n17924, n17925,
         n17926, n17927, n17928, n17929, n17930, n17931, n17932, n17933,
         n17934, n17935, n17936, n17937, n17938, n17939, n17940, n17941,
         n17942, n17943, n17944, n17945, n17946, n17947, n17948, n17949,
         n17950, n17951, n17952, n17953, n17954, n17955, n17956, n17957,
         n17958, n17959, n17960, n17961, n17962, n17963, n17964, n17965,
         n17966, n17967, n17968, n17969, n17970, n17971, n17972, n17973,
         n17974, n17975, n17976, n17977, n17978, n17979, n17980, n17981,
         n17982, n17983, n17984, n17985, n17986, n17987, n17988, n17989,
         n17990, n17991, n17992, n17993, n17994, n17995, n17996, n17997,
         n17998, n17999, n18000, n18001, n18002, n18003, n18004, n18005,
         n18006, n18007, n18008, n18009, n18010, n18011, n18012, n18013,
         n18014, n18015, n18016, n18017, n18018, n18019, n18020, n18021,
         n18022, n18023, n18024, n18025, n18026, n18027, n18028, n18029,
         n18030, n18031, n18032, n18033, n18034, n18035, n18036, n18037,
         n18038, n18039, n18040, n18041, n18042, n18043, n18044, n18045,
         n18046, n18047, n18048, n18049, n18050, n18051, n18052, n18053,
         n18054, n18055, n18056, n18057, n18058, n18059, n18060, n18061,
         n18062, n18063, n18064, n18065, n18066, n18067, n18068, n18069,
         n18070, n18071, n18072, n18073, n18074, n18075, n18076, n18077,
         n18078, n18079, n18080, n18081, n18082, n18083, n18084, n18085,
         n18086, n18087, n18088, n18089, n18090, n18091, n18092, n18093,
         n18094, n18095, n18096, n18097, n18098, n18099, n18100, n18101,
         n18102, n18103, n18104, n18105, n18106, n18107, n18108, n18109,
         n18110, n18111, n18112, n18113, n18114, n18115, n18116, n18117,
         n18118, n18119, n18120, n18121, n18122, n18123, n18124, n18125,
         n18126, n18127, n18128, n18129, n18130, n18131, n18132, n18133,
         n18134, n18135, n18136, n18137, n18138, n18139, n18140, n18141,
         n18142, n18143, n18144, n18145, n18146, n18147, n18148, n18149,
         n18150, n18151, n18152, n18153, n18154, n18155, n18156, n18157,
         n18158, n18159, n18160, n18161, n18162, n18163, n18164, n18165,
         n18166, n18167, n18168, n18169, n18170, n18171, n18172, n18173,
         n18174, n18175, n18176, n18177, n18178, n18179, n18180, n18181,
         n18182, n18183, n18184, n18185, n18186, n18187, n18188, n18189,
         n18190, n18191, n18192, n18193, n18194, n18195, n18196, n18197,
         n18198, n18199, n18200, n18201, n18202, n18203, n18204, n18205,
         n18206, n18207, n18208, n18209, n18210, n18211, n18212, n18213,
         n18214, n18215, n18216, n18217, n18218, n18219, n18220, n18221,
         n18222, n18223, n18224, n18225, n18226, n18227, n18228, n18229,
         n18230, n18231, n18232, n18233, n18234, n18235, n18236, n18237,
         n18238, n18239, n18240, n18241, n18242, n18243, n18244, n18245,
         n18246, n18247, n18248, n18249, n18250, n18251, n18252, n18253,
         n18254, n18255, n18256, n18257, n18258, n18259, n18260, n18261,
         n18262, n18263, n18264, n18265, n18266, n18267, n18268, n18269,
         n18270, n18271, n18272, n18273, n18274, n18275, n18276, n18277,
         n18278, n18279, n18280, n18281, n18282, n18283, n18284, n18285,
         n18286, n18287, n18288, n18289, n18290, n18291, n18292, n18293,
         n18294, n18295, n18296, n18297, n18298, n18299, n18300, n18301,
         n18302, n18303, n18304, n18305, n18306, n18307, n18308, n18309,
         n18310, n18311, n18312, n18313, n18314, n18315, n18316, n18317,
         n18318, n18319, n18320, n18321, n18322, n18323, n18324, n18325,
         n18326, n18327, n18328, n18329, n18330, n18331, n18332, n18333,
         n18334, n18335, n18336, n18337, n18338, n18339, n18340, n18341,
         n18342, n18343, n18344, n18345, n18346, n18347, n18348, n18349,
         n18350, n18351, n18352, n18353, n18354, n18355, n18356, n18357,
         n18358, n18359, n18360, n18361, n18362, n18363, n18364, n18365,
         n18366, n18367, n18368, n18369, n18370, n18371, n18372, n18373,
         n18374, n18375, n18376, n18377, n18378, n18379, n18380, n18381,
         n18382, n18383, n18384, n18385, n18386, n18387, n18388, n18389,
         n18390, n18391, n18392, n18393, n18394, n18395, n18396, n18397,
         n18398, n18399, n18400, n18401, n18402, n18403, n18404, n18405,
         n18406, n18407, n18408, n18409, n18410, n18411, n18412, n18413,
         n18414, n18415, n18416, n18417, n18418, n18419, n18420, n18421,
         n18422, n18423, n18424, n18425, n18426, n18427, n18428, n18429,
         n18430, n18431, n18432, n18433, n18434, n18435, n18436, n18437,
         n18438, n18439, n18440, n18441, n18442, n18443, n18444, n18445,
         n18446, n18447, n18448, n18449, n18450, n18451, n18452, n18453,
         n18454, n18455, n18456, n18457, n18458, n18459, n18460, n18461,
         n18462, n18463, n18464, n18465, n18466, n18467, n18468, n18469,
         n18470, n18471, n18472, n18473, n18474, n18475, n18476, n18477,
         n18478, n18479, n18480, n18481, n18482, n18483, n18484, n18485,
         n18486, n18487, n18488, n18489, n18490, n18491, n18492, n18493,
         n18494, n18495, n18496, n18497, n18498, n18499, n18500, n18501,
         n18502, n18503, n18504, n18505, n18506, n18507, n18508, n18509,
         n18510, n18511, n18512, n18513, n18514, n18515, n18516, n18517,
         n18518, n18519, n18520, n18521, n18522, n18523, n18524, n18525,
         n18526, n18527, n18528, n18529, n18530, n18531, n18532, n18533,
         n18534, n18535, n18536, n18537, n18538, n18539, n18540, n18541,
         n18542, n18543, n18544, n18545, n18546, n18547, n18548, n18549,
         n18550, n18551, n18552, n18553, n18554, n18555, n18556, n18557,
         n18558, n18559, n18560, n18561, n18562, n18563, n18564, n18565,
         n18566, n18567, n18568, n18569, n18570, n18571, n18572, n18573,
         n18574, n18575, n18576, n18577, n18578, n18579, n18580, n18581,
         n18582, n18583, n18584, n18585, n18586, n18587, n18588, n18589,
         n18590, n18591, n18592, n18593, n18594, n18595, n18596, n18597,
         n18598, n18599, n18600, n18601, n18602, n18603, n18604, n18605,
         n18606, n18607, n18608, n18609, n18610, n18611, n18612, n18613,
         n18614, n18615, n18616, n18617, n18618, n18619, n18620, n18621,
         n18622, n18623, n18624, n18625, n18626, n18627, n18628, n18629,
         n18630, n18631, n18632, n18633, n18634, n18635, n18636, n18637,
         n18638, n18639, n18640, n18641, n18642, n18643, n18644, n18645,
         n18646, n18647, n18648, n18649, n18650, n18651, n18652, n18653,
         n18654, n18655, n18656, n18657, n18658, n18659, n18660, n18661,
         n18662, n18663, n18664, n18665, n18666, n18667, n18668, n18669,
         n18670, n18671, n18672, n18673, n18674, n18675, n18676, n18677,
         n18678, n18679, n18680, n18681, n18682, n18683, n18684, n18685,
         n18686, n18687, n18688, n18689, n18690, n18691, n18692, n18693,
         n18694, n18695, n18696, n18697, n18698, n18699, n18700, n18701,
         n18702, n18703, n18704, n18705, n18706, n18707, n18708, n18709,
         n18710, n18711, n18712, n18713, n18714, n18715, n18716, n18717,
         n18718, n18719, n18720, n18721, n18722, n18723, n18724, n18725,
         n18726, n18727, n18728, n18729, n18730, n18731, n18732, n18733,
         n18734, n18735, n18736, n18737, n18738, n18739, n18740, n18741,
         n18742, n18743, n18744, n18745, n18746, n18747, n18748, n18749,
         n18750, n18751, n18752, n18753, n18754, n18755, n18756, n18757,
         n18758, n18759, n18760, n18761, n18762, n18763, n18764, n18765,
         n18766, n18767, n18768, n18769, n18770, n18771, n18772, n18773,
         n18774, n18775, n18776, n18777, n18778, n18779, n18780, n18781,
         n18782, n18783, n18784, n18785, n18786, n18787, n18788, n18789,
         n18790, n18791, n18792, n18793, n18794, n18795, n18796, n18797,
         n18798, n18799, n18800, n18801, n18802, n18803, n18804, n18805,
         n18806, n18807, n18808, n18809, n18810, n18811, n18812, n18813,
         n18814, n18815, n18816, n18817, n18818, n18819, n18820, n18821,
         n18822, n18823, n18824, n18825, n18826, n18827, n18828, n18829,
         n18830, n18831, n18832, n18833, n18834, n18835, n18836, n18837,
         n18838, n18839, n18840, n18841, n18842, n18843, n18844, n18845,
         n18846, n18847, n18848, n18849, n18850, n18851, n18852, n18853,
         n18854, n18855, n18856, n18857, n18858, n18859, n18860, n18861,
         n18862, n18863, n18864, n18865, n18866, n18867, n18868, n18869,
         n18870, n18871, n18872, n18873, n18874, n18875, n18876, n18877,
         n18878, n18879, n18880, n18881, n18882, n18883, n18884, n18885,
         n18886, n18887, n18888, n18889, n18890, n18891, n18892, n18893,
         n18894, n18895, n18896, n18897, n18898, n18899, n18900, n18901,
         n18902, n18903, n18904, n18905, n18906, n18907, n18908, n18909,
         n18910, n18911, n18912, n18913, n18914, n18915, n18916, n18917,
         n18918, n18919, n18920, n18921, n18922, n18923, n18924, n18925,
         n18926, n18927, n18928, n18929, n18930, n18931, n18932, n18933,
         n18934, n18935, n18936, n18937, n18938, n18939, n18940, n18941,
         n18942, n18943, n18944, n18945, n18946, n18947, n18948, n18949,
         n18950, n18951, n18952, n18953, n18954, n18955, n18956, n18957,
         n18958, n18959, n18960, n18961, n18962, n18963, n18964, n18965,
         n18966, n18967, n18968, n18969, n18970, n18971, n18972, n18973,
         n18974, n18975, n18976, n18977, n18978, n18979, n18980, n18981,
         n18982, n18983, n18984, n18985, n18986, n18987, n18988, n18989,
         n18990, n18991, n18992, n18993, n18994, n18995, n18996, n18997,
         n18998, n18999, n19000, n19001, n19002, n19003, n19004, n19005,
         n19006, n19007, n19008, n19009, n19010, n19011, n19012, n19013,
         n19014, n19015, n19016, n19017, n19018, n19019, n19020, n19021,
         n19022, n19023, n19024, n19025, n19026, n19027, n19028, n19029,
         n19030, n19031, n19032, n19033, n19034, n19035, n19036, n19037,
         n19038, n19039, n19040, n19041, n19042, n19043, n19044, n19045,
         n19046, n19047, n19048, n19049, n19050, n19051, n19052, n19053,
         n19054, n19055, n19056, n19057, n19058, n19059, n19060, n19061,
         n19062, n19063, n19064, n19065, n19066, n19067, n19068, n19069,
         n19070, n19071, n19072, n19073, n19074, n19075, n19076, n19077,
         n19078, n19079, n19080, n19081, n19082, n19083, n19084, n19085,
         n19086, n19087, n19088, n19089, n19090, n19091, n19092, n19093,
         n19094, n19095, n19096, n19097, n19098, n19099, n19100, n19101,
         n19102, n19103, n19104, n19105, n19106, n19107, n19108, n19109,
         n19110, n19111, n19112, n19113, n19114, n19115, n19116, n19117,
         n19118, n19119, n19120, n19121, n19122, n19123, n19124, n19125,
         n19126, n19127, n19128, n19129, n19130, n19131, n19132, n19133,
         n19134, n19135, n19136, n19137, n19138, n19139, n19140, n19141,
         n19142, n19143, n19144, n19145, n19146, n19147, n19148, n19149,
         n19150, n19151, n19152, n19153, n19154, n19155, n19156, n19157,
         n19158, n19159, n19160, n19161, n19162, n19163, n19164, n19165,
         n19166, n19167, n19168, n19169, n19170, n19171, n19172, n19173,
         n19174, n19175, n19176, n19177, n19178, n19179, n19180, n19181,
         n19182, n19183, n19184, n19185, n19186, n19187, n19188, n19189,
         n19190, n19191, n19192, n19193, n19194, n19195, n19196, n19197,
         n19198, n19199, n19200, n19201, n19202, n19203, n19204, n19205,
         n19206, n19207, n19208, n19209, n19210, n19211, n19212, n19213,
         n19214, n19215, n19216, n19217, n19218, n19219, n19220, n19221,
         n19222, n19223, n19224, n19225, n19226, n19227, n19228, n19229,
         n19230, n19231, n19232, n19233, n19234, n19235, n19236, n19237,
         n19238, n19239, n19240, n19241, n19242, n19243, n19244, n19245,
         n19246, n19247, n19248, n19249, n19250, n19251, n19252, n19253,
         n19254, n19255, n19256, n19257, n19258, n19259, n19260, n19261,
         n19262, n19263, n19264, n19265, n19266, n19267, n19268, n19269,
         n19270, n19271, n19272, n19273, n19274, n19275, n19276, n19277,
         n19278, n19279, n19280, n19281, n19282, n19283, n19284, n19285,
         n19286, n19287, n19288, n19289, n19290, n19291, n19292, n19293,
         n19294, n19295, n19296, n19297, n19298, n19299, n19300, n19301,
         n19302, n19303, n19304, n19305, n19306, n19307, n19308, n19309,
         n19310, n19311, n19312, n19313, n19314, n19315, n19316, n19317,
         n19318, n19319, n19320, n19321, n19322, n19323, n19324, n19325,
         n19326, n19327, n19328, n19329, n19330, n19331, n19332, n19333,
         n19334, n19335, n19336, n19337, n19338, n19339, n19340, n19341,
         n19342, n19343, n19344, n19345, n19346, n19347, n19348, n19349,
         n19350, n19351, n19352, n19353, n19354, n19355, n19356, n19357,
         n19358, n19359, n19360, n19361, n19362, n19363, n19364, n19365,
         n19366, n19367, n19368, n19369, n19370, n19371, n19372, n19373,
         n19374, n19375, n19376, n19377, n19378, n19379, n19380, n19381,
         n19382, n19383, n19384, n19385, n19386, n19387, n19388, n19389,
         n19390, n19391, n19392, n19393, n19394, n19395, n19396, n19397,
         n19398, n19399, n19400, n19401, n19402, n19403, n19404, n19405,
         n19406, n19407, n19408, n19409, n19410, n19411, n19412, n19413,
         n19414, n19415, n19416, n19417, n19418, n19419, n19420, n19421,
         n19422, n19423, n19424, n19425, n19426, n19427, n19428, n19429,
         n19430, n19431, n19432, n19433, n19434, n19435, n19436, n19437,
         n19438, n19439, n19440, n19441, n19442, n19443, n19444, n19445,
         n19446, n19447, n19448, n19449, n19450, n19451, n19452, n19453,
         n19454, n19455, n19456, n19457, n19458, n19459, n19460, n19461,
         n19462, n19463, n19464, n19465, n19466, n19467, n19468, n19469,
         n19470, n19471, n19472, n19473, n19474, n19475, n19476, n19477,
         n19478, n19479, n19480, n19481, n19482, n19483, n19484, n19485,
         n19486, n19487, n19488, n19489, n19490, n19491, n19492, n19493,
         n19494, n19495, n19496, n19497, n19498, n19499, n19500, n19501,
         n19502, n19503, n19504, n19505, n19506, n19507, n19508, n19509,
         n19510, n19511, n19512, n19513, n19514, n19515, n19516, n19517,
         n19518, n19519, n19520, n19521, n19522, n19523, n19524, n19525,
         n19526, n19527, n19528, n19529, n19530, n19531, n19532, n19533,
         n19534, n19535, n19536, n19537, n19538, n19539, n19540, n19541,
         n19542, n19543, n19544, n19545, n19546, n19547, n19548, n19549,
         n19550, n19551, n19552, n19553, n19554, n19555, n19556, n19557,
         n19558, n19559, n19560, n19561, n19562, n19563, n19564, n19565,
         n19566, n19567, n19568, n19569, n19570, n19571, n19572, n19573,
         n19574, n19575, n19576, n19577, n19578, n19579, n19580, n19581,
         n19582, n19583, n19584, n19585, n19586, n19587, n19588, n19589,
         n19590, n19591, n19592, n19593, n19594, n19595, n19596, n19597,
         n19598, n19599, n19600, n19601, n19602, n19603, n19604, n19605,
         n19606, n19607, n19608, n19609, n19610, n19611, n19612, n19613,
         n19614, n19615, n19616, n19617, n19618, n19619, n19620, n19621,
         n19622, n19623, n19624, n19625, n19626, n19627, n19628, n19629,
         n19630, n19631, n19632, n19633, n19634, n19635, n19636, n19637,
         n19638, n19639, n19640, n19641, n19642, n19643, n19644, n19645,
         n19646, n19647, n19648, n19649, n19650, n19651, n19652, n19653,
         n19654, n19655, n19656, n19657, n19658, n19659, n19660, n19661,
         n19662, n19663, n19664, n19665, n19666, n19667, n19668, n19669,
         n19670, n19671, n19672, n19673, n19674, n19675, n19676, n19677,
         n19678, n19679, n19680, n19681, n19682, n19683, n19684, n19685,
         n19686, n19687, n19688, n19689, n19690, n19691, n19692, n19693,
         n19694, n19695, n19696, n19697, n19698, n19699, n19700, n19701,
         n19702, n19703, n19704, n19705, n19706, n19707, n19708, n19709,
         n19710, n19711, n19712, n19713, n19714, n19715, n19716, n19717,
         n19718, n19719, n19720, n19721, n19722, n19723, n19724, n19725,
         n19726, n19727, n19728, n19729, n19730, n19731, n19732, n19733,
         n19734, n19735, n19736, n19737, n19738, n19739, n19740, n19741,
         n19742, n19743, n19744, n19745, n19746, n19747, n19748, n19749,
         n19750, n19751, n19752, n19753, n19754, n19755, n19756, n19757,
         n19758, n19759, n19760, n19761, n19762, n19763, n19764, n19765,
         n19766, n19767, n19768, n19769, n19770, n19771, n19772, n19773,
         n19774, n19775, n19776, n19777, n19778, n19779, n19780, n19781,
         n19782, n19783, n19784, n19785, n19786, n19787, n19788, n19789,
         n19790, n19791, n19792, n19793, n19794, n19795, n19796, n19797,
         n19798, n19799, n19800, n19801, n19802, n19803, n19804, n19805,
         n19806, n19807, n19808, n19809, n19810, n19811, n19812, n19813,
         n19814, n19815, n19816, n19817, n19818, n19819, n19820, n19821,
         n19822, n19823, n19824, n19825, n19826, n19827, n19828, n19829,
         n19830, n19831, n19832, n19833, n19834, n19835, n19836, n19837,
         n19838, n19839, n19840, n19841, n19842, n19843, n19844, n19845,
         n19846, n19847, n19848, n19849, n19850, n19851, n19852, n19853,
         n19854, n19855, n19856, n19857, n19858, n19859, n19860, n19861,
         n19862, n19863, n19864, n19865, n19866, n19867, n19868, n19869,
         n19870, n19871, n19872, n19873, n19874, n19875, n19876, n19877,
         n19878, n19879, n19880, n19881, n19882, n19883, n19884, n19885,
         n19886, n19887, n19888, n19889, n19890, n19891, n19892, n19893,
         n19894, n19895, n19896, n19897, n19898, n19899, n19900, n19901,
         n19902, n19903, n19904, n19905, n19906, n19907, n19908, n19909,
         n19910, n19911, n19912, n19913, n19914, n19915, n19916, n19917,
         n19918, n19919, n19920, n19921, n19922, n19923, n19924, n19925,
         n19926, n19927, n19928, n19929, n19930, n19931, n19932, n19933,
         n19934, n19935, n19936, n19937, n19938, n19939, n19940, n19941,
         n19942, n19943, n19944, n19945, n19946, n19947, n19948, n19949,
         n19950, n19951, n19952, n19953, n19954, n19955, n19956, n19957,
         n19958, n19959, n19960, n19961, n19962, n19963, n19964, n19965,
         n19966, n19967, n19968, n19969, n19970, n19971, n19972, n19973,
         n19974, n19975, n19976, n19977, n19978, n19979, n19980, n19981,
         n19982, n19983, n19984, n19985, n19986, n19987, n19988, n19989,
         n19990, n19991, n19992, n19993, n19994, n19995, n19996, n19997,
         n19998, n19999, n20000, n20001, n20002, n20003, n20004, n20005,
         n20006, n20007, n20008, n20009, n20010, n20011, n20012, n20013,
         n20014, n20015, n20016, n20017, n20018, n20019, n20020, n20021,
         n20022, n20023, n20024, n20025, n20026, n20027, n20028, n20029,
         n20030, n20031, n20032, n20033, n20034, n20035, n20036, n20037,
         n20038, n20039, n20040, n20041, n20042, n20043, n20044, n20045,
         n20046, n20047, n20048, n20049, n20050, n20051, n20052, n20053,
         n20054, n20055, n20056, n20057, n20058, n20059, n20060, n20061,
         n20062, n20063, n20064, n20065, n20066, n20067, n20068, n20069,
         n20070, n20071, n20072, n20073, n20074, n20075, n20076, n20077,
         n20078, n20079, n20080, n20081, n20082, n20083, n20084, n20085,
         n20086, n20087, n20088, n20089, n20090, n20091, n20092, n20093,
         n20094, n20095, n20096, n20097, n20098, n20099, n20100, n20101,
         n20102, n20103, n20104, n20105, n20106, n20107, n20108, n20109,
         n20110, n20111, n20112, n20113, n20114, n20115, n20116, n20117,
         n20118, n20119, n20120, n20121, n20122, n20123, n20124, n20125,
         n20126, n20127, n20128, n20129, n20130, n20131, n20132, n20133,
         n20134, n20135, n20136, n20137, n20138, n20139, n20140, n20141,
         n20142, n20143, n20144, n20145, n20146, n20147, n20148, n20149,
         n20150, n20151, n20152, n20153, n20154, n20155, n20156, n20157,
         n20158, n20159, n20160, n20161, n20162, n20163, n20164, n20165,
         n20166, n20167, n20168, n20169, n20170, n20171, n20172, n20173,
         n20174, n20175, n20176, n20177, n20178, n20179, n20180, n20181,
         n20182, n20183, n20184, n20185, n20186, n20187, n20188, n20189,
         n20190, n20191, n20192, n20193, n20194, n20195, n20196, n20197,
         n20198, n20199, n20200, n20201, n20202, n20203, n20204, n20205,
         n20206, n20207, n20208, n20209, n20210, n20211, n20212, n20213,
         n20214, n20215, n20216, n20217, n20218, n20219, n20220, n20221,
         n20222, n20223, n20224, n20225, n20226, n20227, n20228, n20229,
         n20230, n20231, n20232, n20233, n20234, n20235, n20236, n20237,
         n20238, n20239, n20240, n20241, n20242, n20243, n20244, n20245,
         n20246, n20247, n20248, n20249, n20250, n20251, n20252, n20253,
         n20254, n20255, n20256, n20257, n20258, n20259, n20260, n20261,
         n20262, n20263, n20264, n20265, n20266, n20267, n20268, n20269,
         n20270, n20271, n20272, n20273, n20274, n20275, n20276, n20277,
         n20278, n20279, n20280, n20281, n20282, n20283, n20284, n20285,
         n20286, n20287, n20288, n20289, n20290, n20291, n20292, n20293,
         n20294, n20295, n20296, n20297, n20298, n20299, n20300, n20301,
         n20302, n20303, n20304, n20305, n20306, n20307, n20308, n20309,
         n20310, n20311, n20312, n20313, n20314, n20315, n20316, n20317,
         n20318, n20319, n20320, n20321, n20322, n20323, n20324, n20325,
         n20326, n20327, n20328, n20329, n20330, n20331, n20332, n20333,
         n20334, n20335, n20336, n20337, n20338, n20339, n20340, n20341,
         n20342, n20343, n20344, n20345, n20346, n20347, n20348, n20349,
         n20350, n20351, n20352, n20353, n20354, n20355, n20356, n20357,
         n20358, n20359, n20360, n20361, n20362, n20363, n20364, n20365,
         n20366, n20367, n20368, n20369, n20370, n20371, n20372, n20373,
         n20374, n20375, n20376, n20377, n20378, n20379, n20380, n20381,
         n20382, n20383, n20384, n20385, n20386, n20387, n20388, n20389,
         n20390, n20391, n20392, n20393, n20394, n20395, n20396, n20397,
         n20398, n20399, n20400, n20401, n20402, n20403, n20404, n20405,
         n20406, n20407, n20408, n20409, n20410, n20411, n20412, n20413,
         n20414, n20415, n20416, n20417, n20418, n20419, n20420, n20421,
         n20422, n20423, n20424, n20425, n20426, n20427, n20428, n20429,
         n20430, n20431, n20432, n20433, n20434, n20435, n20436, n20437,
         n20438, n20439, n20440, n20441, n20442, n20443, n20444, n20445,
         n20446, n20447, n20448, n20449, n20450, n20451, n20452, n20453,
         n20454, n20455, n20456, n20457, n20458, n20459, n20460, n20461,
         n20462, n20463, n20464, n20465, n20466, n20467, n20468, n20469,
         n20470, n20471, n20472, n20473, n20474, n20475, n20476, n20477,
         n20478, n20479, n20480, n20481, n20482, n20483, n20484, n20485,
         n20486, n20487, n20488, n20489, n20490, n20491, n20492, n20493,
         n20494, n20495, n20496, n20497, n20498, n20499, n20500, n20501,
         n20502, n20503, n20504, n20505, n20506, n20507, n20508, n20509,
         n20510, n20511, n20512, n20513, n20514, n20515, n20516, n20517,
         n20518, n20519, n20520, n20521, n20522, n20523, n20524, n20525,
         n20526, n20527, n20528, n20529, n20530, n20531, n20532, n20533,
         n20534, n20535, n20536, n20537, n20538, n20539, n20540, n20541,
         n20542, n20543, n20544, n20545, n20546, n20547, n20548, n20549,
         n20550, n20551, n20552, n20553, n20554, n20555, n20556, n20557,
         n20558, n20559, n20560, n20561, n20562, n20563, n20564, n20565,
         n20566, n20567, n20568, n20569, n20570, n20571, n20572, n20573,
         n20574, n20575, n20576, n20577, n20578, n20579, n20580, n20581,
         n20582, n20583, n20584, n20585, n20586, n20587, n20588, n20589,
         n20590, n20591, n20592, n20593, n20594, n20595, n20596, n20597,
         n20598, n20599, n20600, n20601, n20602, n20603, n20604, n20605,
         n20606, n20607, n20608, n20609, n20610, n20611, n20612, n20613,
         n20614, n20615, n20616, n20617, n20618, n20619, n20620, n20621,
         n20622, n20623, n20624, n20625, n20626, n20627, n20628, n20629,
         n20630, n20631, n20632, n20633, n20634, n20635, n20636, n20637,
         n20638, n20639, n20640, n20641, n20642, n20643, n20644, n20645,
         n20646, n20647, n20648, n20649, n20650, n20651, n20652, n20653,
         n20654, n20655, n20656, n20657, n20658, n20659, n20660, n20661,
         n20662, n20663, n20664, n20665, n20666, n20667, n20668, n20669,
         n20670, n20671, n20672, n20673, n20674, n20675, n20676, n20677,
         n20678, n20679, n20680, n20681, n20682, n20683, n20684, n20685,
         n20686, n20687, n20688, n20689, n20690, n20691, n20692, n20693,
         n20694, n20695, n20696, n20697, n20698, n20699, n20700, n20701,
         n20702, n20703, n20704, n20705, n20706, n20707, n20708, n20709,
         n20710, n20711, n20712, n20713, n20714, n20715, n20716, n20717,
         n20718, n20719, n20720, n20721, n20722, n20723, n20724, n20725,
         n20726, n20727, n20728, n20729, n20730, n20731, n20732, n20733,
         n20734, n20735, n20736, n20737, n20738, n20739, n20740, n20741,
         n20742, n20743, n20744, n20745, n20746, n20747, n20748, n20749,
         n20750, n20751, n20752, n20753, n20754, n20755, n20756, n20757,
         n20758, n20759, n20760, n20761, n20762, n20763, n20764, n20765,
         n20766, n20767, n20768, n20769, n20770, n20771, n20772, n20773,
         n20774, n20775, n20776, n20777, n20778, n20779, n20780, n20781,
         n20782, n20783, n20784, n20785, n20786, n20787, n20788, n20789,
         n20790, n20791, n20792, n20793, n20794, n20795, n20796, n20797,
         n20798, n20799, n20800, n20801, n20802, n20803, n20804, n20805,
         n20806, n20807, n20808, n20809, n20810, n20811, n20812, n20813,
         n20814, n20815, n20816, n20817, n20818, n20819, n20820, n20821,
         n20822, n20823, n20824, n20825, n20826, n20827, n20828, n20829,
         n20830, n20831, n20832, n20833, n20834, n20835, n20836, n20837,
         n20838, n20839, n20840, n20841, n20842, n20843, n20844, n20845,
         n20846, n20847, n20848, n20849, n20850, n20851, n20852, n20853,
         n20854, n20855, n20856, n20857, n20858, n20859, n20860, n20861,
         n20862, n20863, n20864, n20865, n20866, n20867, n20868, n20869,
         n20870, n20871, n20872, n20873, n20874, n20875, n20876, n20877,
         n20878, n20879, n20880, n20881, n20882, n20883, n20884, n20885,
         n20886, n20887, n20888, n20889, n20890, n20891, n20892, n20893,
         n20894, n20895, n20896, n20897, n20898, n20899, n20900, n20901,
         n20902, n20903, n20904, n20905, n20906, n20907, n20908, n20909,
         n20910, n20911, n20912, n20913, n20914, n20915, n20916, n20917,
         n20918, n20919, n20920, n20921, n20922, n20923, n20924, n20925,
         n20926, n20927, n20928, n20929, n20930, n20931, n20932, n20933,
         n20934, n20935, n20936, n20937, n20938, n20939, n20940, n20941,
         n20942, n20943, n20944, n20945, n20946, n20947, n20948, n20949,
         n20950, n20951, n20952, n20953, n20954, n20955, n20956, n20957,
         n20958, n20959, n20960, n20961, n20962, n20963, n20964, n20965,
         n20966, n20967, n20968, n20969, n20970, n20971, n20972, n20973,
         n20974, n20975, n20976, n20977, n20978, n20979, n20980, n20981,
         n20982, n20983, n20984, n20985, n20986, n20987, n20988, n20989,
         n20990, n20991, n20992, n20993, n20994, n20995, n20996, n20997,
         n20998, n20999, n21000, n21001, n21002, n21003, n21004, n21005,
         n21006, n21007, n21008, n21009, n21010, n21011, n21012, n21013,
         n21014, n21015, n21016, n21017, n21018, n21019, n21020, n21021,
         n21022, n21023, n21024, n21025, n21026, n21027, n21028, n21029,
         n21030, n21031, n21032, n21033, n21034, n21035, n21036, n21037,
         n21038, n21039, n21040, n21041, n21042, n21043, n21044, n21045,
         n21046, n21047, n21048, n21049, n21050, n21051, n21052, n21053,
         n21054, n21055, n21056, n21057, n21058, n21059, n21060, n21061,
         n21062, n21063, n21064, n21065, n21066, n21067, n21068, n21069,
         n21070, n21071, n21072, n21073, n21074, n21075, n21076, n21077,
         n21078, n21079, n21080, n21081, n21082, n21083, n21084, n21085,
         n21086, n21087, n21088, n21089, n21090, n21091, n21092, n21093,
         n21094, n21095, n21096, n21097, n21098, n21099, n21100, n21101,
         n21102, n21103, n21104, n21105, n21106, n21107, n21108, n21109,
         n21110, n21111, n21112, n21113, n21114, n21115, n21116, n21117,
         n21118, n21119, n21120, n21121, n21122, n21123, n21124, n21125,
         n21126, n21127, n21128, n21129, n21130, n21131, n21132, n21133,
         n21134, n21135, n21136, n21137, n21138, n21139, n21140, n21141,
         n21142, n21143, n21144, n21145, n21146, n21147, n21148, n21149,
         n21150, n21151, n21152, n21153, n21154, n21155, n21156, n21157,
         n21158, n21159, n21160, n21161, n21162, n21163, n21164, n21165,
         n21166, n21167, n21168, n21169, n21170, n21171, n21172, n21173,
         n21174, n21175, n21176, n21177, n21178, n21179, n21180, n21181,
         n21182, n21183, n21184, n21185, n21186, n21187, n21188, n21189,
         n21190, n21191, n21192, n21193, n21194, n21195, n21196, n21197,
         n21198, n21199, n21200, n21201, n21202, n21203, n21204, n21205,
         n21206, n21207, n21208, n21209, n21210, n21211, n21212, n21213,
         n21214, n21215, n21216, n21217, n21218, n21219, n21220, n21221,
         n21222, n21223, n21224, n21225, n21226, n21227, n21228, n21229,
         n21230, n21231, n21232, n21233, n21234, n21235, n21236, n21237,
         n21238, n21239, n21240, n21241, n21242, n21243, n21244, n21245,
         n21246, n21247, n21248, n21249, n21250, n21251, n21252, n21253,
         n21254, n21255, n21256, n21257, n21258, n21259, n21260, n21261,
         n21262, n21263, n21264, n21265, n21266, n21267, n21268, n21269,
         n21270, n21271, n21272, n21273, n21274, n21275, n21276, n21277,
         n21278, n21279, n21280, n21281, n21282, n21283, n21284, n21285,
         n21286, n21287, n21288, n21289, n21290, n21291, n21292, n21293,
         n21294, n21295, n21296, n21297, n21298, n21299, n21300, n21301,
         n21302, n21303, n21304, n21305, n21306, n21307, n21308, n21309,
         n21310, n21311, n21312, n21313, n21314, n21315, n21316, n21317,
         n21318, n21319, n21320, n21321, n21322, n21323, n21324, n21325,
         n21326, n21327, n21328, n21329, n21330, n21331, n21332, n21333,
         n21334, n21335, n21336, n21337, n21338, n21339, n21340, n21341,
         n21342, n21343, n21344, n21345, n21346, n21347, n21348, n21349,
         n21350, n21351, n21352, n21353, n21354, n21355, n21356, n21357,
         n21358, n21359, n21360, n21361, n21362, n21363, n21364, n21365,
         n21366, n21367, n21368, n21369, n21370, n21371, n21372, n21373,
         n21374, n21375, n21376, n21377, n21378, n21379, n21380, n21381,
         n21382, n21383, n21384, n21385, n21386, n21387, n21388, n21389,
         n21390, n21391, n21392, n21393, n21394, n21395, n21396, n21397,
         n21398, n21399, n21400, n21401, n21402, n21403, n21404, n21405,
         n21406, n21407, n21408, n21409, n21410, n21411, n21412, n21413,
         n21414, n21415, n21416, n21417, n21418, n21419, n21420, n21421,
         n21422, n21423, n21424, n21425, n21426, n21427, n21428, n21429,
         n21430, n21431, n21432, n21433, n21434, n21435, n21436, n21437,
         n21438, n21439, n21440, n21441, n21442, n21443, n21444, n21445,
         n21446, n21447, n21448, n21449, n21450, n21451, n21452, n21453,
         n21454, n21455, n21456, n21457, n21458, n21459, n21460, n21461,
         n21462, n21463, n21464, n21465, n21466, n21467, n21468, n21469,
         n21470, n21471, n21472, n21473, n21474, n21475, n21476, n21477,
         n21478, n21479, n21480, n21481, n21482, n21483, n21484, n21485,
         n21486, n21487, n21488, n21489, n21490, n21491, n21492, n21493,
         n21494, n21495, n21496, n21497, n21498, n21499, n21500, n21501,
         n21502, n21503, n21504, n21505, n21506, n21507, n21508, n21509,
         n21510, n21511, n21512, n21513, n21514, n21515, n21516, n21517,
         n21518, n21519, n21520, n21521, n21522, n21523, n21524, n21525,
         n21526, n21527, n21528, n21529, n21530, n21531, n21532, n21533,
         n21534, n21535, n21536, n21537, n21538, n21539, n21540, n21541,
         n21542, n21543, n21544, n21545, n21546, n21547, n21548, n21549,
         n21550, n21551, n21552, n21553, n21554, n21555, n21556, n21557,
         n21558, n21559, n21560, n21561, n21562, n21563, n21564, n21565,
         n21566, n21567, n21568, n21569, n21570, n21571, n21572, n21573,
         n21574, n21575, n21576, n21577, n21578, n21579, n21580, n21581,
         n21582, n21583, n21584, n21585, n21586, n21587, n21588, n21589,
         n21590, n21591, n21592, n21593, n21594, n21595, n21596, n21597,
         n21598, n21599, n21600, n21601, n21602, n21603, n21604, n21605,
         n21606, n21607, n21608, n21609, n21610, n21611, n21612, n21613,
         n21614, n21615, n21616, n21617, n21618, n21619, n21620, n21621,
         n21622, n21623, n21624, n21625, n21626, n21627, n21628, n21629,
         n21630, n21631, n21632, n21633, n21634, n21635, n21636, n21637,
         n21638, n21639, n21640, n21641, n21642, n21643, n21644, n21645,
         n21646, n21647, n21648, n21649, n21650, n21651, n21652, n21653,
         n21654, n21655, n21656, n21657, n21658, n21659, n21660, n21661,
         n21662, n21663, n21664, n21665, n21666, n21667, n21668, n21669,
         n21670, n21671, n21672, n21673, n21674, n21675, n21676, n21677,
         n21678, n21679, n21680, n21681, n21682, n21683, n21684, n21685,
         n21686, n21687, n21688, n21689, n21690, n21691, n21692, n21693,
         n21694, n21695, n21696, n21697, n21698, n21699, n21700, n21701,
         n21702, n21703, n21704, n21705, n21706, n21707, n21708, n21709,
         n21710, n21711, n21712, n21713, n21714, n21715, n21716, n21717,
         n21718, n21719, n21720, n21721, n21722, n21723, n21724, n21725,
         n21726, n21727, n21728, n21729, n21730, n21731, n21732, n21733,
         n21734, n21735, n21736, n21737, n21738, n21739, n21740, n21741,
         n21742, n21743, n21744, n21745, n21746, n21747, n21748, n21749,
         n21750, n21751, n21752, n21753, n21754, n21755, n21756, n21757,
         n21758, n21759, n21760, n21761, n21762, n21763, n21764, n21765,
         n21766, n21767, n21768, n21769, n21770, n21771, n21772, n21773,
         n21774, n21775, n21776, n21777, n21778, n21779, n21780, n21781,
         n21782, n21783, n21784, n21785, n21786, n21787, n21788, n21789,
         n21790, n21791, n21792, n21793, n21794, n21795, n21796, n21797,
         n21798, n21799, n21800, n21801, n21802, n21803, n21804, n21805,
         n21806, n21807, n21808, n21809, n21810, n21811, n21812, n21813,
         n21814, n21815, n21816, n21817, n21818, n21819, n21820, n21821,
         n21822, n21823, n21824, n21825, n21826, n21827, n21828, n21829,
         n21830, n21831, n21832, n21833, n21834, n21835, n21836, n21837,
         n21838, n21839, n21840, n21841, n21842, n21843, n21844, n21845,
         n21846, n21847, n21848, n21849, n21850, n21851, n21852, n21853,
         n21854, n21855, n21856, n21857, n21858, n21859, n21860, n21861,
         n21862, n21863, n21864, n21865, n21866, n21867, n21868, n21869,
         n21870, n21871, n21872, n21873, n21874, n21875, n21876, n21877,
         n21878, n21879, n21880, n21881, n21882, n21883, n21884, n21885,
         n21886, n21887, n21888, n21889, n21890, n21891, n21892, n21893,
         n21894, n21895, n21896, n21897, n21898, n21899, n21900, n21901,
         n21902, n21903, n21904, n21905, n21906, n21907, n21908, n21909,
         n21910, n21911, n21912, n21913, n21914, n21915, n21916, n21917,
         n21918, n21919, n21920, n21921, n21922, n21923, n21924, n21925,
         n21926, n21927, n21928, n21929, n21930, n21931, n21932, n21933,
         n21934, n21935, n21936, n21937, n21938, n21939, n21940, n21941,
         n21942, n21943, n21944, n21945, n21946, n21947, n21948, n21949,
         n21950, n21951, n21952, n21953, n21954, n21955, n21956, n21957,
         n21958, n21959, n21960, n21961, n21962, n21963, n21964, n21965,
         n21966, n21967, n21968, n21969, n21970, n21971, n21972, n21973,
         n21974, n21975, n21976, n21977, n21978, n21979, n21980, n21981,
         n21982, n21983, n21984, n21985, n21986, n21987, n21988, n21989,
         n21990, n21991, n21992, n21993, n21994, n21995, n21996, n21997,
         n21998, n21999, n22000, n22001, n22002, n22003, n22004, n22005,
         n22006, n22007, n22008, n22009, n22010, n22011, n22012, n22013,
         n22014, n22015, n22016, n22017, n22018, n22019, n22020, n22021,
         n22022, n22023, n22024, n22025, n22026, n22027, n22028, n22029,
         n22030, n22031, n22032, n22033, n22034, n22035, n22036, n22037,
         n22038, n22039, n22040, n22041, n22042, n22043, n22044, n22045,
         n22046, n22047, n22048, n22049, n22050, n22051, n22052, n22053,
         n22054, n22055, n22056, n22057, n22058, n22059, n22060, n22061,
         n22062, n22063, n22064, n22065, n22066, n22067, n22068, n22069,
         n22070, n22071, n22072, n22073, n22074, n22075, n22076, n22077,
         n22078, n22079, n22080, n22081, n22082, n22083, n22084, n22085,
         n22086, n22087, n22088, n22089, n22090, n22091, n22092, n22093,
         n22094, n22095, n22096, n22097, n22098, n22099, n22100, n22101,
         n22102, n22103, n22104, n22105, n22106, n22107, n22108, n22109,
         n22110, n22111, n22112, n22113, n22114, n22115, n22116, n22117,
         n22118, n22119, n22120, n22121, n22122, n22123, n22124, n22125,
         n22126, n22127, n22128, n22129, n22130, n22131, n22132, n22133,
         n22134, n22135, n22136, n22137, n22138, n22139, n22140, n22141,
         n22142, n22143, n22144, n22145, n22146, n22147, n22148, n22149,
         n22150, n22151, n22152, n22153, n22154, n22155, n22156, n22157,
         n22158, n22159, n22160, n22161, n22162, n22163, n22164, n22165,
         n22166, n22167, n22168, n22169, n22170, n22171, n22172, n22173,
         n22174, n22175, n22176, n22177, n22178, n22179, n22180, n22181,
         n22182, n22183, n22184, n22185, n22186, n22187, n22188, n22189,
         n22190, n22191, n22192, n22193, n22194, n22195, n22196, n22197,
         n22198, n22199, n22200, n22201, n22202, n22203, n22204, n22205,
         n22206, n22207, n22208, n22209, n22210, n22211, n22212, n22213,
         n22214, n22215, n22216, n22217, n22218, n22219, n22220, n22221,
         n22222, n22223, n22224, n22225, n22226, n22227, n22228, n22229,
         n22230, n22231, n22232, n22233, n22234, n22235, n22236, n22237,
         n22238, n22239, n22240, n22241, n22242, n22243, n22244, n22245,
         n22246, n22247, n22248, n22249, n22250, n22251, n22252, n22253,
         n22254, n22255, n22256, n22257, n22258, n22259, n22260, n22261,
         n22262, n22263, n22264, n22265, n22266, n22267, n22268, n22269,
         n22270, n22271, n22272, n22273, n22274, n22275, n22276, n22277,
         n22278, n22279, n22280, n22281, n22282, n22283, n22284, n22285,
         n22286, n22287, n22288, n22289, n22290, n22291, n22292, n22293,
         n22294, n22295, n22296, n22297, n22298, n22299, n22300, n22301,
         n22302, n22303, n22304, n22305, n22306, n22307, n22308, n22309,
         n22310, n22311, n22312, n22313, n22314, n22315, n22316, n22317,
         n22318, n22319, n22320, n22321, n22322, n22323, n22324, n22325,
         n22326, n22327, n22328, n22329, n22330, n22331, n22332, n22333,
         n22334, n22335, n22336, n22337, n22338, n22339, n22340, n22341,
         n22342, n22343, n22344, n22345, n22346, n22347, n22348, n22349,
         n22350, n22351, n22352, n22353, n22354, n22355, n22356, n22357,
         n22358, n22359, n22360, n22361, n22362, n22363, n22364, n22365,
         n22366, n22367, n22368, n22369, n22370, n22371, n22372, n22373,
         n22374, n22375, n22376, n22377, n22378, n22379, n22380, n22381,
         n22382, n22383, n22384, n22385, n22386, n22387, n22388, n22389,
         n22390, n22391, n22392, n22393, n22394, n22395, n22396, n22397,
         n22398, n22399, n22400, n22401, n22402, n22403, n22404, n22405,
         n22406, n22407, n22408, n22409, n22410, n22411, n22412, n22413,
         n22414, n22415, n22416, n22417, n22418, n22419, n22420, n22421,
         n22422, n22423, n22424, n22425, n22426, n22427, n22428, n22429,
         n22430, n22431, n22432, n22433, n22434, n22435, n22436, n22437,
         n22438, n22439, n22440, n22441, n22442, n22443, n22444, n22445,
         n22446, n22447, n22448, n22449, n22450, n22451, n22452, n22453,
         n22454, n22455, n22456, n22457, n22458, n22459, n22460, n22461,
         n22462, n22463, n22464, n22465, n22466, n22467, n22468, n22469,
         n22470, n22471, n22472, n22473, n22474, n22475, n22476, n22477,
         n22478, n22479, n22480, n22481, n22482, n22483, n22484, n22485,
         n22486, n22487, n22488, n22489, n22490, n22491, n22492, n22493,
         n22494, n22495, n22496, n22497, n22498, n22499, n22500, n22501,
         n22502, n22503, n22504, n22505, n22506, n22507, n22508, n22509,
         n22510, n22511, n22512, n22513, n22514, n22515, n22516, n22517,
         n22518, n22519, n22520, n22521, n22522, n22523, n22524, n22525,
         n22526, n22527, n22528, n22529, n22530, n22531, n22532, n22533,
         n22534, n22535, n22536, n22537, n22538, n22539, n22540, n22541,
         n22542, n22543, n22544, n22545, n22546, n22547, n22548, n22549,
         n22550, n22551, n22552, n22553, n22554, n22555, n22556, n22557,
         n22558, n22559, n22560, n22561, n22562, n22563, n22564, n22565,
         n22566, n22567, n22568, n22569, n22570, n22571, n22572, n22573,
         n22574, n22575, n22576, n22577, n22578, n22579, n22580, n22581,
         n22582, n22583, n22584, n22585, n22586, n22587, n22588, n22589,
         n22590, n22591, n22592, n22593, n22594, n22595, n22596, n22597,
         n22598, n22599, n22600, n22601, n22602, n22603, n22604, n22605,
         n22606, n22607, n22608, n22609, n22610, n22611, n22612, n22613,
         n22614, n22615, n22616, n22617, n22618, n22619, n22620, n22621,
         n22622, n22623, n22624, n22625, n22626, n22627, n22628, n22629,
         n22630, n22631, n22632, n22633, n22634, n22635, n22636, n22637,
         n22638, n22639, n22640, n22641, n22642, n22643, n22644, n22645,
         n22646, n22647, n22648, n22649, n22650, n22651, n22652, n22653,
         n22654, n22655, n22656, n22657, n22658, n22659, n22660, n22661,
         n22662, n22663, n22664, n22665, n22666, n22667, n22668, n22669,
         n22670, n22671, n22672, n22673, n22674, n22675, n22676, n22677,
         n22678, n22679, n22680, n22681, n22682, n22683, n22684, n22685,
         n22686, n22687, n22688, n22689, n22690, n22691, n22692, n22693,
         n22694, n22695, n22696, n22697, n22698, n22699, n22700, n22701,
         n22702, n22703, n22704, n22705, n22706, n22707, n22708, n22709,
         n22710, n22711, n22712, n22713, n22714, n22715, n22716, n22717,
         n22718, n22719, n22720, n22721, n22722, n22723, n22724, n22725,
         n22726, n22727, n22728, n22729, n22730, n22731, n22732, n22733,
         n22734, n22735, n22736, n22737, n22738, n22739, n22740, n22741,
         n22742, n22743, n22744, n22745, n22746, n22747, n22748, n22749,
         n22750, n22751, n22752, n22753, n22754, n22755, n22756, n22757,
         n22758, n22759, n22760, n22761, n22762, n22763, n22764, n22765,
         n22766, n22767, n22768, n22769, n22770, n22771, n22772, n22773,
         n22774, n22775, n22776, n22777, n22778, n22779, n22780, n22781,
         n22782, n22783, n22784, n22785, n22786, n22787, n22788, n22789,
         n22790, n22791, n22792, n22793, n22794, n22795, n22796, n22797,
         n22798, n22799, n22800, n22801, n22802, n22803, n22804, n22805,
         n22806, n22807, n22808, n22809, n22810, n22811, n22812, n22813,
         n22814, n22815, n22816, n22817, n22818, n22819, n22820, n22821,
         n22822, n22823, n22824, n22825, n22826, n22827, n22828, n22829,
         n22830, n22831, n22832, n22833, n22834, n22835, n22836, n22837,
         n22838, n22839, n22840, n22841, n22842, n22843, n22844, n22845,
         n22846, n22847, n22848, n22849, n22850, n22851, n22852, n22853,
         n22854, n22855, n22856, n22857, n22858, n22859, n22860, n22861,
         n22862, n22863, n22864, n22865, n22866, n22867, n22868, n22869,
         n22870, n22871, n22872, n22873, n22874, n22875, n22876, n22877,
         n22878, n22879, n22880, n22881, n22882, n22883, n22884, n22885,
         n22886, n22887, n22888, n22889, n22890, n22891, n22892, n22893,
         n22894, n22895, n22896, n22897, n22898, n22899, n22900, n22901,
         n22902, n22903, n22904, n22905, n22906, n22907, n22908, n22909,
         n22910, n22911, n22912, n22913, n22914, n22915, n22916, n22917,
         n22918, n22919, n22920, n22921, n22922, n22923, n22924, n22925,
         n22926, n22927, n22928, n22929, n22930, n22931, n22932, n22933,
         n22934, n22935, n22936, n22937, n22938, n22939, n22940, n22941,
         n22942, n22943, n22944, n22945, n22946, n22947, n22948, n22949,
         n22950, n22951, n22952, n22953, n22954, n22955, n22956, n22957,
         n22958, n22959, n22960, n22961, n22962, n22963, n22964, n22965,
         n22966, n22967, n22968, n22969, n22970, n22971, n22972, n22973,
         n22974, n22975, n22976, n22977, n22978, n22979, n22980, n22981,
         n22982, n22983, n22984, n22985, n22986, n22987, n22988, n22989,
         n22990, n22991, n22992, n22993, n22994, n22995, n22996, n22997,
         n22998, n22999, n23000, n23001, n23002, n23003, n23004, n23005,
         n23006, n23007, n23008, n23009, n23010, n23011, n23012, n23013,
         n23014, n23015, n23016, n23017, n23018, n23019, n23020, n23021,
         n23022, n23023, n23024, n23025, n23026, n23027, n23028, n23029,
         n23030, n23031, n23032, n23033, n23034, n23035, n23036, n23037,
         n23038, n23039, n23040, n23041, n23042, n23043, n23044, n23045,
         n23046, n23047, n23048, n23049, n23050, n23051, n23052, n23053,
         n23054, n23055, n23056, n23057, n23058, n23059, n23060, n23061,
         n23062, n23063, n23064, n23065, n23066, n23067, n23068, n23069,
         n23070, n23071, n23072, n23073, n23074, n23075, n23076, n23077,
         n23078, n23079, n23080, n23081, n23082, n23083, n23084, n23085,
         n23086, n23087, n23088, n23089, n23090, n23091, n23092, n23093,
         n23094, n23095, n23096, n23097, n23098, n23099, n23100, n23101,
         n23102, n23103, n23104, n23105, n23106, n23107, n23108, n23109,
         n23110, n23111, n23112, n23113, n23114, n23115, n23116, n23117,
         n23118, n23119, n23120, n23121, n23122, n23123, n23124, n23125,
         n23126, n23127, n23128, n23129, n23130, n23131, n23132, n23133,
         n23134, n23135, n23136, n23137, n23138, n23139, n23140, n23141,
         n23142, n23143, n23144, n23145, n23146, n23147, n23148, n23149,
         n23150, n23151, n23152, n23153, n23154, n23155, n23156, n23157,
         n23158, n23159, n23160, n23161, n23162, n23163, n23164, n23165,
         n23166, n23167, n23168, n23169, n23170, n23171, n23172, n23173,
         n23174, n23175, n23176, n23177, n23178, n23179, n23180, n23181,
         n23182, n23183, n23184, n23185, n23186, n23187, n23188, n23189,
         n23190, n23191, n23192, n23193, n23194, n23195, n23196, n23197,
         n23198, n23199, n23200, n23201, n23202, n23203, n23204, n23205,
         n23206, n23207, n23208, n23209, n23210, n23211, n23212, n23213,
         n23214, n23215, n23216, n23217, n23218, n23219, n23220, n23221,
         n23222, n23223, n23224, n23225, n23226, n23227, n23228, n23229,
         n23230, n23231, n23232, n23233, n23234, n23235, n23236, n23237,
         n23238, n23239, n23240, n23241, n23242, n23243, n23244, n23245,
         n23246, n23247, n23248, n23249, n23250, n23251, n23252, n23253,
         n23254, n23255, n23256, n23257, n23258, n23259, n23260, n23261,
         n23262, n23263, n23264, n23265, n23266, n23267, n23268, n23269,
         n23270, n23271, n23272, n23273, n23274, n23275, n23276, n23277,
         n23278, n23279, n23280, n23281, n23282, n23283, n23284, n23285,
         n23286, n23287, n23288, n23289, n23290, n23291, n23292, n23293,
         n23294, n23295, n23296, n23297, n23298, n23299, n23300, n23301,
         n23302, n23303, n23304, n23305, n23306, n23307, n23308, n23309,
         n23310, n23311, n23312, n23313, n23314, n23315, n23316, n23317,
         n23318, n23319, n23320, n23321, n23322, n23323, n23324, n23325,
         n23326, n23327, n23328, n23329, n23330, n23331, n23332, n23333,
         n23334, n23335, n23336, n23337, n23338, n23339, n23340, n23341,
         n23342, n23343, n23344, n23345, n23346, n23347, n23348, n23349,
         n23350, n23351, n23352, n23353, n23354, n23355, n23356, n23357,
         n23358, n23359, n23360, n23361, n23362, n23363, n23364, n23365,
         n23366, n23367, n23368, n23369, n23370, n23371, n23372, n23373,
         n23374, n23375, n23376, n23377, n23378, n23379, n23380, n23381,
         n23382, n23383, n23384, n23385, n23386, n23387, n23388, n23389,
         n23390, n23391, n23392, n23393, n23394, n23395, n23396, n23397,
         n23398, n23399, n23400, n23401, n23402, n23403, n23404, n23405,
         n23406, n23407, n23408, n23409, n23410, n23411, n23412, n23413,
         n23414, n23415, n23416, n23417, n23418, n23419, n23420, n23421,
         n23422, n23423, n23424, n23425, n23426, n23427, n23428, n23429,
         n23430, n23431, n23432, n23433, n23434, n23435, n23436, n23437,
         n23438, n23439, n23440, n23441, n23442, n23443, n23444, n23445,
         n23446, n23447, n23448, n23449, n23450, n23451, n23452, n23453,
         n23454, n23455, n23456, n23457, n23458, n23459, n23460, n23461,
         n23462, n23463, n23464, n23465, n23466, n23467, n23468, n23469,
         n23470, n23471, n23472, n23473, n23474, n23475, n23476, n23477,
         n23478, n23479, n23480, n23481, n23482, n23483, n23484, n23485,
         n23486, n23487, n23488, n23489, n23490, n23491, n23492, n23493,
         n23494, n23495, n23496, n23497, n23498, n23499, n23500, n23501,
         n23502, n23503, n23504, n23505, n23506, n23507, n23508, n23509,
         n23510, n23511, n23512, n23513, n23514, n23515, n23516, n23517,
         n23518, n23519, n23520, n23521, n23522, n23523, n23524, n23525,
         n23526, n23527, n23528, n23529, n23530, n23531, n23532, n23533,
         n23534, n23535, n23536, n23537, n23538, n23539, n23540, n23541,
         n23542, n23543, n23544, n23545, n23546, n23547, n23548, n23549,
         n23550, n23551, n23552, n23553, n23554, n23555, n23556, n23557,
         n23558, n23559, n23560, n23561, n23562, n23563, n23564, n23565,
         n23566, n23567, n23568, n23569, n23570, n23571, n23572, n23573,
         n23574, n23575, n23576, n23577, n23578, n23579, n23580, n23581,
         n23582, n23583, n23584, n23585, n23586, n23587, n23588, n23589,
         n23590, n23591, n23592, n23593, n23594, n23595, n23596, n23597,
         n23598, n23599, n23600, n23601, n23602, n23603, n23604, n23605,
         n23606, n23607, n23608, n23609, n23610, n23611, n23612, n23613,
         n23614, n23615, n23616, n23617, n23618, n23619, n23620, n23621,
         n23622, n23623, n23624, n23625, n23626, n23627, n23628, n23629,
         n23630, n23631, n23632, n23633, n23634, n23635, n23636, n23637,
         n23638, n23639, n23640, n23641, n23642, n23643, n23644, n23645,
         n23646, n23647, n23648, n23649, n23650, n23651, n23652, n23653,
         n23654, n23655, n23656, n23657, n23658, n23659, n23660, n23661,
         n23662, n23663, n23664, n23665, n23666, n23667, n23668, n23669,
         n23670, n23671, n23672, n23673, n23674, n23675, n23676, n23677,
         n23678, n23679, n23680, n23681, n23682, n23683, n23684, n23685,
         n23686, n23687, n23688, n23689, n23690, n23691, n23692, n23693,
         n23694, n23695, n23696, n23697, n23698, n23699, n23700, n23701,
         n23702, n23703, n23704, n23705, n23706, n23707, n23708, n23709,
         n23710, n23711, n23712, n23713, n23714, n23715, n23716, n23717,
         n23718, n23719, n23720, n23721, n23722, n23723, n23724, n23725,
         n23726, n23727, n23728, n23729, n23730, n23731, n23732, n23733,
         n23734, n23735, n23736, n23737, n23738, n23739, n23740, n23741,
         n23742, n23743, n23744, n23745, n23746, n23747, n23748, n23749,
         n23750, n23751, n23752, n23753, n23754, n23755, n23756, n23757,
         n23758, n23759, n23760, n23761, n23762, n23763, n23764, n23765,
         n23766, n23767, n23768, n23769, n23770, n23771, n23772, n23773,
         n23774, n23775, n23776, n23777, n23778, n23779, n23780, n23781,
         n23782, n23783, n23784, n23785, n23786, n23787, n23788, n23789,
         n23790, n23791, n23792, n23793, n23794, n23795, n23796, n23797,
         n23798, n23799, n23800, n23801, n23802, n23803, n23804, n23805,
         n23806, n23807, n23808, n23809, n23810, n23811, n23812, n23813,
         n23814, n23815, n23816, n23817, n23818, n23819, n23820, n23821,
         n23822, n23823, n23824, n23825, n23826, n23827, n23828, n23829,
         n23830, n23831, n23832, n23833, n23834, n23835, n23836, n23837,
         n23838, n23839, n23840, n23841, n23842, n23843, n23844, n23845,
         n23846, n23847, n23848, n23849, n23850, n23851, n23852, n23853,
         n23854, n23855, n23856, n23857, n23858, n23859, n23860, n23861,
         n23862, n23863, n23864, n23865, n23866, n23867, n23868, n23869,
         n23870, n23871, n23872, n23873, n23874, n23875, n23876, n23877,
         n23878, n23879, n23880, n23881, n23882, n23883, n23884, n23885,
         n23886, n23887, n23888, n23889, n23890, n23891, n23892, n23893,
         n23894, n23895, n23896, n23897, n23898, n23899, n23900, n23901,
         n23902, n23903, n23904, n23905, n23906, n23907, n23908, n23909,
         n23910, n23911, n23912, n23913, n23914, n23915, n23916, n23917,
         n23918, n23919, n23920, n23921, n23922, n23923, n23924, n23925,
         n23926, n23927, n23928, n23929, n23930, n23931, n23932, n23933,
         n23934, n23935, n23936, n23937, n23938, n23939, n23940, n23941,
         n23942, n23943, n23944, n23945, n23946, n23947, n23948, n23949,
         n23950, n23951, n23952, n23953, n23954, n23955, n23956, n23957,
         n23958, n23959, n23960, n23961, n23962, n23963, n23964, n23965,
         n23966, n23967, n23968, n23969, n23970, n23971, n23972, n23973,
         n23974, n23975, n23976, n23977, n23978, n23979, n23980, n23981,
         n23982, n23983, n23984, n23985, n23986, n23987, n23988, n23989,
         n23990, n23991, n23992, n23993, n23994, n23995, n23996, n23997,
         n23998, n23999, n24000, n24001, n24002, n24003, n24004, n24005,
         n24006, n24007, n24008, n24009, n24010, n24011, n24012, n24013,
         n24014, n24015, n24016, n24017, n24018, n24019, n24020, n24021,
         n24022, n24023, n24024, n24025, n24026, n24027, n24028, n24029,
         n24030, n24031, n24032, n24033, n24034, n24035, n24036, n24037,
         n24038, n24039, n24040, n24041, n24042, n24043, n24044, n24045,
         n24046, n24047, n24048, n24049, n24050, n24051, n24052, n24053,
         n24054, n24055, n24056, n24057, n24058, n24059, n24060, n24061,
         n24062, n24063, n24064, n24065, n24066, n24067, n24068, n24069,
         n24070, n24071, n24072, n24073, n24074, n24075, n24076, n24077,
         n24078, n24079, n24080, n24081, n24082, n24083, n24084, n24085,
         n24086, n24087, n24088, n24089, n24090, n24091, n24092, n24093,
         n24094, n24095, n24096, n24097, n24098, n24099, n24100, n24101,
         n24102, n24103, n24104, n24105, n24106, n24107, n24108, n24109,
         n24110, n24111, n24112, n24113, n24114, n24115, n24116, n24117,
         n24118, n24119, n24120, n24121, n24122, n24123, n24124, n24125,
         n24126, n24127, n24128, n24129, n24130, n24131, n24132, n24133,
         n24134, n24135, n24136, n24137, n24138, n24139, n24140, n24141,
         n24142, n24143, n24144, n24145, n24146, n24147, n24148, n24149,
         n24150, n24151, n24152, n24153, n24154, n24155, n24156, n24157,
         n24158, n24159, n24160, n24161, n24162, n24163, n24164, n24165,
         n24166, n24167, n24168, n24169, n24170, n24171, n24172, n24173,
         n24174, n24175, n24176, n24177, n24178, n24179, n24180, n24181,
         n24182, n24183, n24184, n24185, n24186, n24187, n24188, n24189,
         n24190, n24191, n24192, n24193, n24194, n24195, n24196, n24197,
         n24198, n24199, n24200, n24201, n24202, n24203, n24204, n24205,
         n24206, n24207, n24208, n24209, n24210, n24211, n24212, n24213,
         n24214, n24215, n24216, n24217, n24218, n24219, n24220, n24221,
         n24222, n24223, n24224, n24225, n24226, n24227, n24228, n24229,
         n24230, n24231, n24232, n24233, n24234, n24235, n24236, n24237,
         n24238, n24239, n24240, n24241, n24242, n24243, n24244, n24245,
         n24246, n24247, n24248, n24249, n24250, n24251, n24252, n24253,
         n24254, n24255, n24256, n24257, n24258, n24259, n24260, n24261,
         n24262, n24263, n24264, n24265, n24266, n24267, n24268, n24269,
         n24270, n24271, n24272, n24273, n24274, n24275, n24276, n24277,
         n24278, n24279, n24280, n24281, n24282, n24283, n24284, n24285,
         n24286, n24287, n24288, n24289, n24290, n24291, n24292, n24293,
         n24294, n24295, n24296, n24297, n24298, n24299, n24300, n24301,
         n24302, n24303, n24304, n24305, n24306, n24307, n24308, n24309,
         n24310, n24311, n24312, n24313, n24314, n24315, n24316, n24317,
         n24318, n24319, n24320, n24321, n24322, n24323, n24324, n24325,
         n24326, n24327, n24328, n24329, n24330, n24331, n24332, n24333,
         n24334, n24335, n24336, n24337, n24338, n24339, n24340, n24341,
         n24342, n24343, n24344, n24345, n24346, n24347, n24348, n24349,
         n24350, n24351, n24352, n24353, n24354, n24355, n24356, n24357,
         n24358, n24359, n24360, n24361, n24362, n24363, n24364, n24365,
         n24366, n24367, n24368, n24369, n24370, n24371, n24372, n24373,
         n24374, n24375, n24376, n24377, n24378, n24379, n24380, n24381,
         n24382, n24383, n24384, n24385, n24386, n24387, n24388, n24389,
         n24390, n24391, n24392, n24393, n24394, n24395, n24396, n24397,
         n24398, n24399, n24400, n24401, n24402, n24403, n24404, n24405,
         n24406, n24407, n24408, n24409, n24410, n24411, n24412, n24413,
         n24414, n24415, n24416, n24417, n24418, n24419, n24420, n24421,
         n24422, n24423, n24424, n24425, n24426, n24427, n24428, n24429,
         n24430, n24431, n24432, n24433, n24434, n24435, n24436, n24437,
         n24438, n24439, n24440, n24441, n24442, n24443, n24444, n24445,
         n24446, n24447, n24448, n24449, n24450, n24451, n24452, n24453,
         n24454, n24455, n24456, n24457, n24458, n24459, n24460, n24461,
         n24462, n24463, n24464, n24465, n24466, n24467, n24468, n24469,
         n24470, n24471, n24472, n24473, n24474, n24475, n24476, n24477,
         n24478, n24479, n24480, n24481, n24482, n24483, n24484, n24485,
         n24486, n24487, n24488, n24489, n24490, n24491, n24492, n24493,
         n24494, n24495, n24496, n24497, n24498, n24499, n24500, n24501,
         n24502, n24503, n24504, n24505, n24506, n24507, n24508, n24509,
         n24510, n24511, n24512, n24513, n24514, n24515, n24516, n24517,
         n24518, n24519, n24520, n24521, n24522, n24523, n24524, n24525,
         n24526, n24527, n24528, n24529, n24530, n24531, n24532, n24533,
         n24534, n24535, n24536, n24537, n24538, n24539, n24540, n24541,
         n24542, n24543, n24544, n24545, n24546, n24547, n24548, n24549,
         n24550, n24551, n24552, n24553, n24554, n24555, n24556, n24557,
         n24558, n24559, n24560, n24561, n24562, n24563, n24564, n24565,
         n24566, n24567, n24568, n24569, n24570, n24571, n24572, n24573,
         n24574, n24575, n24576, n24577, n24578, n24579, n24580, n24581,
         n24582, n24583, n24584, n24585, n24586, n24587, n24588, n24589,
         n24590, n24591, n24592, n24593, n24594, n24595, n24596, n24597,
         n24598, n24599, n24600, n24601, n24602, n24603, n24604, n24605,
         n24606, n24607, n24608, n24609, n24610, n24611, n24612, n24613,
         n24614, n24615, n24616, n24617, n24618, n24619, n24620, n24621,
         n24622, n24623, n24624, n24625, n24626, n24627, n24628, n24629,
         n24630, n24631, n24632, n24633, n24634, n24635, n24636, n24637,
         n24638, n24639, n24640, n24641, n24642, n24643, n24644, n24645,
         n24646, n24647, n24648, n24649, n24650, n24651, n24652, n24653,
         n24654, n24655, n24656, n24657, n24658, n24659, n24660, n24661,
         n24662, n24663, n24664, n24665, n24666, n24667, n24668, n24669,
         n24670, n24671, n24672, n24673, n24674, n24675, n24676, n24677,
         n24678, n24679, n24680, n24681, n24682, n24683, n24684, n24685,
         n24686, n24687, n24688, n24689, n24690, n24691, n24692, n24693,
         n24694, n24695, n24696, n24697, n24698, n24699, n24700, n24701,
         n24702, n24703, n24704, n24705, n24706, n24707, n24708, n24709,
         n24710, n24711, n24712, n24713, n24714, n24715, n24716, n24717,
         n24718, n24719, n24720, n24721, n24722, n24723, n24724, n24725,
         n24726, n24727, n24728, n24729, n24730, n24731, n24732, n24733,
         n24734, n24735, n24736, n24737, n24738, n24739, n24740, n24741,
         n24742, n24743, n24744, n24745, n24746, n24747, n24748, n24749,
         n24750, n24751, n24752, n24753, n24754, n24755, n24756, n24757,
         n24758, n24759, n24760, n24761, n24762, n24763, n24764, n24765,
         n24766, n24767, n24768, n24769, n24770, n24771, n24772, n24773,
         n24774, n24775, n24776, n24777, n24778, n24779, n24780, n24781,
         n24782, n24783, n24784, n24785, n24786, n24787, n24788, n24789,
         n24790, n24791, n24792, n24793, n24794, n24795, n24796, n24797,
         n24798, n24799, n24800, n24801, n24802, n24803, n24804, n24805,
         n24806, n24807, n24808, n24809, n24810, n24811, n24812, n24813,
         n24814, n24815, n24816, n24817, n24818, n24819, n24820, n24821,
         n24822, n24823, n24824, n24825, n24826, n24827, n24828, n24829,
         n24830, n24831, n24832, n24833, n24834, n24835, n24836, n24837,
         n24838, n24839, n24840, n24841, n24842, n24843, n24844, n24845,
         n24846, n24847, n24848, n24849, n24850, n24851, n24852, n24853,
         n24854, n24855, n24856, n24857, n24858, n24859, n24860, n24861,
         n24862, n24863, n24864, n24865, n24866, n24867, n24868, n24869,
         n24870, n24871, n24872, n24873, n24874, n24875, n24876, n24877,
         n24878, n24879, n24880, n24881, n24882, n24883, n24884, n24885,
         n24886, n24887, n24888, n24889, n24890, n24891, n24892, n24893,
         n24894, n24895, n24896, n24897, n24898, n24899, n24900, n24901,
         n24902, n24903, n24904, n24905, n24906, n24907, n24908, n24909,
         n24910, n24911, n24912, n24913, n24914, n24915, n24916, n24917,
         n24918, n24919, n24920, n24921, n24922, n24923, n24924, n24925,
         n24926, n24927, n24928, n24929, n24930, n24931, n24932, n24933,
         n24934, n24935, n24936, n24937, n24938, n24939, n24940, n24941,
         n24942, n24943, n24944, n24945, n24946, n24947, n24948, n24949,
         n24950, n24951, n24952, n24953, n24954, n24955, n24956, n24957,
         n24958, n24959, n24960, n24961, n24962, n24963, n24964, n24965,
         n24966, n24967, n24968, n24969, n24970, n24971, n24972, n24973,
         n24974, n24975, n24976, n24977, n24978, n24979, n24980, n24981,
         n24982, n24983, n24984, n24985, n24986, n24987, n24988, n24989,
         n24990, n24991, n24992, n24993, n24994, n24995, n24996, n24997,
         n24998, n24999, n25000, n25001, n25002, n25003, n25004, n25005,
         n25006, n25007, n25008, n25009, n25010, n25011, n25012, n25013,
         n25014, n25015, n25016, n25017, n25018, n25019, n25020, n25021,
         n25022, n25023, n25024, n25025, n25026, n25027, n25028, n25029,
         n25030, n25031, n25032, n25033, n25034, n25035, n25036, n25037,
         n25038, n25039, n25040, n25041, n25042, n25043, n25044, n25045,
         n25046, n25047, n25048, n25049, n25050, n25051, n25052, n25053,
         n25054, n25055, n25056, n25057, n25058, n25059, n25060, n25061,
         n25062, n25063, n25064, n25065, n25066, n25067, n25068, n25069,
         n25070, n25071, n25072, n25073, n25074, n25075, n25076, n25077,
         n25078, n25079, n25080, n25081, n25082, n25083, n25084, n25085,
         n25086, n25087, n25088, n25089, n25090, n25091, n25092, n25093,
         n25094, n25095, n25096, n25097, n25098, n25099, n25100, n25101,
         n25102, n25103, n25104, n25105, n25106, n25107, n25108, n25109,
         n25110, n25111, n25112, n25113, n25114, n25115, n25116, n25117,
         n25118, n25119, n25120, n25121, n25122, n25123, n25124, n25125,
         n25126, n25127, n25128, n25129, n25130, n25131, n25132, n25133,
         n25134, n25135, n25136, n25137, n25138, n25139, n25140, n25141,
         n25142, n25143, n25144, n25145, n25146, n25147, n25148, n25149,
         n25150, n25151, n25152, n25153, n25154, n25155, n25156, n25157,
         n25158, n25159, n25160, n25161, n25162, n25163, n25164, n25165,
         n25166, n25167, n25168, n25169, n25170, n25171, n25172, n25173,
         n25174, n25175, n25176, n25177, n25178, n25179, n25180, n25181,
         n25182, n25183, n25184, n25185, n25186, n25187, n25188, n25189,
         n25190, n25191, n25192, n25193, n25194, n25195, n25196, n25197,
         n25198, n25199, n25200, n25201, n25202, n25203, n25204, n25205,
         n25206, n25207, n25208, n25209, n25210, n25211, n25212, n25213,
         n25214, n25215, n25216, n25217, n25218, n25219, n25220, n25221,
         n25222, n25223, n25224, n25225, n25226, n25227, n25228, n25229,
         n25230, n25231, n25232, n25233, n25234, n25235, n25236, n25237,
         n25238, n25239, n25240, n25241, n25242, n25243, n25244, n25245,
         n25246, n25247, n25248, n25249, n25250, n25251, n25252, n25253,
         n25254, n25255, n25256, n25257, n25258, n25259, n25260, n25261,
         n25262, n25263, n25264, n25265, n25266, n25267, n25268, n25269,
         n25270, n25271, n25272, n25273, n25274, n25275, n25276, n25277,
         n25278, n25279, n25280, n25281, n25282, n25283, n25284, n25285,
         n25286, n25287, n25288, n25289, n25290, n25291, n25292, n25293,
         n25294, n25295, n25296, n25297, n25298, n25299, n25300, n25301,
         n25302, n25303, n25304, n25305, n25306, n25307, n25308, n25309,
         n25310, n25311, n25312, n25313, n25314, n25315, n25316, n25317,
         n25318, n25319, n25320, n25321, n25322, n25323, n25324, n25325,
         n25326, n25327, n25328, n25329, n25330, n25331, n25332, n25333,
         n25334, n25335, n25336, n25337, n25338, n25339, n25340, n25341,
         n25342, n25343, n25344, n25345, n25346, n25347, n25348, n25349,
         n25350, n25351, n25352, n25353, n25354, n25355, n25356, n25357,
         n25358, n25359, n25360, n25361, n25362, n25363, n25364, n25365,
         n25366, n25367, n25368, n25369, n25370, n25371, n25372, n25373,
         n25374, n25375, n25376, n25377, n25378, n25379, n25380, n25381,
         n25382, n25383, n25384, n25385, n25386, n25387, n25388, n25389,
         n25390, n25391, n25392, n25393, n25394, n25395, n25396, n25397,
         n25398, n25399, n25400, n25401, n25402, n25403, n25404, n25405,
         n25406, n25407, n25408, n25409, n25410, n25411, n25412, n25413,
         n25414, n25415, n25416, n25417, n25418, n25419, n25420, n25421,
         n25422, n25423, n25424, n25425, n25426, n25427, n25428, n25429,
         n25430, n25431, n25432, n25433, n25434, n25435, n25436, n25437,
         n25438, n25439, n25440, n25441, n25442, n25443, n25444, n25445,
         n25446, n25447, n25448, n25449, n25450, n25451, n25452, n25453,
         n25454, n25455, n25456, n25457, n25458, n25459, n25460, n25461,
         n25462, n25463, n25464, n25465, n25466, n25467, n25468, n25469,
         n25470, n25471, n25472, n25473, n25474, n25475, n25476, n25477,
         n25478, n25479, n25480, n25481, n25482, n25483, n25484, n25485,
         n25486, n25487, n25488, n25489, n25490, n25491, n25492, n25493,
         n25494, n25495, n25496, n25497, n25498, n25499, n25500, n25501,
         n25502, n25503, n25504, n25505, n25506, n25507, n25508, n25509,
         n25510, n25511, n25512, n25513, n25514, n25515, n25516, n25517,
         n25518, n25519, n25520, n25521, n25522, n25523, n25524, n25525,
         n25526, n25527, n25528, n25529, n25530, n25531, n25532, n25533,
         n25534, n25535, n25536, n25537, n25538, n25539, n25540, n25541,
         n25542, n25543, n25544, n25545, n25546, n25547, n25548, n25549,
         n25550, n25551, n25552, n25553, n25554, n25555, n25556, n25557,
         n25558, n25559, n25560, n25561, n25562, n25563, n25564, n25565,
         n25566, n25567, n25568, n25569, n25570, n25571, n25572, n25573,
         n25574, n25575, n25576, n25577, n25578, n25579, n25580, n25581,
         n25582, n25583, n25584, n25585, n25586, n25587, n25588, n25589,
         n255901, n25591, n25592, n25593, n25594, n25595, n25596, n25597,
         n25598, n25599, n256001, n25601, n25602, n25603, n25604, n25605,
         n25606, n25607, n25608, n25609, n256101, n25611, n25612, n25613,
         n25614, n25615, n25616, n25617, n25618, n25619, n256201, n25621,
         n25622, n25623, n25624, n25625, n25626, n25627, n25628, n25629,
         n256301, n25631, n25632, n25633, n25634, n25635, n25636, n25637,
         n25638, n25639, n256401, n25641, n25642, n25643, n25644, n25645,
         n25646, n25647, n25648, n25649, n256501, n25651, n25652, n25653,
         n25654, n25655, n25656, n25657, n25658, n25659, n256601, n25661,
         n25662, n25663, n25664, n25665, n25666, n25667, n25668, n25669,
         n256701, n25671, n25672, n25673, n25674, n25675, n25676, n25677,
         n25678, n25679, n256801, n25681, n25682, n25683, n25684, n25685,
         n25686, n25687, n25688, n25689, n256901, n25691, n25692, n25693,
         n25694, n25695, n25696, n25697, n25698, n25699, n257001, n25701,
         n25702, n25703, n25704, n25705, n25706, n25707, n25708, n25709,
         n257101, n25711, n25712, n25713, n25714, n25715, n25716, n25717,
         n25718, n25719, n257201, n25721, n25722, n25723, n25724, n25725,
         n25726, n25727, n25728, n25729, n257301, n25731, n25732, n25733,
         n25734, n25735, n25736, n25737, n25738, n25739, n257401, n25741,
         n25742, n25743, n25744, n25745, n25746, n25747, n25748, n25749,
         n25750, n25751, n25752, n25753, n25754, n25755, n25756, n25757,
         n25758, n25759, n25760, n25761, n25762, n25763, n25764, n25765,
         n25766, n25767, n25768, n25769, n25770, n25771, n25772, n25773,
         n25774, n25775, n25776, n25777, n25778, n25779, n25780, n25781,
         n25782, n25783, n25784, n25785, n25786, n25787, n25788, n25789,
         n25790, n25791, n25792, n25793, n25794, n25795, n25796, n25797,
         n25798, n25799, n25800, n25801, n25802, n25803, n25804, n25805,
         n25806, n25807, n25808, n25809, n25810, n25811, n25812, n25813,
         n25814, n25815, n25816, n25817, n25818, n25819, n25820, n25821,
         n25822, n25823, n25824, n25825, n25826, n25827, n25828, n25829,
         n25830, n25831, n25832, n25833, n25834, n25835, n25836, n25837,
         n25838, n25839, n25840, n25841, n25842, n25843, n25844, n25845,
         n25846, n25847, n25848, n25849, n25850, n25851, n25852, n25853,
         n25854, n25855, n25856, n25857, n25858, n25859, n25860, n25861,
         n25862, n25863, n25864, n25865, n25866, n25867, n25868, n25869,
         n25870, n25871, n25872, n25873, n25874, n25875, n25876, n25877,
         n25878, n25879, n25880, n25881, n25882, n25883, n25884, n25885,
         n25886, n25887, n25888, n25889, n25890, n25891, n25892, n25893,
         n25894, n25895, n25896, n25897, n25898, n25899, n25900, n25901,
         n25902, n25903, n25904, n25905, n25906, n25907, n25908, n25909,
         n25910, n25911, n25912, n25913, n25914, n25915, n25916, n25917,
         n25918, n25919, n259201, n25921, n25922, n25923, n25924, n25925,
         n25926, n25927, n25928, n25929, n259301, n25931, n25932, n25933,
         n25934, n25935, n25936, n25937, n25938, n25939, n259401, n25941,
         n25942, n25943, n25944, n25945, n25946, n25947, n25948, n25949,
         n259501, n25951, n25952, n25953, n25954, n25955, n25956, n25957,
         n25958, n25959, n259601, n25961, n25962, n25963, n25964, n25965,
         n25966, n25967, n25968, n25969, n259701, n25971, n25972, n25973,
         n25974, n25975, n25976, n25977, n25978, n25979, n259801, n25981,
         n25982, n25983, n25984, n25985, n25986, n25987, n25988, n25989,
         n259901, n25991, n25992, n25993, n25994, n25995, n25996, n25997,
         n25998, n25999, n260001, n26001, n26002, n26003, n26004, n26005,
         n26006, n26007, n26008, n26009, n260101, n26011, n26012, n26013,
         n26014, n26015, n26016, n26017, n26018, n26019, n260201, n26021,
         n26022, n26023, n26024, n26025, n26026, n26027, n26028, n26029,
         n260301, n26031, n26032, n26033, n26034, n26035, n26036, n26037,
         n26038, n26039, n260401, n26041, n26042, n26043, n26044, n26045,
         n26046, n26047, n26048, n26049, n260501, n26051, n26052, n26053,
         n26054, n26055, n26056, n26057, n26058, n26059, n260601, n26061,
         n26062, n26063, n26064, n26065, n26066, n26067, n26068, n26069,
         n260701, n26071, n26072, n26073, n26074, n26075, n26076, n26077,
         n26078, n26079, n260801, n26081, n26082, n26083, n26084, n26085,
         n26086, n26087, n26088, n26089, n260901, n26091, n26092, n26093,
         n26094, n26095, n26096, n26097, n26098, n26099, n261001, n26101,
         n26102, n26103, n26104, n26105, n26106, n26107, n26108, n26109,
         n261101, n26111, n26112, n26113, n26114, n26115, n26116, n26117,
         n26118, n26119, n261201, n26121, n26122, n26123, n26124, n26125,
         n26126, n26127, n26128, n26129, n26130, n26131, n26132, n26133,
         n26134, n26135, n26136, n26137, n26138, n26139, n26140, n26141,
         n26142, n26143, n26144, n26145, n26146, n26147, n26148, n26149,
         n26150, n26151, n26152, n26153, n26154, n26155, n26156, n26157,
         n26158, n26159, n26160, n26161, n26162, n26163, n26164, n26165,
         n26166, n26167, n26168, n26169, n26170, n26171, n26172, n26173,
         n26174, n26175, n26176, n26177, n26178, n26179, n26180, n26181,
         n26182, n26183, n26184, n26185, n26186, n26187, n26188, n26189,
         n26190, n26191, n26192, n26193, n26194, n26195, n26196, n26197,
         n26198, n26199, n26200, n26201, n26202, n26203, n26204, n26205,
         n26206, n26207, n26208, n26209, n26210, n26211, n26212, n26213,
         n26214, n26215, n26216, n26217, n26218, n26219, n26220, n26221,
         n26222, n26223, n26224, n26225, n26226, n26227, n26228, n26229,
         n26230, n26231, n26232, n26233, n26234, n26235, n26236, n26237,
         n26238, n26239, n26240, n26241, n26242, n26243, n26244, n26245,
         n26246, n26247, n26248, n26249, n26250, n26251, n26252, n26253,
         n26254, n26255, n26256, n26257, n26258, n26259, n26260, n26261,
         n26262, n26263, n26264, n26265, n26266, n26267, n26268, n26269,
         n26270, n26271, n26272, n26273, n26274, n26275, n26276, n26277,
         n26278, n26279, n26280, n26281, n26282, n26283, n26284, n26285,
         n26286, n26287, n26288, n26289, n26290, n26291, n26292, n26293,
         n26294, n26295, n26296, n26297, n26298, n26299, n26300, n26301,
         n26302, n26303, n26304, n26305, n26306, n26307, n26308, n26309,
         n26310, n26311, n26312, n26313, n26314, n26315, n26316, n26317,
         n26318, n26319, n26320, n26321, n26322, n26323, n26324, n26325,
         n26326, n26327, n26328, n26329, n26330, n26331, n26332, n26333,
         n26334, n26335, n26336, n26337, n26338, n26339, n26340, n26341,
         n26342, n26343, n26344, n26345, n26346, n26347, n26348, n26349,
         n26350, n26351, n26352, n26353, n26354, n26355, n26356, n26357,
         n26358, n26359, n26360, n26361, n26362, n26363, n26364, n26365,
         n26366, n26367, n26368, n26369, n263701, n26371, n26372, n26373,
         n26374, n26375, n26376, n26377, n26378, n26379, n26380, n26381,
         n26382, n26383, n26384, n26385, n26386, n26387, n26388, n26389,
         n26390, n26391, n26392, n26393, n26394, n26395, n26396, n26397,
         n26398, n26399, n26400, n26401, n26402, n26403, n26404, n26405,
         n26406, n26407, n26408, n26409, n264101, n26411, n26412, n26413,
         n26414, n26415, n26416, n26417, n26418, n26419, n264201, n26421,
         n26422, n26423, n26424, n26425, n26426, n26427, n26428, n26429,
         n264301, n26431, n26432, n26433, n26434, n26435, n26436, n26437,
         n26438, n26439, n264401, n26441, n26442, n26443, n26444, n26445,
         n26446, n26447, n26448, n26449, n264501, n26451, n26452, n26453,
         n26454, n26455, n26456, n26457, n26458, n26459, n264601, n26461,
         n26462, n26463, n26464, n26465, n26466, n26467, n26468, n26469,
         n264701, n26471, n26472, n26473, n26474, n26475, n26476, n26477,
         n26478, n26479, n264801, n26481, n26482, n26483, n26484, n26485,
         n26486, n26487, n26488, n26489, n264901, n26491, n26492, n26493,
         n26494, n26495, n26496, n26497, n26498, n26499, n265001, n26501,
         n26502, n26503, n26504, n26505, n26506, n26507, n26508, n26509,
         n265101, n26511, n26512, n26513, n26514, n26515, n26516, n26517,
         n26518, n26519, n265201, n26521, n26522, n26523, n26524, n26525,
         n26526, n26527, n26528, n26529, n265301, n26531, n26532, n26533,
         n26534, n26535, n26536, n26537, n26538, n26539, n265401, n26541,
         n26542, n26543, n26544, n26545, n26546, n26547, n26548, n26549,
         n265501, n26551, n26552, n26553, n26554, n26555, n26556, n26557,
         n26558, n26559, n265601, n26561, n26562, n26563, n26564, n26565,
         n26566, n26567, n26568, n26569, n26570, n26571, n26572, n26573,
         n26574, n26575, n26576, n26577, n26578, n26579, n26580, n26581,
         n26582, n26583, n26584, n26585, n26586, n26587, n26588, n26589,
         n26590, n26591, n26592, n26593, n26594, n26595, n26596, n26597,
         n26598, n26599, n26600, n26601, n26602, n26603, n26604, n26605,
         n26606, n26607, n26608, n26609, n26610, n26611, n26612, n26613,
         n26614, n26615, n26616, n26617, n26618, n26619, n26620, n26621,
         n26622, n26623, n26624, n26625, n26626, n26627, n26628, n26629,
         n26630, n26631, n26632, n26633, n26634, n26635, n26636, n26637,
         n26638, n26639, n26640, n26641, n26642, n26643, n26644, n26645,
         n26646, n26647, n26648, n26649, n26650, n26651, n26652, n26653,
         n26654, n26655, n26656, n26657, n26658, n26659, n26660, n26661,
         n26662, n26663, n26664, n26665, n26666, n26667, n26668, n26669,
         n26670, n26671, n26672, n26673, n26674, n26675, n26676, n26677,
         n26678, n26679, n26680, n26681, n26682, n26683, n26684, n26685,
         n26686, n26687, n26688, n26689, n26690, n26691, n26692, n26693,
         n26694, n26695, n26696, n26697, n26698, n26699, n26700, n26701,
         n26702, n26703, n26704, n26705, n26706, n26707, n26708, n26709,
         n26710, n26711, n26712, n26713, n26714, n26715, n26716, n26717,
         n26718, n26719, n26720, n26721, n26722, n26723, n26724, n26725,
         n26726, n26727, n26728, n26729, n26730, n26731, n26732, n26733,
         n26734, n26735, n26736, n26737, n26738, n26739, n267401, n26741,
         n26742, n26743, n26744, n26745, n26746, n26747, n26748, n26749,
         n267501, n26751, n26752, n26753, n26754, n26755, n26756, n26757,
         n26758, n26759, n267601, n26761, n26762, n26763, n26764, n26765,
         n26766, n26767, n26768, n26769, n267701, n26771, n26772, n26773,
         n26774, n26775, n26776, n26777, n26778, n26779, n267801, n26781,
         n26782, n26783, n26784, n26785, n26786, n26787, n26788, n26789,
         n267901, n26791, n26792, n26793, n26794, n26795, n26796, n26797,
         n26798, n26799, n268001, n26801, n26802, n26803, n26804, n26805,
         n26806, n26807, n26808, n26809, n268101, n26811, n26812, n26813,
         n26814, n26815, n26816, n26817, n26818, n26819, n268201, n26821,
         n26822, n26823, n26824, n26825, n26826, n26827, n26828, n26829,
         n268301, n26831, n26832, n26833, n26834, n26835, n26836, n26837,
         n26838, n26839, n268401, n26841, n26842, n26843, n26844, n26845,
         n26846, n26847, n26848, n26849, n268501, n26851, n26852, n26853,
         n26854, n26855, n26856, n26857, n26858, n26859, n268601, n26861,
         n26862, n26863, n26864, n26865, n26866, n26867, n26868, n26869,
         n268701, n26871, n26872, n26873, n26874, n26875, n26876, n26877,
         n26878, n26879, n268801, n26881, n26882, n26883, n26884, n26885,
         n26886, n26887, n26888, n26889, n268901, n26891, n26892, n26893,
         n26894, n26895, n26896, n26897, n26898, n26899, n269001, n26901,
         n26902, n26903, n26904, n26905, n26906, n26907, n26908, n26909,
         n269101, n26911, n26912, n26913, n26914, n26915, n26916, n26917,
         n26918, n26919, n269201, n26921, n26922, n26923, n26924, n26925,
         n26926, n26927, n26928, n26929, n269301, n26931, n26932, n26933,
         n26934, n26935, n26936, n26937, n26938, n26939, n269401, n26941,
         n26942, n26943, n26944, n26945, n26946, n26947, n26948, n26949,
         n26950, n26951, n26952, n26953, n26954, n26955, n26956, n26957,
         n26958, n26959, n26960, n26961, n26962, n26963, n26964, n26965,
         n26966, n26967, n26968, n26969, n26970, n26971, n26972, n26973,
         n26974, n26975, n26976, n26977, n26978, n26979, n26980, n26981,
         n26982, n26983, n26984, n26985, n26986, n26987, n26988, n26989,
         n26990, n26991, n26992, n26993, n26994, n26995, n26996, n26997,
         n26998, n26999, n27000, n27001, n27002, n27003, n27004, n27005,
         n27006, n27007, n27008, n27009, n27010, n27011, n27012, n27013,
         n27014, n27015, n27016, n27017, n27018, n27019, n27020, n27021,
         n27022, n27023, n27024, n27025, n27026, n27027, n27028, n27029,
         n27030, n27031, n27032, n27033, n27034, n27035, n27036, n27037,
         n27038, n27039, n27040, n27041, n27042, n27043, n27044, n27045,
         n27046, n27047, n27048, n27049, n27050, n27051, n27052, n27053,
         n27054, n27055, n27056, n27057, n27058, n27059, n27060, n27061,
         n27062, n27063, n27064, n27065, n27066, n27067, n27068, n27069,
         n27070, n27071, n27072, n27073, n27074, n27075, n27076, n27077,
         n27078, n27079, n27080, n27081, n27082, n27083, n27084, n27085,
         n27086, n27087, n27088, n27089, n27090, n27091, n27092, n27093,
         n27094, n27095, n27096, n27097, n27098, n27099, n27100, n27101,
         n27102, n27103, n27104, n27105, n27106, n27107, n27108, n27109,
         n27110, n27111, n27112, n27113, n27114, n27115, n27116, n27117,
         n27118, n27119, n27120, n27121, n27122, n27123, n27124, n27125,
         n27126, n27127, n27128, n27129, n27130, n27131, n27132, n27133,
         n27134, n27135, n27136, n27137, n27138, n27139, n27140, n27141,
         n27142, n27143, n27144, n27145, n27146, n27147, n27148, n27149,
         n27150, n27151, n27152, n27153, n27154, n27155, n27156, n27157,
         n27158, n27159, n27160, n27161, n27162, n27163, n27164, n27165,
         n27166, n27167, n27168, n27169, n27170, n27171, n27172, n27173,
         n27174, n27175, n27176, n27177, n27178, n27179, n27180, n27181,
         n27182, n27183, n27184, n27185, n27186, n27187, n27188, n27189,
         n27190, n27191, n27192, n27193, n27194, n27195, n27196, n27197,
         n27198, n27199, n27200, n27201, n27202, n27203, n27204, n27205,
         n27206, n27207, n27208, n27209, n27210, n27211, n27212, n27213,
         n27214, n27215, n27216, n27217, n27218, n27219, n27220, n27221,
         n27222, n27223, n27224, n27225, n27226, n27227, n27228, n27229,
         n27230, n27231, n27232, n27233, n27234, n27235, n27236, n27237,
         n27238, n27239, n27240, n27241, n27242, n27243, n27244, n27245,
         n27246, n27247, n27248, n27249, n27250, n27251, n27252, n27253,
         n27254, n27255, n27256, n27257, n27258, n27259, n27260, n27261,
         n27262, n27263, n27264, n27265, n27266, n27267, n27268, n27269,
         n27270, n27271, n27272, n27273, n27274, n27275, n27276, n27277,
         n27278, n27279, n27280, n27281, n27282, n27283, n27284, n27285,
         n27286, n27287, n27288, n27289, n272901, n27291, n27292, n27293,
         n27294, n27295, n27296, n27297, n27298, n27299, n27300, n27301,
         n27302, n27303, n27304, n27305, n27306, n27307, n27308, n27309,
         n27310, n27311, n27312, n27313, n27314, n27315, n27316, n27317,
         n27318, n27319, n27320, n27321, n27322, n27323, n27324, n27325,
         n27326, n27327, n27328, n27329, n273301, n27331, n27332, n27333,
         n27334, n27335, n27336, n27337, n27338, n27339, n273401, n27341,
         n27342, n27343, n27344, n27345, n27346, n27347, n27348, n27349,
         n273501, n27351, n27352, n27353, n27354, n27355, n27356, n27357,
         n27358, n27359, n273601, n27361, n27362, n27363, n27364, n27365,
         n27366, n27367, n27368, n27369, n273701, n27371, n27372, n27373,
         n27374, n27375, n27376, n27377, n27378, n27379, n273801, n27381,
         n27382, n27383, n27384, n27385, n27386, n27387, n27388, n27389,
         n273901, n27391, n27392, n27393, n27394, n27395, n27396, n27397,
         n27398, n27399, n274001, n27401, n27402, n27403, n27404, n27405,
         n27406, n27407, n27408, n27409, n274101, n27411, n27412, n27413,
         n27414, n27415, n27416, n27417, n27418, n27419, n274201, n27421,
         n27422, n27423, n27424, n27425, n27426, n27427, n27428, n27429,
         n274301, n27431, n27432, n27433, n27434, n27435, n27436, n27437,
         n27438, n27439, n274401, n27441, n27442, n27443, n27444, n27445,
         n27446, n27447, n27448, n27449, n274501, n27451, n27452, n27453,
         n27454, n27455, n27456, n27457, n27458, n27459, n274601, n27461,
         n27462, n27463, n27464, n27465, n27466, n27467, n27468, n27469,
         n274701, n27471, n27472, n27473, n27474, n27475, n27476, n27477,
         n27478, n27479, n274801, n27481, n27482, n27483, n27484, n27485,
         n27486, n27487, n27488, n27489, n27490, n27491, n27492, n27493,
         n27494, n27495, n27496, n27497, n27498, n27499, n27500, n27501,
         n27502, n27503, n27504, n27505, n27506, n27507, n27508, n27509,
         n27510, n27511, n27512, n27513, n27514, n27515, n27516, n27517,
         n27518, n27519, n27520, n27521, n27522, n27523, n27524, n27525,
         n27526, n27527, n27528, n27529, n27530, n27531, n27532, n27533,
         n27534, n27535, n27536, n27537, n27538, n27539, n27540, n27541,
         n27542, n27543, n27544, n27545, n27546, n27547, n27548, n27549,
         n27550, n27551, n27552, n27553, n27554, n27555, n27556, n27557,
         n27558, n27559, n27560, n27561, n27562, n27563, n27564, n27565,
         n27566, n27567, n27568, n27569, n27570, n27571, n27572, n27573,
         n27574, n27575, n27576, n27577, n27578, n27579, n27580, n27581,
         n27582, n27583, n27584, n27585, n27586, n27587, n27588, n27589,
         n27590, n27591, n27592, n27593, n27594, n27595, n27596, n27597,
         n27598, n27599, n27600, n27601, n27602, n27603, n27604, n27605,
         n27606, n27607, n27608, n27609, n27610, n27611, n27612, n27613,
         n27614, n27615, n27616, n27617, n27618, n27619, n27620, n27621,
         n27622, n27623, n27624, n27625, n27626, n27627, n27628, n27629,
         n27630, n27631, n27632, n27633, n27634, n27635, n27636, n27637,
         n27638, n27639, n27640, n27641, n27642, n27643, n27644, n27645,
         n27646, n27647, n27648, n27649, n27650, n27651, n27652, n27653,
         n27654, n27655, n27656, n27657, n27658, n27659, n276601, n27661,
         n27662, n27663, n27664, n27665, n27666, n27667, n27668, n27669,
         n276701, n27671, n27672, n27673, n27674, n27675, n27676, n27677,
         n27678, n27679, n276801, n27681, n27682, n27683, n27684, n27685,
         n27686, n27687, n27688, n27689, n276901, n27691, n27692, n27693,
         n27694, n27695, n27696, n27697, n27698, n27699, n277001, n27701,
         n27702, n27703, n27704, n27705, n27706, n27707, n27708, n27709,
         n277101, n27711, n27712, n27713, n27714, n27715, n27716, n27717,
         n27718, n27719, n277201, n27721, n27722, n27723, n27724, n27725,
         n27726, n27727, n27728, n27729, n277301, n27731, n27732, n27733,
         n27734, n27735, n27736, n27737, n27738, n27739, n277401, n27741,
         n27742, n27743, n27744, n27745, n27746, n27747, n27748, n27749,
         n277501, n27751, n27752, n27753, n27754, n27755, n27756, n27757,
         n27758, n27759, n277601, n27761, n27762, n27763, n27764, n27765,
         n27766, n27767, n27768, n27769, n277701, n27771, n27772, n27773,
         n27774, n27775, n27776, n27777, n27778, n27779, n277801, n27781,
         n27782, n27783, n27784, n27785, n27786, n27787, n27788, n27789,
         n277901, n27791, n27792, n27793, n27794, n27795, n27796, n27797,
         n27798, n27799, n278001, n27801, n27802, n27803, n27804, n27805,
         n27806, n27807, n27808, n27809, n278101, n27811, n27812, n27813,
         n27814, n27815, n27816, n27817, n27818, n27819, n278201, n27821,
         n27822, n27823, n27824, n27825, n27826, n27827, n27828, n27829,
         n278301, n27831, n27832, n27833, n27834, n27835, n27836, n27837,
         n27838, n27839, n278401, n27841, n27842, n27843, n27844, n27845,
         n27846, n27847, n27848, n27849, n278501, n27851, n27852, n27853,
         n27854, n27855, n27856, n27857, n27858, n27859, n278601, n27861,
         n27862, n27863, n27864, n27865, n27866, n27867, n27868, n27869,
         n27870, n27871, n27872, n27873, n27874, n27875, n27876, n27877,
         n27878, n27879, n27880, n27881, n27882, n27883, n27884, n27885,
         n27886, n27887, n27888, n27889, n27890, n27891, n27892, n27893,
         n27894, n27895, n27896, n27897, n27898, n27899, n27900, n27901,
         n27902, n27903, n27904, n27905, n27906, n27907, n27908, n27909,
         n27910, n27911, n27912, n27913, n27914, n27915, n27916, n27917,
         n27918, n27919, n27920, n27921, n27922, n27923, n27924, n27925,
         n27926, n27927, n27928, n27929, n27930, n27931, n27932, n27933,
         n27934, n27935, n27936, n27937, n27938, n27939, n27940, n27941,
         n27942, n27943, n27944, n27945, n27946, n27947, n27948;
  wire   [5:3] upper_bound;
  wire   [5:4] sub_127_aco_carry;

  DFF_X1 data_queue_reg_0__0__7_ ( .D(n16772), .CK(clk), .Q(
        data_queue_0__0__7_), .QN(n949) );
  DFF_X1 data_queue_reg_0__0__6_ ( .D(n16767), .CK(clk), .Q(
        data_queue_0__0__6_), .QN(n950) );
  DFF_X1 data_queue_reg_0__0__5_ ( .D(n16762), .CK(clk), .Q(
        data_queue_0__0__5_), .QN(n951) );
  DFF_X1 data_queue_reg_0__0__4_ ( .D(n16757), .CK(clk), .Q(
        data_queue_0__0__4_), .QN(n952) );
  DFF_X1 data_queue_reg_0__0__3_ ( .D(n16752), .CK(clk), .Q(
        data_queue_0__0__3_), .QN(n953) );
  DFF_X1 data_queue_reg_0__0__2_ ( .D(n16747), .CK(clk), .Q(
        data_queue_0__0__2_), .QN(n954) );
  DFF_X1 data_queue_reg_0__0__1_ ( .D(n16742), .CK(clk), .Q(
        data_queue_0__0__1_), .QN(n955) );
  DFF_X1 data_queue_reg_0__0__0_ ( .D(n16737), .CK(clk), .Q(
        data_queue_0__0__0_), .QN(n956) );
  DFF_X1 data_queue_reg_0__1__7_ ( .D(n16732), .CK(clk), .Q(
        data_queue_0__1__7_), .QN(n957) );
  DFF_X1 data_queue_reg_0__1__6_ ( .D(n16727), .CK(clk), .Q(
        data_queue_0__1__6_), .QN(n958) );
  DFF_X1 data_queue_reg_0__1__5_ ( .D(n16722), .CK(clk), .Q(
        data_queue_0__1__5_), .QN(n959) );
  DFF_X1 data_queue_reg_0__1__4_ ( .D(n16717), .CK(clk), .Q(
        data_queue_0__1__4_), .QN(n960) );
  DFF_X1 data_queue_reg_0__1__3_ ( .D(n16712), .CK(clk), .Q(
        data_queue_0__1__3_), .QN(n961) );
  DFF_X1 data_queue_reg_0__1__2_ ( .D(n16707), .CK(clk), .Q(
        data_queue_0__1__2_), .QN(n962) );
  DFF_X1 data_queue_reg_0__1__1_ ( .D(n16702), .CK(clk), .Q(
        data_queue_0__1__1_), .QN(n963) );
  DFF_X1 data_queue_reg_0__1__0_ ( .D(n16697), .CK(clk), .Q(
        data_queue_0__1__0_), .QN(n964) );
  DFF_X1 data_queue_reg_0__2__7_ ( .D(n16692), .CK(clk), .Q(
        data_queue_0__2__7_), .QN(n965) );
  DFF_X1 data_queue_reg_0__2__6_ ( .D(n16687), .CK(clk), .Q(
        data_queue_0__2__6_), .QN(n966) );
  DFF_X1 data_queue_reg_0__2__5_ ( .D(n16682), .CK(clk), .Q(
        data_queue_0__2__5_), .QN(n967) );
  DFF_X1 data_queue_reg_0__2__4_ ( .D(n16677), .CK(clk), .Q(
        data_queue_0__2__4_), .QN(n968) );
  DFF_X1 data_queue_reg_0__2__3_ ( .D(n16672), .CK(clk), .Q(
        data_queue_0__2__3_), .QN(n969) );
  DFF_X1 data_queue_reg_0__2__2_ ( .D(n16667), .CK(clk), .Q(
        data_queue_0__2__2_), .QN(n970) );
  DFF_X1 data_queue_reg_0__2__1_ ( .D(n16662), .CK(clk), .Q(
        data_queue_0__2__1_), .QN(n971) );
  DFF_X1 data_queue_reg_0__2__0_ ( .D(n16657), .CK(clk), .Q(
        data_queue_0__2__0_), .QN(n972) );
  DFF_X1 data_queue_reg_0__3__7_ ( .D(n16652), .CK(clk), .Q(
        data_queue_0__3__7_), .QN(n973) );
  DFF_X1 data_queue_reg_0__3__6_ ( .D(n16647), .CK(clk), .Q(
        data_queue_0__3__6_), .QN(n974) );
  DFF_X1 data_queue_reg_0__3__5_ ( .D(n16642), .CK(clk), .Q(
        data_queue_0__3__5_), .QN(n975) );
  DFF_X1 data_queue_reg_0__3__4_ ( .D(n16637), .CK(clk), .Q(
        data_queue_0__3__4_), .QN(n976) );
  DFF_X1 data_queue_reg_0__3__3_ ( .D(n16632), .CK(clk), .Q(
        data_queue_0__3__3_), .QN(n977) );
  DFF_X1 data_queue_reg_0__3__2_ ( .D(n16627), .CK(clk), .Q(
        data_queue_0__3__2_), .QN(n978) );
  DFF_X1 data_queue_reg_0__3__1_ ( .D(n16622), .CK(clk), .Q(
        data_queue_0__3__1_), .QN(n979) );
  DFF_X1 data_queue_reg_0__3__0_ ( .D(n16617), .CK(clk), .Q(
        data_queue_0__3__0_), .QN(n980) );
  DFF_X1 data_queue_reg_0__4__7_ ( .D(n16612), .CK(clk), .Q(
        data_queue_0__4__7_), .QN(n981) );
  DFF_X1 data_queue_reg_0__4__6_ ( .D(n16607), .CK(clk), .Q(
        data_queue_0__4__6_), .QN(n982) );
  DFF_X1 data_queue_reg_0__4__5_ ( .D(n16602), .CK(clk), .Q(
        data_queue_0__4__5_), .QN(n983) );
  DFF_X1 data_queue_reg_0__4__4_ ( .D(n16597), .CK(clk), .Q(
        data_queue_0__4__4_), .QN(n984) );
  DFF_X1 data_queue_reg_0__4__3_ ( .D(n16592), .CK(clk), .Q(
        data_queue_0__4__3_), .QN(n985) );
  DFF_X1 data_queue_reg_0__4__2_ ( .D(n16587), .CK(clk), .Q(
        data_queue_0__4__2_), .QN(n986) );
  DFF_X1 data_queue_reg_0__4__1_ ( .D(n16582), .CK(clk), .Q(
        data_queue_0__4__1_), .QN(n987) );
  DFF_X1 data_queue_reg_0__4__0_ ( .D(n16577), .CK(clk), .Q(
        data_queue_0__4__0_), .QN(n988) );
  DFF_X1 data_queue_reg_0__5__7_ ( .D(n16572), .CK(clk), .Q(
        data_queue_0__5__7_), .QN(n989) );
  DFF_X1 data_queue_reg_0__5__6_ ( .D(n16567), .CK(clk), .Q(
        data_queue_0__5__6_), .QN(n990) );
  DFF_X1 data_queue_reg_0__5__5_ ( .D(n16562), .CK(clk), .Q(
        data_queue_0__5__5_), .QN(n991) );
  DFF_X1 data_queue_reg_0__5__4_ ( .D(n16557), .CK(clk), .Q(
        data_queue_0__5__4_), .QN(n992) );
  DFF_X1 data_queue_reg_0__5__3_ ( .D(n16552), .CK(clk), .Q(
        data_queue_0__5__3_), .QN(n993) );
  DFF_X1 data_queue_reg_0__5__2_ ( .D(n16547), .CK(clk), .Q(
        data_queue_0__5__2_), .QN(n994) );
  DFF_X1 data_queue_reg_0__5__1_ ( .D(n16542), .CK(clk), .Q(
        data_queue_0__5__1_), .QN(n995) );
  DFF_X1 data_queue_reg_0__5__0_ ( .D(n16537), .CK(clk), .Q(
        data_queue_0__5__0_), .QN(n996) );
  DFF_X1 data_queue_reg_0__6__7_ ( .D(n16530), .CK(clk), .Q(
        data_queue_0__6__7_), .QN(n997) );
  DFF_X1 data_queue_reg_0__6__6_ ( .D(n16523), .CK(clk), .Q(
        data_queue_0__6__6_), .QN(n998) );
  DFF_X1 data_queue_reg_0__6__5_ ( .D(n16516), .CK(clk), .Q(
        data_queue_0__6__5_), .QN(n999) );
  DFF_X1 data_queue_reg_0__6__4_ ( .D(n16509), .CK(clk), .Q(
        data_queue_0__6__4_), .QN(n1000) );
  DFF_X1 data_queue_reg_0__6__3_ ( .D(n16502), .CK(clk), .Q(
        data_queue_0__6__3_), .QN(n1001) );
  DFF_X1 data_queue_reg_0__6__2_ ( .D(n16495), .CK(clk), .Q(
        data_queue_0__6__2_), .QN(n1002) );
  DFF_X1 data_queue_reg_0__6__1_ ( .D(n16488), .CK(clk), .Q(
        data_queue_0__6__1_), .QN(n1003) );
  DFF_X1 data_queue_reg_0__6__0_ ( .D(n16481), .CK(clk), .Q(
        data_queue_0__6__0_), .QN(n1004) );
  DFF_X1 data_queue_reg_0__7__7_ ( .D(n16480), .CK(clk), .Q(
        data_queue_0__7__7_), .QN(n17264) );
  DFF_X1 data_queue_reg_0__7__6_ ( .D(n16477), .CK(clk), .Q(
        data_queue_0__7__6_), .QN(n17263) );
  DFF_X1 data_queue_reg_0__7__5_ ( .D(n16474), .CK(clk), .Q(
        data_queue_0__7__5_), .QN(n17262) );
  DFF_X1 data_queue_reg_0__7__4_ ( .D(n16471), .CK(clk), .Q(
        data_queue_0__7__4_), .QN(n17261) );
  DFF_X1 data_queue_reg_0__7__3_ ( .D(n16468), .CK(clk), .Q(
        data_queue_0__7__3_), .QN(n17260) );
  DFF_X1 data_queue_reg_0__7__2_ ( .D(n16465), .CK(clk), .Q(
        data_queue_0__7__2_), .QN(n17259) );
  DFF_X1 data_queue_reg_0__7__1_ ( .D(n16462), .CK(clk), .Q(
        data_queue_0__7__1_), .QN(n17258) );
  DFF_X1 data_queue_reg_0__7__0_ ( .D(n16459), .CK(clk), .Q(
        data_queue_0__7__0_), .QN(n17257) );
  DFF_X1 data_queue_reg_1__0__7_ ( .D(n16452), .CK(clk), .Q(
        data_queue_1__0__7_), .QN(n1005) );
  DFF_X1 data_queue_reg_1__0__6_ ( .D(n16447), .CK(clk), .Q(
        data_queue_1__0__6_), .QN(n1006) );
  DFF_X1 data_queue_reg_1__0__5_ ( .D(n16442), .CK(clk), .Q(
        data_queue_1__0__5_), .QN(n1007) );
  DFF_X1 data_queue_reg_1__0__4_ ( .D(n16437), .CK(clk), .Q(
        data_queue_1__0__4_), .QN(n1008) );
  DFF_X1 data_queue_reg_1__0__3_ ( .D(n16432), .CK(clk), .Q(
        data_queue_1__0__3_), .QN(n1009) );
  DFF_X1 data_queue_reg_1__0__2_ ( .D(n16427), .CK(clk), .Q(
        data_queue_1__0__2_), .QN(n1010) );
  DFF_X1 data_queue_reg_1__0__1_ ( .D(n16422), .CK(clk), .Q(
        data_queue_1__0__1_), .QN(n1011) );
  DFF_X1 data_queue_reg_1__0__0_ ( .D(n16417), .CK(clk), .Q(
        data_queue_1__0__0_), .QN(n1012) );
  DFF_X1 data_queue_reg_1__1__7_ ( .D(n16412), .CK(clk), .Q(
        data_queue_1__1__7_), .QN(n1013) );
  DFF_X1 data_queue_reg_1__1__6_ ( .D(n16407), .CK(clk), .Q(
        data_queue_1__1__6_), .QN(n1014) );
  DFF_X1 data_queue_reg_1__1__5_ ( .D(n16402), .CK(clk), .Q(
        data_queue_1__1__5_), .QN(n1015) );
  DFF_X1 data_queue_reg_1__1__4_ ( .D(n16397), .CK(clk), .Q(
        data_queue_1__1__4_), .QN(n1016) );
  DFF_X1 data_queue_reg_1__1__3_ ( .D(n16392), .CK(clk), .Q(
        data_queue_1__1__3_), .QN(n1017) );
  DFF_X1 data_queue_reg_1__1__2_ ( .D(n16387), .CK(clk), .Q(
        data_queue_1__1__2_), .QN(n1018) );
  DFF_X1 data_queue_reg_1__1__1_ ( .D(n16382), .CK(clk), .Q(
        data_queue_1__1__1_), .QN(n1019) );
  DFF_X1 data_queue_reg_1__1__0_ ( .D(n16377), .CK(clk), .Q(
        data_queue_1__1__0_), .QN(n1020) );
  DFF_X1 data_queue_reg_1__2__7_ ( .D(n16372), .CK(clk), .Q(
        data_queue_1__2__7_), .QN(n1021) );
  DFF_X1 data_queue_reg_1__2__6_ ( .D(n16367), .CK(clk), .Q(
        data_queue_1__2__6_), .QN(n1022) );
  DFF_X1 data_queue_reg_1__2__5_ ( .D(n16362), .CK(clk), .Q(
        data_queue_1__2__5_), .QN(n1023) );
  DFF_X1 data_queue_reg_1__2__4_ ( .D(n16357), .CK(clk), .Q(
        data_queue_1__2__4_), .QN(n1024) );
  DFF_X1 data_queue_reg_1__2__3_ ( .D(n16352), .CK(clk), .Q(
        data_queue_1__2__3_), .QN(n1025) );
  DFF_X1 data_queue_reg_1__2__2_ ( .D(n16347), .CK(clk), .Q(
        data_queue_1__2__2_), .QN(n1026) );
  DFF_X1 data_queue_reg_1__2__1_ ( .D(n16342), .CK(clk), .Q(
        data_queue_1__2__1_), .QN(n1027) );
  DFF_X1 data_queue_reg_1__2__0_ ( .D(n16337), .CK(clk), .Q(
        data_queue_1__2__0_), .QN(n1028) );
  DFF_X1 data_queue_reg_1__3__7_ ( .D(n16332), .CK(clk), .Q(
        data_queue_1__3__7_), .QN(n1029) );
  DFF_X1 data_queue_reg_1__3__6_ ( .D(n16327), .CK(clk), .Q(
        data_queue_1__3__6_), .QN(n1030) );
  DFF_X1 data_queue_reg_1__3__5_ ( .D(n16322), .CK(clk), .Q(
        data_queue_1__3__5_), .QN(n1031) );
  DFF_X1 data_queue_reg_1__3__4_ ( .D(n16317), .CK(clk), .Q(
        data_queue_1__3__4_), .QN(n1032) );
  DFF_X1 data_queue_reg_1__3__3_ ( .D(n16312), .CK(clk), .Q(
        data_queue_1__3__3_), .QN(n1033) );
  DFF_X1 data_queue_reg_1__3__2_ ( .D(n16307), .CK(clk), .Q(
        data_queue_1__3__2_), .QN(n1034) );
  DFF_X1 data_queue_reg_1__3__1_ ( .D(n16302), .CK(clk), .Q(
        data_queue_1__3__1_), .QN(n1035) );
  DFF_X1 data_queue_reg_1__3__0_ ( .D(n16297), .CK(clk), .Q(
        data_queue_1__3__0_), .QN(n1036) );
  DFF_X1 data_queue_reg_1__4__7_ ( .D(n16292), .CK(clk), .Q(
        data_queue_1__4__7_), .QN(n1037) );
  DFF_X1 data_queue_reg_1__4__6_ ( .D(n16287), .CK(clk), .Q(
        data_queue_1__4__6_), .QN(n1038) );
  DFF_X1 data_queue_reg_1__4__5_ ( .D(n16282), .CK(clk), .Q(
        data_queue_1__4__5_), .QN(n1039) );
  DFF_X1 data_queue_reg_1__4__4_ ( .D(n16277), .CK(clk), .Q(
        data_queue_1__4__4_), .QN(n1040) );
  DFF_X1 data_queue_reg_1__4__3_ ( .D(n16272), .CK(clk), .Q(
        data_queue_1__4__3_), .QN(n1041) );
  DFF_X1 data_queue_reg_1__4__2_ ( .D(n16267), .CK(clk), .Q(
        data_queue_1__4__2_), .QN(n1042) );
  DFF_X1 data_queue_reg_1__4__1_ ( .D(n16262), .CK(clk), .Q(
        data_queue_1__4__1_), .QN(n1043) );
  DFF_X1 data_queue_reg_1__4__0_ ( .D(n16257), .CK(clk), .Q(
        data_queue_1__4__0_), .QN(n1044) );
  DFF_X1 data_queue_reg_1__5__7_ ( .D(n16252), .CK(clk), .Q(
        data_queue_1__5__7_), .QN(n1045) );
  DFF_X1 data_queue_reg_1__5__6_ ( .D(n16247), .CK(clk), .Q(
        data_queue_1__5__6_), .QN(n1046) );
  DFF_X1 data_queue_reg_1__5__5_ ( .D(n16242), .CK(clk), .Q(
        data_queue_1__5__5_), .QN(n1047) );
  DFF_X1 data_queue_reg_1__5__4_ ( .D(n16237), .CK(clk), .Q(
        data_queue_1__5__4_), .QN(n1048) );
  DFF_X1 data_queue_reg_1__5__3_ ( .D(n16232), .CK(clk), .Q(
        data_queue_1__5__3_), .QN(n1049) );
  DFF_X1 data_queue_reg_1__5__2_ ( .D(n16227), .CK(clk), .Q(
        data_queue_1__5__2_), .QN(n1050) );
  DFF_X1 data_queue_reg_1__5__1_ ( .D(n16222), .CK(clk), .Q(
        data_queue_1__5__1_), .QN(n1051) );
  DFF_X1 data_queue_reg_1__5__0_ ( .D(n16217), .CK(clk), .Q(
        data_queue_1__5__0_), .QN(n1052) );
  DFF_X1 data_queue_reg_1__6__7_ ( .D(n16210), .CK(clk), .Q(
        data_queue_1__6__7_), .QN(n1053) );
  DFF_X1 data_queue_reg_1__6__6_ ( .D(n16203), .CK(clk), .Q(
        data_queue_1__6__6_), .QN(n1054) );
  DFF_X1 data_queue_reg_1__6__5_ ( .D(n16196), .CK(clk), .Q(
        data_queue_1__6__5_), .QN(n1055) );
  DFF_X1 data_queue_reg_1__6__4_ ( .D(n16189), .CK(clk), .Q(
        data_queue_1__6__4_), .QN(n1056) );
  DFF_X1 data_queue_reg_1__6__3_ ( .D(n16182), .CK(clk), .Q(
        data_queue_1__6__3_), .QN(n1057) );
  DFF_X1 data_queue_reg_1__6__2_ ( .D(n16175), .CK(clk), .Q(
        data_queue_1__6__2_), .QN(n1058) );
  DFF_X1 data_queue_reg_1__6__1_ ( .D(n16168), .CK(clk), .Q(
        data_queue_1__6__1_), .QN(n1059) );
  DFF_X1 data_queue_reg_1__6__0_ ( .D(n16161), .CK(clk), .Q(
        data_queue_1__6__0_), .QN(n1060) );
  DFF_X1 data_queue_reg_1__7__7_ ( .D(n16160), .CK(clk), .Q(
        data_queue_1__7__7_), .QN(n17256) );
  DFF_X1 data_queue_reg_1__7__6_ ( .D(n16157), .CK(clk), .Q(
        data_queue_1__7__6_), .QN(n17255) );
  DFF_X1 data_queue_reg_1__7__5_ ( .D(n16154), .CK(clk), .Q(
        data_queue_1__7__5_), .QN(n17254) );
  DFF_X1 data_queue_reg_1__7__4_ ( .D(n16151), .CK(clk), .Q(
        data_queue_1__7__4_), .QN(n17253) );
  DFF_X1 data_queue_reg_1__7__3_ ( .D(n16148), .CK(clk), .Q(
        data_queue_1__7__3_), .QN(n17252) );
  DFF_X1 data_queue_reg_1__7__2_ ( .D(n16145), .CK(clk), .Q(
        data_queue_1__7__2_), .QN(n17251) );
  DFF_X1 data_queue_reg_1__7__1_ ( .D(n16142), .CK(clk), .Q(
        data_queue_1__7__1_), .QN(n17250) );
  DFF_X1 data_queue_reg_1__7__0_ ( .D(n16139), .CK(clk), .Q(
        data_queue_1__7__0_), .QN(n17249) );
  DFF_X1 data_queue_reg_2__0__7_ ( .D(n16132), .CK(clk), .Q(
        data_queue_2__0__7_), .QN(n1061) );
  DFF_X1 data_queue_reg_2__0__6_ ( .D(n16127), .CK(clk), .Q(
        data_queue_2__0__6_), .QN(n1062) );
  DFF_X1 data_queue_reg_2__0__5_ ( .D(n16122), .CK(clk), .Q(
        data_queue_2__0__5_), .QN(n1063) );
  DFF_X1 data_queue_reg_2__0__4_ ( .D(n16117), .CK(clk), .Q(
        data_queue_2__0__4_), .QN(n1064) );
  DFF_X1 data_queue_reg_2__0__3_ ( .D(n16112), .CK(clk), .Q(
        data_queue_2__0__3_), .QN(n1065) );
  DFF_X1 data_queue_reg_2__0__2_ ( .D(n16107), .CK(clk), .Q(
        data_queue_2__0__2_), .QN(n1066) );
  DFF_X1 data_queue_reg_2__0__1_ ( .D(n16102), .CK(clk), .Q(
        data_queue_2__0__1_), .QN(n1067) );
  DFF_X1 data_queue_reg_2__0__0_ ( .D(n16097), .CK(clk), .Q(
        data_queue_2__0__0_), .QN(n1068) );
  DFF_X1 data_queue_reg_2__1__7_ ( .D(n16092), .CK(clk), .Q(
        data_queue_2__1__7_), .QN(n1069) );
  DFF_X1 data_queue_reg_2__1__6_ ( .D(n16087), .CK(clk), .Q(
        data_queue_2__1__6_), .QN(n1070) );
  DFF_X1 data_queue_reg_2__1__5_ ( .D(n16082), .CK(clk), .Q(
        data_queue_2__1__5_), .QN(n1071) );
  DFF_X1 data_queue_reg_2__1__4_ ( .D(n16077), .CK(clk), .Q(
        data_queue_2__1__4_), .QN(n1072) );
  DFF_X1 data_queue_reg_2__1__3_ ( .D(n16072), .CK(clk), .Q(
        data_queue_2__1__3_), .QN(n1073) );
  DFF_X1 data_queue_reg_2__1__2_ ( .D(n16067), .CK(clk), .Q(
        data_queue_2__1__2_), .QN(n1074) );
  DFF_X1 data_queue_reg_2__1__1_ ( .D(n16062), .CK(clk), .Q(
        data_queue_2__1__1_), .QN(n1075) );
  DFF_X1 data_queue_reg_2__1__0_ ( .D(n16057), .CK(clk), .Q(
        data_queue_2__1__0_), .QN(n1076) );
  DFF_X1 data_queue_reg_2__2__7_ ( .D(n16052), .CK(clk), .Q(
        data_queue_2__2__7_), .QN(n1077) );
  DFF_X1 data_queue_reg_2__2__6_ ( .D(n16047), .CK(clk), .Q(
        data_queue_2__2__6_), .QN(n1078) );
  DFF_X1 data_queue_reg_2__2__5_ ( .D(n16042), .CK(clk), .Q(
        data_queue_2__2__5_), .QN(n1079) );
  DFF_X1 data_queue_reg_2__2__4_ ( .D(n16037), .CK(clk), .Q(
        data_queue_2__2__4_), .QN(n1080) );
  DFF_X1 data_queue_reg_2__2__3_ ( .D(n16032), .CK(clk), .Q(
        data_queue_2__2__3_), .QN(n1081) );
  DFF_X1 data_queue_reg_2__2__2_ ( .D(n16027), .CK(clk), .Q(
        data_queue_2__2__2_), .QN(n1082) );
  DFF_X1 data_queue_reg_2__2__1_ ( .D(n16022), .CK(clk), .Q(
        data_queue_2__2__1_), .QN(n1083) );
  DFF_X1 data_queue_reg_2__2__0_ ( .D(n16017), .CK(clk), .Q(
        data_queue_2__2__0_), .QN(n1084) );
  DFF_X1 data_queue_reg_2__3__7_ ( .D(n16012), .CK(clk), .Q(
        data_queue_2__3__7_), .QN(n1085) );
  DFF_X1 data_queue_reg_2__3__6_ ( .D(n16007), .CK(clk), .Q(
        data_queue_2__3__6_), .QN(n1086) );
  DFF_X1 data_queue_reg_2__3__5_ ( .D(n16002), .CK(clk), .Q(
        data_queue_2__3__5_), .QN(n1087) );
  DFF_X1 data_queue_reg_2__3__4_ ( .D(n15997), .CK(clk), .Q(
        data_queue_2__3__4_), .QN(n1088) );
  DFF_X1 data_queue_reg_2__3__3_ ( .D(n15992), .CK(clk), .Q(
        data_queue_2__3__3_), .QN(n1089) );
  DFF_X1 data_queue_reg_2__3__2_ ( .D(n15987), .CK(clk), .Q(
        data_queue_2__3__2_), .QN(n1090) );
  DFF_X1 data_queue_reg_2__3__1_ ( .D(n15982), .CK(clk), .Q(
        data_queue_2__3__1_), .QN(n1091) );
  DFF_X1 data_queue_reg_2__3__0_ ( .D(n15977), .CK(clk), .Q(
        data_queue_2__3__0_), .QN(n1092) );
  DFF_X1 data_queue_reg_2__4__7_ ( .D(n15972), .CK(clk), .Q(
        data_queue_2__4__7_), .QN(n1093) );
  DFF_X1 data_queue_reg_2__4__6_ ( .D(n15967), .CK(clk), .Q(
        data_queue_2__4__6_), .QN(n1094) );
  DFF_X1 data_queue_reg_2__4__5_ ( .D(n15962), .CK(clk), .Q(
        data_queue_2__4__5_), .QN(n1095) );
  DFF_X1 data_queue_reg_2__4__4_ ( .D(n15957), .CK(clk), .Q(
        data_queue_2__4__4_), .QN(n1096) );
  DFF_X1 data_queue_reg_2__4__3_ ( .D(n15952), .CK(clk), .Q(
        data_queue_2__4__3_), .QN(n1097) );
  DFF_X1 data_queue_reg_2__4__2_ ( .D(n15947), .CK(clk), .Q(
        data_queue_2__4__2_), .QN(n1098) );
  DFF_X1 data_queue_reg_2__4__1_ ( .D(n15942), .CK(clk), .Q(
        data_queue_2__4__1_), .QN(n1099) );
  DFF_X1 data_queue_reg_2__4__0_ ( .D(n15937), .CK(clk), .Q(
        data_queue_2__4__0_), .QN(n1100) );
  DFF_X1 data_queue_reg_2__5__7_ ( .D(n15932), .CK(clk), .Q(
        data_queue_2__5__7_), .QN(n1101) );
  DFF_X1 data_queue_reg_2__5__6_ ( .D(n15927), .CK(clk), .Q(
        data_queue_2__5__6_), .QN(n1102) );
  DFF_X1 data_queue_reg_2__5__5_ ( .D(n15922), .CK(clk), .Q(
        data_queue_2__5__5_), .QN(n1103) );
  DFF_X1 data_queue_reg_2__5__4_ ( .D(n15917), .CK(clk), .Q(
        data_queue_2__5__4_), .QN(n1104) );
  DFF_X1 data_queue_reg_2__5__3_ ( .D(n15912), .CK(clk), .Q(
        data_queue_2__5__3_), .QN(n1105) );
  DFF_X1 data_queue_reg_2__5__2_ ( .D(n15907), .CK(clk), .Q(
        data_queue_2__5__2_), .QN(n1106) );
  DFF_X1 data_queue_reg_2__5__1_ ( .D(n15902), .CK(clk), .Q(
        data_queue_2__5__1_), .QN(n1107) );
  DFF_X1 data_queue_reg_2__5__0_ ( .D(n15897), .CK(clk), .Q(
        data_queue_2__5__0_), .QN(n1108) );
  DFF_X1 data_queue_reg_2__6__7_ ( .D(n15890), .CK(clk), .Q(
        data_queue_2__6__7_), .QN(n1109) );
  DFF_X1 data_queue_reg_2__6__6_ ( .D(n15883), .CK(clk), .Q(
        data_queue_2__6__6_), .QN(n1110) );
  DFF_X1 data_queue_reg_2__6__5_ ( .D(n15876), .CK(clk), .Q(
        data_queue_2__6__5_), .QN(n1111) );
  DFF_X1 data_queue_reg_2__6__4_ ( .D(n15869), .CK(clk), .Q(
        data_queue_2__6__4_), .QN(n1112) );
  DFF_X1 data_queue_reg_2__6__3_ ( .D(n15862), .CK(clk), .Q(
        data_queue_2__6__3_), .QN(n1113) );
  DFF_X1 data_queue_reg_2__6__2_ ( .D(n15855), .CK(clk), .Q(
        data_queue_2__6__2_), .QN(n1114) );
  DFF_X1 data_queue_reg_2__6__1_ ( .D(n15848), .CK(clk), .Q(
        data_queue_2__6__1_), .QN(n1115) );
  DFF_X1 data_queue_reg_2__6__0_ ( .D(n15841), .CK(clk), .Q(
        data_queue_2__6__0_), .QN(n1116) );
  DFF_X1 data_queue_reg_2__7__7_ ( .D(n15840), .CK(clk), .Q(
        data_queue_2__7__7_), .QN(n17248) );
  DFF_X1 data_queue_reg_2__7__6_ ( .D(n15837), .CK(clk), .Q(
        data_queue_2__7__6_), .QN(n17247) );
  DFF_X1 data_queue_reg_2__7__5_ ( .D(n15834), .CK(clk), .Q(
        data_queue_2__7__5_), .QN(n17246) );
  DFF_X1 data_queue_reg_2__7__4_ ( .D(n15831), .CK(clk), .Q(
        data_queue_2__7__4_), .QN(n17245) );
  DFF_X1 data_queue_reg_2__7__3_ ( .D(n15828), .CK(clk), .Q(
        data_queue_2__7__3_), .QN(n17244) );
  DFF_X1 data_queue_reg_2__7__2_ ( .D(n15825), .CK(clk), .Q(
        data_queue_2__7__2_), .QN(n17243) );
  DFF_X1 data_queue_reg_2__7__1_ ( .D(n15822), .CK(clk), .Q(
        data_queue_2__7__1_), .QN(n17242) );
  DFF_X1 data_queue_reg_2__7__0_ ( .D(n15819), .CK(clk), .Q(
        data_queue_2__7__0_), .QN(n17241) );
  DFF_X1 data_queue_reg_3__0__7_ ( .D(n15812), .CK(clk), .Q(
        data_queue_3__0__7_), .QN(n1117) );
  DFF_X1 data_queue_reg_3__0__6_ ( .D(n15807), .CK(clk), .Q(
        data_queue_3__0__6_), .QN(n1118) );
  DFF_X1 data_queue_reg_3__0__5_ ( .D(n15802), .CK(clk), .Q(
        data_queue_3__0__5_), .QN(n1119) );
  DFF_X1 data_queue_reg_3__0__4_ ( .D(n15797), .CK(clk), .Q(
        data_queue_3__0__4_), .QN(n1120) );
  DFF_X1 data_queue_reg_3__0__3_ ( .D(n15792), .CK(clk), .Q(
        data_queue_3__0__3_), .QN(n1121) );
  DFF_X1 data_queue_reg_3__0__2_ ( .D(n15787), .CK(clk), .Q(
        data_queue_3__0__2_), .QN(n1122) );
  DFF_X1 data_queue_reg_3__0__1_ ( .D(n15782), .CK(clk), .Q(
        data_queue_3__0__1_), .QN(n1123) );
  DFF_X1 data_queue_reg_3__0__0_ ( .D(n15777), .CK(clk), .Q(
        data_queue_3__0__0_), .QN(n1124) );
  DFF_X1 data_queue_reg_3__1__7_ ( .D(n15772), .CK(clk), .Q(
        data_queue_3__1__7_), .QN(n1125) );
  DFF_X1 data_queue_reg_3__1__6_ ( .D(n15767), .CK(clk), .Q(
        data_queue_3__1__6_), .QN(n1126) );
  DFF_X1 data_queue_reg_3__1__5_ ( .D(n15762), .CK(clk), .Q(
        data_queue_3__1__5_), .QN(n1127) );
  DFF_X1 data_queue_reg_3__1__4_ ( .D(n15757), .CK(clk), .Q(
        data_queue_3__1__4_), .QN(n1128) );
  DFF_X1 data_queue_reg_3__1__3_ ( .D(n15752), .CK(clk), .Q(
        data_queue_3__1__3_), .QN(n1129) );
  DFF_X1 data_queue_reg_3__1__2_ ( .D(n15747), .CK(clk), .Q(
        data_queue_3__1__2_), .QN(n1130) );
  DFF_X1 data_queue_reg_3__1__1_ ( .D(n15742), .CK(clk), .Q(
        data_queue_3__1__1_), .QN(n1131) );
  DFF_X1 data_queue_reg_3__1__0_ ( .D(n15737), .CK(clk), .Q(
        data_queue_3__1__0_), .QN(n1132) );
  DFF_X1 data_queue_reg_3__2__7_ ( .D(n15732), .CK(clk), .Q(
        data_queue_3__2__7_), .QN(n1133) );
  DFF_X1 data_queue_reg_3__2__6_ ( .D(n15727), .CK(clk), .Q(
        data_queue_3__2__6_), .QN(n1134) );
  DFF_X1 data_queue_reg_3__2__5_ ( .D(n15722), .CK(clk), .Q(
        data_queue_3__2__5_), .QN(n1135) );
  DFF_X1 data_queue_reg_3__2__4_ ( .D(n15717), .CK(clk), .Q(
        data_queue_3__2__4_), .QN(n1136) );
  DFF_X1 data_queue_reg_3__2__3_ ( .D(n15712), .CK(clk), .Q(
        data_queue_3__2__3_), .QN(n1137) );
  DFF_X1 data_queue_reg_3__2__2_ ( .D(n15707), .CK(clk), .Q(
        data_queue_3__2__2_), .QN(n1138) );
  DFF_X1 data_queue_reg_3__2__1_ ( .D(n15702), .CK(clk), .Q(
        data_queue_3__2__1_), .QN(n1139) );
  DFF_X1 data_queue_reg_3__2__0_ ( .D(n15697), .CK(clk), .Q(
        data_queue_3__2__0_), .QN(n1140) );
  DFF_X1 data_queue_reg_3__3__7_ ( .D(n15692), .CK(clk), .Q(
        data_queue_3__3__7_), .QN(n1141) );
  DFF_X1 data_queue_reg_3__3__6_ ( .D(n15687), .CK(clk), .Q(
        data_queue_3__3__6_), .QN(n1142) );
  DFF_X1 data_queue_reg_3__3__5_ ( .D(n15682), .CK(clk), .Q(
        data_queue_3__3__5_), .QN(n1143) );
  DFF_X1 data_queue_reg_3__3__4_ ( .D(n15677), .CK(clk), .Q(
        data_queue_3__3__4_), .QN(n1144) );
  DFF_X1 data_queue_reg_3__3__3_ ( .D(n15672), .CK(clk), .Q(
        data_queue_3__3__3_), .QN(n1145) );
  DFF_X1 data_queue_reg_3__3__2_ ( .D(n15667), .CK(clk), .Q(
        data_queue_3__3__2_), .QN(n1146) );
  DFF_X1 data_queue_reg_3__3__1_ ( .D(n15662), .CK(clk), .Q(
        data_queue_3__3__1_), .QN(n1147) );
  DFF_X1 data_queue_reg_3__3__0_ ( .D(n15657), .CK(clk), .Q(
        data_queue_3__3__0_), .QN(n1148) );
  DFF_X1 data_queue_reg_3__4__7_ ( .D(n15652), .CK(clk), .Q(
        data_queue_3__4__7_), .QN(n1149) );
  DFF_X1 data_queue_reg_3__4__6_ ( .D(n15647), .CK(clk), .Q(
        data_queue_3__4__6_), .QN(n1150) );
  DFF_X1 data_queue_reg_3__4__5_ ( .D(n15642), .CK(clk), .Q(
        data_queue_3__4__5_), .QN(n1151) );
  DFF_X1 data_queue_reg_3__4__4_ ( .D(n15637), .CK(clk), .Q(
        data_queue_3__4__4_), .QN(n1152) );
  DFF_X1 data_queue_reg_3__4__3_ ( .D(n15632), .CK(clk), .Q(
        data_queue_3__4__3_), .QN(n1153) );
  DFF_X1 data_queue_reg_3__4__2_ ( .D(n15627), .CK(clk), .Q(
        data_queue_3__4__2_), .QN(n1154) );
  DFF_X1 data_queue_reg_3__4__1_ ( .D(n15622), .CK(clk), .Q(
        data_queue_3__4__1_), .QN(n1155) );
  DFF_X1 data_queue_reg_3__4__0_ ( .D(n15617), .CK(clk), .Q(
        data_queue_3__4__0_), .QN(n1156) );
  DFF_X1 data_queue_reg_3__5__7_ ( .D(n15612), .CK(clk), .Q(
        data_queue_3__5__7_), .QN(n1157) );
  DFF_X1 data_queue_reg_3__5__6_ ( .D(n15607), .CK(clk), .Q(
        data_queue_3__5__6_), .QN(n1158) );
  DFF_X1 data_queue_reg_3__5__5_ ( .D(n15602), .CK(clk), .Q(
        data_queue_3__5__5_), .QN(n1159) );
  DFF_X1 data_queue_reg_3__5__4_ ( .D(n15597), .CK(clk), .Q(
        data_queue_3__5__4_), .QN(n1160) );
  DFF_X1 data_queue_reg_3__5__3_ ( .D(n15592), .CK(clk), .Q(
        data_queue_3__5__3_), .QN(n1161) );
  DFF_X1 data_queue_reg_3__5__2_ ( .D(n15587), .CK(clk), .Q(
        data_queue_3__5__2_), .QN(n1162) );
  DFF_X1 data_queue_reg_3__5__1_ ( .D(n15582), .CK(clk), .Q(
        data_queue_3__5__1_), .QN(n1163) );
  DFF_X1 data_queue_reg_3__5__0_ ( .D(n15577), .CK(clk), .Q(
        data_queue_3__5__0_), .QN(n1164) );
  DFF_X1 data_queue_reg_3__6__7_ ( .D(n15570), .CK(clk), .Q(
        data_queue_3__6__7_), .QN(n1165) );
  DFF_X1 data_queue_reg_3__6__6_ ( .D(n15563), .CK(clk), .Q(
        data_queue_3__6__6_), .QN(n1166) );
  DFF_X1 data_queue_reg_3__6__5_ ( .D(n15556), .CK(clk), .Q(
        data_queue_3__6__5_), .QN(n1167) );
  DFF_X1 data_queue_reg_3__6__4_ ( .D(n15549), .CK(clk), .Q(
        data_queue_3__6__4_), .QN(n1168) );
  DFF_X1 data_queue_reg_3__6__3_ ( .D(n15542), .CK(clk), .Q(
        data_queue_3__6__3_), .QN(n1169) );
  DFF_X1 data_queue_reg_3__6__2_ ( .D(n15535), .CK(clk), .Q(
        data_queue_3__6__2_), .QN(n1170) );
  DFF_X1 data_queue_reg_3__6__1_ ( .D(n15528), .CK(clk), .Q(
        data_queue_3__6__1_), .QN(n1171) );
  DFF_X1 data_queue_reg_3__6__0_ ( .D(n15521), .CK(clk), .Q(
        data_queue_3__6__0_), .QN(n1172) );
  DFF_X1 data_queue_reg_3__7__7_ ( .D(n15520), .CK(clk), .Q(
        data_queue_3__7__7_), .QN(n17240) );
  DFF_X1 data_queue_reg_3__7__6_ ( .D(n15517), .CK(clk), .Q(
        data_queue_3__7__6_), .QN(n17239) );
  DFF_X1 data_queue_reg_3__7__5_ ( .D(n15514), .CK(clk), .Q(
        data_queue_3__7__5_), .QN(n17238) );
  DFF_X1 data_queue_reg_3__7__4_ ( .D(n15511), .CK(clk), .Q(
        data_queue_3__7__4_), .QN(n17237) );
  DFF_X1 data_queue_reg_3__7__3_ ( .D(n15508), .CK(clk), .Q(
        data_queue_3__7__3_), .QN(n17236) );
  DFF_X1 data_queue_reg_3__7__2_ ( .D(n15505), .CK(clk), .Q(
        data_queue_3__7__2_), .QN(n17235) );
  DFF_X1 data_queue_reg_3__7__1_ ( .D(n15502), .CK(clk), .Q(
        data_queue_3__7__1_), .QN(n17234) );
  DFF_X1 data_queue_reg_3__7__0_ ( .D(n15499), .CK(clk), .Q(
        data_queue_3__7__0_), .QN(n17233) );
  DFF_X1 data_queue_reg_4__0__7_ ( .D(n15492), .CK(clk), .Q(
        data_queue_4__0__7_), .QN(n1173) );
  DFF_X1 data_queue_reg_4__0__6_ ( .D(n15487), .CK(clk), .Q(
        data_queue_4__0__6_), .QN(n1174) );
  DFF_X1 data_queue_reg_4__0__5_ ( .D(n15482), .CK(clk), .Q(
        data_queue_4__0__5_), .QN(n1175) );
  DFF_X1 data_queue_reg_4__0__4_ ( .D(n15477), .CK(clk), .Q(
        data_queue_4__0__4_), .QN(n1176) );
  DFF_X1 data_queue_reg_4__0__3_ ( .D(n15472), .CK(clk), .Q(
        data_queue_4__0__3_), .QN(n1177) );
  DFF_X1 data_queue_reg_4__0__2_ ( .D(n15467), .CK(clk), .Q(
        data_queue_4__0__2_), .QN(n1178) );
  DFF_X1 data_queue_reg_4__0__1_ ( .D(n15462), .CK(clk), .Q(
        data_queue_4__0__1_), .QN(n1179) );
  DFF_X1 data_queue_reg_4__0__0_ ( .D(n15457), .CK(clk), .Q(
        data_queue_4__0__0_), .QN(n1180) );
  DFF_X1 data_queue_reg_4__1__7_ ( .D(n15452), .CK(clk), .Q(
        data_queue_4__1__7_), .QN(n1181) );
  DFF_X1 data_queue_reg_4__1__6_ ( .D(n15447), .CK(clk), .Q(
        data_queue_4__1__6_), .QN(n1182) );
  DFF_X1 data_queue_reg_4__1__5_ ( .D(n15442), .CK(clk), .Q(
        data_queue_4__1__5_), .QN(n1183) );
  DFF_X1 data_queue_reg_4__1__4_ ( .D(n15437), .CK(clk), .Q(
        data_queue_4__1__4_), .QN(n1184) );
  DFF_X1 data_queue_reg_4__1__3_ ( .D(n15432), .CK(clk), .Q(
        data_queue_4__1__3_), .QN(n1185) );
  DFF_X1 data_queue_reg_4__1__2_ ( .D(n15427), .CK(clk), .Q(
        data_queue_4__1__2_), .QN(n1186) );
  DFF_X1 data_queue_reg_4__1__1_ ( .D(n15422), .CK(clk), .Q(
        data_queue_4__1__1_), .QN(n1187) );
  DFF_X1 data_queue_reg_4__1__0_ ( .D(n15417), .CK(clk), .Q(
        data_queue_4__1__0_), .QN(n1188) );
  DFF_X1 data_queue_reg_4__2__7_ ( .D(n15412), .CK(clk), .Q(
        data_queue_4__2__7_), .QN(n1189) );
  DFF_X1 data_queue_reg_4__2__6_ ( .D(n15407), .CK(clk), .Q(
        data_queue_4__2__6_), .QN(n1190) );
  DFF_X1 data_queue_reg_4__2__5_ ( .D(n15402), .CK(clk), .Q(
        data_queue_4__2__5_), .QN(n1191) );
  DFF_X1 data_queue_reg_4__2__4_ ( .D(n15397), .CK(clk), .Q(
        data_queue_4__2__4_), .QN(n1192) );
  DFF_X1 data_queue_reg_4__2__3_ ( .D(n15392), .CK(clk), .Q(
        data_queue_4__2__3_), .QN(n1193) );
  DFF_X1 data_queue_reg_4__2__2_ ( .D(n15387), .CK(clk), .Q(
        data_queue_4__2__2_), .QN(n1194) );
  DFF_X1 data_queue_reg_4__2__1_ ( .D(n15382), .CK(clk), .Q(
        data_queue_4__2__1_), .QN(n1195) );
  DFF_X1 data_queue_reg_4__2__0_ ( .D(n15377), .CK(clk), .Q(
        data_queue_4__2__0_), .QN(n1196) );
  DFF_X1 data_queue_reg_4__3__7_ ( .D(n15372), .CK(clk), .Q(
        data_queue_4__3__7_), .QN(n1197) );
  DFF_X1 data_queue_reg_4__3__6_ ( .D(n15367), .CK(clk), .Q(
        data_queue_4__3__6_), .QN(n1198) );
  DFF_X1 data_queue_reg_4__3__5_ ( .D(n15362), .CK(clk), .Q(
        data_queue_4__3__5_), .QN(n1199) );
  DFF_X1 data_queue_reg_4__3__4_ ( .D(n15357), .CK(clk), .Q(
        data_queue_4__3__4_), .QN(n1200) );
  DFF_X1 data_queue_reg_4__3__3_ ( .D(n15352), .CK(clk), .Q(
        data_queue_4__3__3_), .QN(n1201) );
  DFF_X1 data_queue_reg_4__3__2_ ( .D(n15347), .CK(clk), .Q(
        data_queue_4__3__2_), .QN(n1202) );
  DFF_X1 data_queue_reg_4__3__1_ ( .D(n15342), .CK(clk), .Q(
        data_queue_4__3__1_), .QN(n1203) );
  DFF_X1 data_queue_reg_4__3__0_ ( .D(n15337), .CK(clk), .Q(
        data_queue_4__3__0_), .QN(n1204) );
  DFF_X1 data_queue_reg_4__4__7_ ( .D(n15332), .CK(clk), .Q(
        data_queue_4__4__7_), .QN(n1205) );
  DFF_X1 data_queue_reg_4__4__6_ ( .D(n15327), .CK(clk), .Q(
        data_queue_4__4__6_), .QN(n1206) );
  DFF_X1 data_queue_reg_4__4__5_ ( .D(n15322), .CK(clk), .Q(
        data_queue_4__4__5_), .QN(n1207) );
  DFF_X1 data_queue_reg_4__4__4_ ( .D(n15317), .CK(clk), .Q(
        data_queue_4__4__4_), .QN(n1208) );
  DFF_X1 data_queue_reg_4__4__3_ ( .D(n15312), .CK(clk), .Q(
        data_queue_4__4__3_), .QN(n1209) );
  DFF_X1 data_queue_reg_4__4__2_ ( .D(n15307), .CK(clk), .Q(
        data_queue_4__4__2_), .QN(n1210) );
  DFF_X1 data_queue_reg_4__4__1_ ( .D(n15302), .CK(clk), .Q(
        data_queue_4__4__1_), .QN(n1211) );
  DFF_X1 data_queue_reg_4__4__0_ ( .D(n15297), .CK(clk), .Q(
        data_queue_4__4__0_), .QN(n1212) );
  DFF_X1 data_queue_reg_4__5__7_ ( .D(n15292), .CK(clk), .Q(
        data_queue_4__5__7_), .QN(n1213) );
  DFF_X1 data_queue_reg_4__5__6_ ( .D(n15287), .CK(clk), .Q(
        data_queue_4__5__6_), .QN(n1214) );
  DFF_X1 data_queue_reg_4__5__5_ ( .D(n15282), .CK(clk), .Q(
        data_queue_4__5__5_), .QN(n1215) );
  DFF_X1 data_queue_reg_4__5__4_ ( .D(n15277), .CK(clk), .Q(
        data_queue_4__5__4_), .QN(n1216) );
  DFF_X1 data_queue_reg_4__5__3_ ( .D(n15272), .CK(clk), .Q(
        data_queue_4__5__3_), .QN(n1217) );
  DFF_X1 data_queue_reg_4__5__2_ ( .D(n15267), .CK(clk), .Q(
        data_queue_4__5__2_), .QN(n1218) );
  DFF_X1 data_queue_reg_4__5__1_ ( .D(n15262), .CK(clk), .Q(
        data_queue_4__5__1_), .QN(n1219) );
  DFF_X1 data_queue_reg_4__5__0_ ( .D(n15257), .CK(clk), .Q(
        data_queue_4__5__0_), .QN(n1220) );
  DFF_X1 data_queue_reg_4__6__7_ ( .D(n15250), .CK(clk), .Q(
        data_queue_4__6__7_), .QN(n1221) );
  DFF_X1 data_queue_reg_4__6__6_ ( .D(n15243), .CK(clk), .Q(
        data_queue_4__6__6_), .QN(n1222) );
  DFF_X1 data_queue_reg_4__6__5_ ( .D(n15236), .CK(clk), .Q(
        data_queue_4__6__5_), .QN(n1223) );
  DFF_X1 data_queue_reg_4__6__4_ ( .D(n15229), .CK(clk), .Q(
        data_queue_4__6__4_), .QN(n1224) );
  DFF_X1 data_queue_reg_4__6__3_ ( .D(n15222), .CK(clk), .Q(
        data_queue_4__6__3_), .QN(n1225) );
  DFF_X1 data_queue_reg_4__6__2_ ( .D(n15215), .CK(clk), .Q(
        data_queue_4__6__2_), .QN(n1226) );
  DFF_X1 data_queue_reg_4__6__1_ ( .D(n15208), .CK(clk), .Q(
        data_queue_4__6__1_), .QN(n1227) );
  DFF_X1 data_queue_reg_4__6__0_ ( .D(n15201), .CK(clk), .Q(
        data_queue_4__6__0_), .QN(n1228) );
  DFF_X1 data_queue_reg_4__7__7_ ( .D(n15200), .CK(clk), .Q(
        data_queue_4__7__7_), .QN(n17232) );
  DFF_X1 data_queue_reg_4__7__6_ ( .D(n15197), .CK(clk), .Q(
        data_queue_4__7__6_), .QN(n17231) );
  DFF_X1 data_queue_reg_4__7__5_ ( .D(n15194), .CK(clk), .Q(
        data_queue_4__7__5_), .QN(n17230) );
  DFF_X1 data_queue_reg_4__7__4_ ( .D(n15191), .CK(clk), .Q(
        data_queue_4__7__4_), .QN(n17229) );
  DFF_X1 data_queue_reg_4__7__3_ ( .D(n15188), .CK(clk), .Q(
        data_queue_4__7__3_), .QN(n17228) );
  DFF_X1 data_queue_reg_4__7__2_ ( .D(n15185), .CK(clk), .Q(
        data_queue_4__7__2_), .QN(n17227) );
  DFF_X1 data_queue_reg_4__7__1_ ( .D(n15182), .CK(clk), .Q(
        data_queue_4__7__1_), .QN(n17226) );
  DFF_X1 data_queue_reg_4__7__0_ ( .D(n15179), .CK(clk), .Q(
        data_queue_4__7__0_), .QN(n17225) );
  DFF_X1 data_queue_reg_5__0__7_ ( .D(n15172), .CK(clk), .Q(
        data_queue_5__0__7_), .QN(n1229) );
  DFF_X1 data_queue_reg_5__0__6_ ( .D(n15167), .CK(clk), .Q(
        data_queue_5__0__6_), .QN(n1230) );
  DFF_X1 data_queue_reg_5__0__5_ ( .D(n15162), .CK(clk), .Q(
        data_queue_5__0__5_), .QN(n1231) );
  DFF_X1 data_queue_reg_5__0__4_ ( .D(n15157), .CK(clk), .Q(
        data_queue_5__0__4_), .QN(n1232) );
  DFF_X1 data_queue_reg_5__0__3_ ( .D(n15152), .CK(clk), .Q(
        data_queue_5__0__3_), .QN(n1233) );
  DFF_X1 data_queue_reg_5__0__2_ ( .D(n15147), .CK(clk), .Q(
        data_queue_5__0__2_), .QN(n1234) );
  DFF_X1 data_queue_reg_5__0__1_ ( .D(n15142), .CK(clk), .Q(
        data_queue_5__0__1_), .QN(n1235) );
  DFF_X1 data_queue_reg_5__0__0_ ( .D(n15137), .CK(clk), .Q(
        data_queue_5__0__0_), .QN(n1236) );
  DFF_X1 data_queue_reg_5__1__7_ ( .D(n15132), .CK(clk), .Q(
        data_queue_5__1__7_), .QN(n1237) );
  DFF_X1 data_queue_reg_5__1__6_ ( .D(n15127), .CK(clk), .Q(
        data_queue_5__1__6_), .QN(n1238) );
  DFF_X1 data_queue_reg_5__1__5_ ( .D(n15122), .CK(clk), .Q(
        data_queue_5__1__5_), .QN(n1239) );
  DFF_X1 data_queue_reg_5__1__4_ ( .D(n15117), .CK(clk), .Q(
        data_queue_5__1__4_), .QN(n1240) );
  DFF_X1 data_queue_reg_5__1__3_ ( .D(n15112), .CK(clk), .Q(
        data_queue_5__1__3_), .QN(n1241) );
  DFF_X1 data_queue_reg_5__1__2_ ( .D(n15107), .CK(clk), .Q(
        data_queue_5__1__2_), .QN(n1242) );
  DFF_X1 data_queue_reg_5__1__1_ ( .D(n15102), .CK(clk), .Q(
        data_queue_5__1__1_), .QN(n1243) );
  DFF_X1 data_queue_reg_5__1__0_ ( .D(n15097), .CK(clk), .Q(
        data_queue_5__1__0_), .QN(n1244) );
  DFF_X1 data_queue_reg_5__2__7_ ( .D(n15092), .CK(clk), .Q(
        data_queue_5__2__7_), .QN(n1245) );
  DFF_X1 data_queue_reg_5__2__6_ ( .D(n15087), .CK(clk), .Q(
        data_queue_5__2__6_), .QN(n1246) );
  DFF_X1 data_queue_reg_5__2__5_ ( .D(n15082), .CK(clk), .Q(
        data_queue_5__2__5_), .QN(n1247) );
  DFF_X1 data_queue_reg_5__2__4_ ( .D(n15077), .CK(clk), .Q(
        data_queue_5__2__4_), .QN(n1248) );
  DFF_X1 data_queue_reg_5__2__3_ ( .D(n15072), .CK(clk), .Q(
        data_queue_5__2__3_), .QN(n1249) );
  DFF_X1 data_queue_reg_5__2__2_ ( .D(n15067), .CK(clk), .Q(
        data_queue_5__2__2_), .QN(n1250) );
  DFF_X1 data_queue_reg_5__2__1_ ( .D(n15062), .CK(clk), .Q(
        data_queue_5__2__1_), .QN(n1251) );
  DFF_X1 data_queue_reg_5__2__0_ ( .D(n15057), .CK(clk), .Q(
        data_queue_5__2__0_), .QN(n1252) );
  DFF_X1 data_queue_reg_5__3__7_ ( .D(n15052), .CK(clk), .Q(
        data_queue_5__3__7_), .QN(n1253) );
  DFF_X1 data_queue_reg_5__3__6_ ( .D(n15047), .CK(clk), .Q(
        data_queue_5__3__6_), .QN(n1254) );
  DFF_X1 data_queue_reg_5__3__5_ ( .D(n15042), .CK(clk), .Q(
        data_queue_5__3__5_), .QN(n1255) );
  DFF_X1 data_queue_reg_5__3__4_ ( .D(n15037), .CK(clk), .Q(
        data_queue_5__3__4_), .QN(n1256) );
  DFF_X1 data_queue_reg_5__3__3_ ( .D(n15032), .CK(clk), .Q(
        data_queue_5__3__3_), .QN(n1257) );
  DFF_X1 data_queue_reg_5__3__2_ ( .D(n15027), .CK(clk), .Q(
        data_queue_5__3__2_), .QN(n1258) );
  DFF_X1 data_queue_reg_5__3__1_ ( .D(n15022), .CK(clk), .Q(
        data_queue_5__3__1_), .QN(n1259) );
  DFF_X1 data_queue_reg_5__3__0_ ( .D(n15017), .CK(clk), .Q(
        data_queue_5__3__0_), .QN(n1260) );
  DFF_X1 data_queue_reg_5__4__7_ ( .D(n15012), .CK(clk), .Q(
        data_queue_5__4__7_), .QN(n1261) );
  DFF_X1 data_queue_reg_5__4__6_ ( .D(n15007), .CK(clk), .Q(
        data_queue_5__4__6_), .QN(n1262) );
  DFF_X1 data_queue_reg_5__4__5_ ( .D(n15002), .CK(clk), .Q(
        data_queue_5__4__5_), .QN(n1263) );
  DFF_X1 data_queue_reg_5__4__4_ ( .D(n14997), .CK(clk), .Q(
        data_queue_5__4__4_), .QN(n1264) );
  DFF_X1 data_queue_reg_5__4__3_ ( .D(n14992), .CK(clk), .Q(
        data_queue_5__4__3_), .QN(n1265) );
  DFF_X1 data_queue_reg_5__4__2_ ( .D(n14987), .CK(clk), .Q(
        data_queue_5__4__2_), .QN(n1266) );
  DFF_X1 data_queue_reg_5__4__1_ ( .D(n14982), .CK(clk), .Q(
        data_queue_5__4__1_), .QN(n1267) );
  DFF_X1 data_queue_reg_5__4__0_ ( .D(n14977), .CK(clk), .Q(
        data_queue_5__4__0_), .QN(n1268) );
  DFF_X1 data_queue_reg_5__5__7_ ( .D(n14972), .CK(clk), .Q(
        data_queue_5__5__7_), .QN(n1269) );
  DFF_X1 data_queue_reg_5__5__6_ ( .D(n14967), .CK(clk), .Q(
        data_queue_5__5__6_), .QN(n1270) );
  DFF_X1 data_queue_reg_5__5__5_ ( .D(n14962), .CK(clk), .Q(
        data_queue_5__5__5_), .QN(n1271) );
  DFF_X1 data_queue_reg_5__5__4_ ( .D(n14957), .CK(clk), .Q(
        data_queue_5__5__4_), .QN(n1272) );
  DFF_X1 data_queue_reg_5__5__3_ ( .D(n14952), .CK(clk), .Q(
        data_queue_5__5__3_), .QN(n1273) );
  DFF_X1 data_queue_reg_5__5__2_ ( .D(n14947), .CK(clk), .Q(
        data_queue_5__5__2_), .QN(n1274) );
  DFF_X1 data_queue_reg_5__5__1_ ( .D(n14942), .CK(clk), .Q(
        data_queue_5__5__1_), .QN(n1275) );
  DFF_X1 data_queue_reg_5__5__0_ ( .D(n14937), .CK(clk), .Q(
        data_queue_5__5__0_), .QN(n1276) );
  DFF_X1 data_queue_reg_5__6__7_ ( .D(n14930), .CK(clk), .Q(
        data_queue_5__6__7_), .QN(n1277) );
  DFF_X1 data_queue_reg_5__6__6_ ( .D(n14923), .CK(clk), .Q(
        data_queue_5__6__6_), .QN(n1278) );
  DFF_X1 data_queue_reg_5__6__5_ ( .D(n14916), .CK(clk), .Q(
        data_queue_5__6__5_), .QN(n1279) );
  DFF_X1 data_queue_reg_5__6__4_ ( .D(n14909), .CK(clk), .Q(
        data_queue_5__6__4_), .QN(n1280) );
  DFF_X1 data_queue_reg_5__6__3_ ( .D(n14902), .CK(clk), .Q(
        data_queue_5__6__3_), .QN(n1281) );
  DFF_X1 data_queue_reg_5__6__2_ ( .D(n14895), .CK(clk), .Q(
        data_queue_5__6__2_), .QN(n1282) );
  DFF_X1 data_queue_reg_5__6__1_ ( .D(n14888), .CK(clk), .Q(
        data_queue_5__6__1_), .QN(n1283) );
  DFF_X1 data_queue_reg_5__6__0_ ( .D(n14881), .CK(clk), .Q(
        data_queue_5__6__0_), .QN(n1284) );
  DFF_X1 data_queue_reg_5__7__7_ ( .D(n14880), .CK(clk), .Q(
        data_queue_5__7__7_), .QN(n17224) );
  DFF_X1 data_queue_reg_5__7__6_ ( .D(n14877), .CK(clk), .Q(
        data_queue_5__7__6_), .QN(n17223) );
  DFF_X1 data_queue_reg_5__7__5_ ( .D(n14874), .CK(clk), .Q(
        data_queue_5__7__5_), .QN(n17222) );
  DFF_X1 data_queue_reg_5__7__4_ ( .D(n14871), .CK(clk), .Q(
        data_queue_5__7__4_), .QN(n17221) );
  DFF_X1 data_queue_reg_5__7__3_ ( .D(n14868), .CK(clk), .Q(
        data_queue_5__7__3_), .QN(n17220) );
  DFF_X1 data_queue_reg_5__7__2_ ( .D(n14865), .CK(clk), .Q(
        data_queue_5__7__2_), .QN(n17219) );
  DFF_X1 data_queue_reg_5__7__1_ ( .D(n14862), .CK(clk), .Q(
        data_queue_5__7__1_), .QN(n17218) );
  DFF_X1 data_queue_reg_5__7__0_ ( .D(n14859), .CK(clk), .Q(
        data_queue_5__7__0_), .QN(n17217) );
  DFF_X1 data_queue_reg_6__0__7_ ( .D(n14852), .CK(clk), .Q(
        data_queue_6__0__7_), .QN(n1285) );
  DFF_X1 data_queue_reg_6__0__6_ ( .D(n14847), .CK(clk), .Q(
        data_queue_6__0__6_), .QN(n1286) );
  DFF_X1 data_queue_reg_6__0__5_ ( .D(n14842), .CK(clk), .Q(
        data_queue_6__0__5_), .QN(n1287) );
  DFF_X1 data_queue_reg_6__0__4_ ( .D(n14837), .CK(clk), .Q(
        data_queue_6__0__4_), .QN(n1288) );
  DFF_X1 data_queue_reg_6__0__3_ ( .D(n14832), .CK(clk), .Q(
        data_queue_6__0__3_), .QN(n1289) );
  DFF_X1 data_queue_reg_6__0__2_ ( .D(n14827), .CK(clk), .Q(
        data_queue_6__0__2_), .QN(n1290) );
  DFF_X1 data_queue_reg_6__0__1_ ( .D(n14822), .CK(clk), .Q(
        data_queue_6__0__1_), .QN(n1291) );
  DFF_X1 data_queue_reg_6__0__0_ ( .D(n14817), .CK(clk), .Q(
        data_queue_6__0__0_), .QN(n1292) );
  DFF_X1 data_queue_reg_6__1__7_ ( .D(n14812), .CK(clk), .Q(
        data_queue_6__1__7_), .QN(n1293) );
  DFF_X1 data_queue_reg_6__1__6_ ( .D(n14807), .CK(clk), .Q(
        data_queue_6__1__6_), .QN(n1294) );
  DFF_X1 data_queue_reg_6__1__5_ ( .D(n14802), .CK(clk), .Q(
        data_queue_6__1__5_), .QN(n1295) );
  DFF_X1 data_queue_reg_6__1__4_ ( .D(n14797), .CK(clk), .Q(
        data_queue_6__1__4_), .QN(n1296) );
  DFF_X1 data_queue_reg_6__1__3_ ( .D(n14792), .CK(clk), .Q(
        data_queue_6__1__3_), .QN(n1297) );
  DFF_X1 data_queue_reg_6__1__2_ ( .D(n14787), .CK(clk), .Q(
        data_queue_6__1__2_), .QN(n1298) );
  DFF_X1 data_queue_reg_6__1__1_ ( .D(n14782), .CK(clk), .Q(
        data_queue_6__1__1_), .QN(n1299) );
  DFF_X1 data_queue_reg_6__1__0_ ( .D(n14777), .CK(clk), .Q(
        data_queue_6__1__0_), .QN(n1300) );
  DFF_X1 data_queue_reg_6__2__7_ ( .D(n14772), .CK(clk), .Q(
        data_queue_6__2__7_), .QN(n1301) );
  DFF_X1 data_queue_reg_6__2__6_ ( .D(n14767), .CK(clk), .Q(
        data_queue_6__2__6_), .QN(n1302) );
  DFF_X1 data_queue_reg_6__2__5_ ( .D(n14762), .CK(clk), .Q(
        data_queue_6__2__5_), .QN(n1303) );
  DFF_X1 data_queue_reg_6__2__4_ ( .D(n14757), .CK(clk), .Q(
        data_queue_6__2__4_), .QN(n1304) );
  DFF_X1 data_queue_reg_6__2__3_ ( .D(n14752), .CK(clk), .Q(
        data_queue_6__2__3_), .QN(n1305) );
  DFF_X1 data_queue_reg_6__2__2_ ( .D(n14747), .CK(clk), .Q(
        data_queue_6__2__2_), .QN(n1306) );
  DFF_X1 data_queue_reg_6__2__1_ ( .D(n14742), .CK(clk), .Q(
        data_queue_6__2__1_), .QN(n1307) );
  DFF_X1 data_queue_reg_6__2__0_ ( .D(n14737), .CK(clk), .Q(
        data_queue_6__2__0_), .QN(n1308) );
  DFF_X1 data_queue_reg_6__3__7_ ( .D(n14732), .CK(clk), .Q(
        data_queue_6__3__7_), .QN(n1309) );
  DFF_X1 data_queue_reg_6__3__6_ ( .D(n14727), .CK(clk), .Q(
        data_queue_6__3__6_), .QN(n1310) );
  DFF_X1 data_queue_reg_6__3__5_ ( .D(n14722), .CK(clk), .Q(
        data_queue_6__3__5_), .QN(n1311) );
  DFF_X1 data_queue_reg_6__3__4_ ( .D(n14717), .CK(clk), .Q(
        data_queue_6__3__4_), .QN(n1312) );
  DFF_X1 data_queue_reg_6__3__3_ ( .D(n14712), .CK(clk), .Q(
        data_queue_6__3__3_), .QN(n1313) );
  DFF_X1 data_queue_reg_6__3__2_ ( .D(n14707), .CK(clk), .Q(
        data_queue_6__3__2_), .QN(n1314) );
  DFF_X1 data_queue_reg_6__3__1_ ( .D(n14702), .CK(clk), .Q(
        data_queue_6__3__1_), .QN(n1315) );
  DFF_X1 data_queue_reg_6__3__0_ ( .D(n14697), .CK(clk), .Q(
        data_queue_6__3__0_), .QN(n1316) );
  DFF_X1 data_queue_reg_6__4__7_ ( .D(n14692), .CK(clk), .Q(
        data_queue_6__4__7_), .QN(n1317) );
  DFF_X1 data_queue_reg_6__4__6_ ( .D(n14687), .CK(clk), .Q(
        data_queue_6__4__6_), .QN(n1318) );
  DFF_X1 data_queue_reg_6__4__5_ ( .D(n14682), .CK(clk), .Q(
        data_queue_6__4__5_), .QN(n1319) );
  DFF_X1 data_queue_reg_6__4__4_ ( .D(n14677), .CK(clk), .Q(
        data_queue_6__4__4_), .QN(n1320) );
  DFF_X1 data_queue_reg_6__4__3_ ( .D(n14672), .CK(clk), .Q(
        data_queue_6__4__3_), .QN(n1321) );
  DFF_X1 data_queue_reg_6__4__2_ ( .D(n14667), .CK(clk), .Q(
        data_queue_6__4__2_), .QN(n1322) );
  DFF_X1 data_queue_reg_6__4__1_ ( .D(n14662), .CK(clk), .Q(
        data_queue_6__4__1_), .QN(n1323) );
  DFF_X1 data_queue_reg_6__4__0_ ( .D(n14657), .CK(clk), .Q(
        data_queue_6__4__0_), .QN(n1324) );
  DFF_X1 data_queue_reg_6__5__7_ ( .D(n14652), .CK(clk), .Q(
        data_queue_6__5__7_), .QN(n1325) );
  DFF_X1 data_queue_reg_6__5__6_ ( .D(n14647), .CK(clk), .Q(
        data_queue_6__5__6_), .QN(n1326) );
  DFF_X1 data_queue_reg_6__5__5_ ( .D(n14642), .CK(clk), .Q(
        data_queue_6__5__5_), .QN(n1327) );
  DFF_X1 data_queue_reg_6__5__4_ ( .D(n14637), .CK(clk), .Q(
        data_queue_6__5__4_), .QN(n1328) );
  DFF_X1 data_queue_reg_6__5__3_ ( .D(n14632), .CK(clk), .Q(
        data_queue_6__5__3_), .QN(n1329) );
  DFF_X1 data_queue_reg_6__5__2_ ( .D(n14627), .CK(clk), .Q(
        data_queue_6__5__2_), .QN(n1330) );
  DFF_X1 data_queue_reg_6__5__1_ ( .D(n14622), .CK(clk), .Q(
        data_queue_6__5__1_), .QN(n1331) );
  DFF_X1 data_queue_reg_6__5__0_ ( .D(n14617), .CK(clk), .Q(
        data_queue_6__5__0_), .QN(n1332) );
  DFF_X1 data_queue_reg_6__6__7_ ( .D(n14610), .CK(clk), .Q(
        data_queue_6__6__7_), .QN(n1333) );
  DFF_X1 data_queue_reg_6__6__6_ ( .D(n14603), .CK(clk), .Q(
        data_queue_6__6__6_), .QN(n1334) );
  DFF_X1 data_queue_reg_6__6__5_ ( .D(n14596), .CK(clk), .Q(
        data_queue_6__6__5_), .QN(n1335) );
  DFF_X1 data_queue_reg_6__6__4_ ( .D(n14589), .CK(clk), .Q(
        data_queue_6__6__4_), .QN(n1336) );
  DFF_X1 data_queue_reg_6__6__3_ ( .D(n14582), .CK(clk), .Q(
        data_queue_6__6__3_), .QN(n1337) );
  DFF_X1 data_queue_reg_6__6__2_ ( .D(n14575), .CK(clk), .Q(
        data_queue_6__6__2_), .QN(n1338) );
  DFF_X1 data_queue_reg_6__6__1_ ( .D(n14568), .CK(clk), .Q(
        data_queue_6__6__1_), .QN(n1339) );
  DFF_X1 data_queue_reg_6__6__0_ ( .D(n14561), .CK(clk), .Q(
        data_queue_6__6__0_), .QN(n1340) );
  DFF_X1 data_queue_reg_6__7__7_ ( .D(n14560), .CK(clk), .Q(
        data_queue_6__7__7_), .QN(n17216) );
  DFF_X1 data_queue_reg_6__7__6_ ( .D(n14557), .CK(clk), .Q(
        data_queue_6__7__6_), .QN(n17215) );
  DFF_X1 data_queue_reg_6__7__5_ ( .D(n14554), .CK(clk), .Q(
        data_queue_6__7__5_), .QN(n17214) );
  DFF_X1 data_queue_reg_6__7__4_ ( .D(n14551), .CK(clk), .Q(
        data_queue_6__7__4_), .QN(n17213) );
  DFF_X1 data_queue_reg_6__7__3_ ( .D(n14548), .CK(clk), .Q(
        data_queue_6__7__3_), .QN(n17212) );
  DFF_X1 data_queue_reg_6__7__2_ ( .D(n14545), .CK(clk), .Q(
        data_queue_6__7__2_), .QN(n17211) );
  DFF_X1 data_queue_reg_6__7__1_ ( .D(n14542), .CK(clk), .Q(
        data_queue_6__7__1_), .QN(n17210) );
  DFF_X1 data_queue_reg_6__7__0_ ( .D(n14539), .CK(clk), .Q(
        data_queue_6__7__0_), .QN(n17209) );
  DFF_X1 data_queue_reg_7__0__7_ ( .D(n14532), .CK(clk), .Q(
        data_queue_7__0__7_), .QN(n1341) );
  DFF_X1 data_queue_reg_7__0__6_ ( .D(n14527), .CK(clk), .Q(
        data_queue_7__0__6_), .QN(n1342) );
  DFF_X1 data_queue_reg_7__0__5_ ( .D(n14522), .CK(clk), .Q(
        data_queue_7__0__5_), .QN(n1343) );
  DFF_X1 data_queue_reg_7__0__4_ ( .D(n14517), .CK(clk), .Q(
        data_queue_7__0__4_), .QN(n1344) );
  DFF_X1 data_queue_reg_7__0__3_ ( .D(n14512), .CK(clk), .Q(
        data_queue_7__0__3_), .QN(n1345) );
  DFF_X1 data_queue_reg_7__0__2_ ( .D(n14507), .CK(clk), .Q(
        data_queue_7__0__2_), .QN(n1346) );
  DFF_X1 data_queue_reg_7__0__1_ ( .D(n14502), .CK(clk), .Q(
        data_queue_7__0__1_), .QN(n1347) );
  DFF_X1 data_queue_reg_7__0__0_ ( .D(n14497), .CK(clk), .Q(
        data_queue_7__0__0_), .QN(n1348) );
  DFF_X1 data_queue_reg_7__1__7_ ( .D(n14492), .CK(clk), .Q(
        data_queue_7__1__7_), .QN(n1349) );
  DFF_X1 data_queue_reg_7__1__6_ ( .D(n14487), .CK(clk), .Q(
        data_queue_7__1__6_), .QN(n1350) );
  DFF_X1 data_queue_reg_7__1__5_ ( .D(n14482), .CK(clk), .Q(
        data_queue_7__1__5_), .QN(n1351) );
  DFF_X1 data_queue_reg_7__1__4_ ( .D(n14477), .CK(clk), .Q(
        data_queue_7__1__4_), .QN(n1352) );
  DFF_X1 data_queue_reg_7__1__3_ ( .D(n14472), .CK(clk), .Q(
        data_queue_7__1__3_), .QN(n1353) );
  DFF_X1 data_queue_reg_7__1__2_ ( .D(n14467), .CK(clk), .Q(
        data_queue_7__1__2_), .QN(n1354) );
  DFF_X1 data_queue_reg_7__1__1_ ( .D(n14462), .CK(clk), .Q(
        data_queue_7__1__1_), .QN(n1355) );
  DFF_X1 data_queue_reg_7__1__0_ ( .D(n14457), .CK(clk), .Q(
        data_queue_7__1__0_), .QN(n1356) );
  DFF_X1 data_queue_reg_7__2__7_ ( .D(n14452), .CK(clk), .Q(
        data_queue_7__2__7_), .QN(n1357) );
  DFF_X1 data_queue_reg_7__2__6_ ( .D(n14447), .CK(clk), .Q(
        data_queue_7__2__6_), .QN(n1358) );
  DFF_X1 data_queue_reg_7__2__5_ ( .D(n14442), .CK(clk), .Q(
        data_queue_7__2__5_), .QN(n1359) );
  DFF_X1 data_queue_reg_7__2__4_ ( .D(n14437), .CK(clk), .Q(
        data_queue_7__2__4_), .QN(n1360) );
  DFF_X1 data_queue_reg_7__2__3_ ( .D(n14432), .CK(clk), .Q(
        data_queue_7__2__3_), .QN(n1361) );
  DFF_X1 data_queue_reg_7__2__2_ ( .D(n14427), .CK(clk), .Q(
        data_queue_7__2__2_), .QN(n1362) );
  DFF_X1 data_queue_reg_7__2__1_ ( .D(n14422), .CK(clk), .Q(
        data_queue_7__2__1_), .QN(n1363) );
  DFF_X1 data_queue_reg_7__2__0_ ( .D(n14417), .CK(clk), .Q(
        data_queue_7__2__0_), .QN(n1364) );
  DFF_X1 data_queue_reg_7__3__7_ ( .D(n14412), .CK(clk), .Q(
        data_queue_7__3__7_), .QN(n1365) );
  DFF_X1 data_queue_reg_7__3__6_ ( .D(n14407), .CK(clk), .Q(
        data_queue_7__3__6_), .QN(n1366) );
  DFF_X1 data_queue_reg_7__3__5_ ( .D(n14402), .CK(clk), .Q(
        data_queue_7__3__5_), .QN(n1367) );
  DFF_X1 data_queue_reg_7__3__4_ ( .D(n14397), .CK(clk), .Q(
        data_queue_7__3__4_), .QN(n1368) );
  DFF_X1 data_queue_reg_7__3__3_ ( .D(n14392), .CK(clk), .Q(
        data_queue_7__3__3_), .QN(n1369) );
  DFF_X1 data_queue_reg_7__3__2_ ( .D(n14387), .CK(clk), .Q(
        data_queue_7__3__2_), .QN(n1370) );
  DFF_X1 data_queue_reg_7__3__1_ ( .D(n14382), .CK(clk), .Q(
        data_queue_7__3__1_), .QN(n1371) );
  DFF_X1 data_queue_reg_7__3__0_ ( .D(n14377), .CK(clk), .Q(
        data_queue_7__3__0_), .QN(n1372) );
  DFF_X1 data_queue_reg_7__4__7_ ( .D(n14372), .CK(clk), .Q(
        data_queue_7__4__7_), .QN(n1373) );
  DFF_X1 data_queue_reg_7__4__6_ ( .D(n14367), .CK(clk), .Q(
        data_queue_7__4__6_), .QN(n1374) );
  DFF_X1 data_queue_reg_7__4__5_ ( .D(n14362), .CK(clk), .Q(
        data_queue_7__4__5_), .QN(n1375) );
  DFF_X1 data_queue_reg_7__4__4_ ( .D(n14357), .CK(clk), .Q(
        data_queue_7__4__4_), .QN(n1376) );
  DFF_X1 data_queue_reg_7__4__3_ ( .D(n14352), .CK(clk), .Q(
        data_queue_7__4__3_), .QN(n1377) );
  DFF_X1 data_queue_reg_7__4__2_ ( .D(n14347), .CK(clk), .Q(
        data_queue_7__4__2_), .QN(n1378) );
  DFF_X1 data_queue_reg_7__4__1_ ( .D(n14342), .CK(clk), .Q(
        data_queue_7__4__1_), .QN(n1379) );
  DFF_X1 data_queue_reg_7__4__0_ ( .D(n14337), .CK(clk), .Q(
        data_queue_7__4__0_), .QN(n1380) );
  DFF_X1 data_queue_reg_7__5__7_ ( .D(n14332), .CK(clk), .Q(
        data_queue_7__5__7_), .QN(n1381) );
  DFF_X1 data_queue_reg_7__5__6_ ( .D(n14327), .CK(clk), .Q(
        data_queue_7__5__6_), .QN(n1382) );
  DFF_X1 data_queue_reg_7__5__5_ ( .D(n14322), .CK(clk), .Q(
        data_queue_7__5__5_), .QN(n1383) );
  DFF_X1 data_queue_reg_7__5__4_ ( .D(n14317), .CK(clk), .Q(
        data_queue_7__5__4_), .QN(n1384) );
  DFF_X1 data_queue_reg_7__5__3_ ( .D(n14312), .CK(clk), .Q(
        data_queue_7__5__3_), .QN(n1385) );
  DFF_X1 data_queue_reg_7__5__2_ ( .D(n14307), .CK(clk), .Q(
        data_queue_7__5__2_), .QN(n1386) );
  DFF_X1 data_queue_reg_7__5__1_ ( .D(n14302), .CK(clk), .Q(
        data_queue_7__5__1_), .QN(n1387) );
  DFF_X1 data_queue_reg_7__5__0_ ( .D(n14297), .CK(clk), .Q(
        data_queue_7__5__0_), .QN(n1388) );
  DFF_X1 data_queue_reg_7__6__7_ ( .D(n14290), .CK(clk), .Q(
        data_queue_7__6__7_), .QN(n1389) );
  DFF_X1 data_queue_reg_7__6__6_ ( .D(n14283), .CK(clk), .Q(
        data_queue_7__6__6_), .QN(n1390) );
  DFF_X1 data_queue_reg_7__6__5_ ( .D(n14276), .CK(clk), .Q(
        data_queue_7__6__5_), .QN(n1391) );
  DFF_X1 data_queue_reg_7__6__4_ ( .D(n14269), .CK(clk), .Q(
        data_queue_7__6__4_), .QN(n1392) );
  DFF_X1 data_queue_reg_7__6__3_ ( .D(n14262), .CK(clk), .Q(
        data_queue_7__6__3_), .QN(n1393) );
  DFF_X1 data_queue_reg_7__6__2_ ( .D(n14255), .CK(clk), .Q(
        data_queue_7__6__2_), .QN(n1394) );
  DFF_X1 data_queue_reg_7__6__1_ ( .D(n14248), .CK(clk), .Q(
        data_queue_7__6__1_), .QN(n1395) );
  DFF_X1 data_queue_reg_7__6__0_ ( .D(n14241), .CK(clk), .Q(
        data_queue_7__6__0_), .QN(n1396) );
  DFF_X1 data_queue_reg_7__7__7_ ( .D(n14240), .CK(clk), .Q(
        data_queue_7__7__7_), .QN(n17208) );
  DFF_X1 data_queue_reg_7__7__6_ ( .D(n14237), .CK(clk), .Q(
        data_queue_7__7__6_), .QN(n17207) );
  DFF_X1 data_queue_reg_7__7__5_ ( .D(n14234), .CK(clk), .Q(
        data_queue_7__7__5_), .QN(n17206) );
  DFF_X1 data_queue_reg_7__7__4_ ( .D(n14231), .CK(clk), .Q(
        data_queue_7__7__4_), .QN(n17205) );
  DFF_X1 data_queue_reg_7__7__3_ ( .D(n14228), .CK(clk), .Q(
        data_queue_7__7__3_), .QN(n17204) );
  DFF_X1 data_queue_reg_7__7__2_ ( .D(n14225), .CK(clk), .Q(
        data_queue_7__7__2_), .QN(n17203) );
  DFF_X1 data_queue_reg_7__7__1_ ( .D(n14222), .CK(clk), .Q(
        data_queue_7__7__1_), .QN(n17202) );
  DFF_X1 data_queue_reg_7__7__0_ ( .D(n14219), .CK(clk), .Q(
        data_queue_7__7__0_), .QN(n17201) );
  DFF_X1 weight_queue_reg_0__0__7_ ( .D(n14212), .CK(clk), .Q(
        weight_queue_0__0__7_), .QN(n1397) );
  DFF_X1 weight_queue_reg_0__0__6_ ( .D(n14207), .CK(clk), .Q(
        weight_queue_0__0__6_), .QN(n1398) );
  DFF_X1 weight_queue_reg_0__0__5_ ( .D(n14202), .CK(clk), .Q(
        weight_queue_0__0__5_), .QN(n1399) );
  DFF_X1 weight_queue_reg_0__0__4_ ( .D(n14197), .CK(clk), .Q(
        weight_queue_0__0__4_), .QN(n1400) );
  DFF_X1 weight_queue_reg_0__0__3_ ( .D(n14192), .CK(clk), .Q(
        weight_queue_0__0__3_), .QN(n1401) );
  DFF_X1 weight_queue_reg_0__0__2_ ( .D(n14187), .CK(clk), .Q(
        weight_queue_0__0__2_), .QN(n1402) );
  DFF_X1 weight_queue_reg_0__0__1_ ( .D(n14182), .CK(clk), .Q(
        weight_queue_0__0__1_), .QN(n1403) );
  DFF_X1 weight_queue_reg_0__0__0_ ( .D(n14177), .CK(clk), .Q(
        weight_queue_0__0__0_), .QN(n1404) );
  DFF_X1 weight_queue_reg_0__1__7_ ( .D(n14172), .CK(clk), .Q(
        weight_queue_0__1__7_), .QN(n1405) );
  DFF_X1 weight_queue_reg_0__1__6_ ( .D(n14167), .CK(clk), .Q(
        weight_queue_0__1__6_), .QN(n1406) );
  DFF_X1 weight_queue_reg_0__1__5_ ( .D(n14162), .CK(clk), .Q(
        weight_queue_0__1__5_), .QN(n1407) );
  DFF_X1 weight_queue_reg_0__1__4_ ( .D(n14157), .CK(clk), .Q(
        weight_queue_0__1__4_), .QN(n1408) );
  DFF_X1 weight_queue_reg_0__1__3_ ( .D(n14152), .CK(clk), .Q(
        weight_queue_0__1__3_), .QN(n1409) );
  DFF_X1 weight_queue_reg_0__1__2_ ( .D(n14147), .CK(clk), .Q(
        weight_queue_0__1__2_), .QN(n1410) );
  DFF_X1 weight_queue_reg_0__1__1_ ( .D(n14142), .CK(clk), .Q(
        weight_queue_0__1__1_), .QN(n1411) );
  DFF_X1 weight_queue_reg_0__1__0_ ( .D(n14137), .CK(clk), .Q(
        weight_queue_0__1__0_), .QN(n1412) );
  DFF_X1 weight_queue_reg_0__2__7_ ( .D(n14132), .CK(clk), .Q(
        weight_queue_0__2__7_), .QN(n1413) );
  DFF_X1 weight_queue_reg_0__2__6_ ( .D(n14127), .CK(clk), .Q(
        weight_queue_0__2__6_), .QN(n1414) );
  DFF_X1 weight_queue_reg_0__2__5_ ( .D(n14122), .CK(clk), .Q(
        weight_queue_0__2__5_), .QN(n1415) );
  DFF_X1 weight_queue_reg_0__2__4_ ( .D(n14117), .CK(clk), .Q(
        weight_queue_0__2__4_), .QN(n1416) );
  DFF_X1 weight_queue_reg_0__2__3_ ( .D(n14112), .CK(clk), .Q(
        weight_queue_0__2__3_), .QN(n1417) );
  DFF_X1 weight_queue_reg_0__2__2_ ( .D(n14107), .CK(clk), .Q(
        weight_queue_0__2__2_), .QN(n1418) );
  DFF_X1 weight_queue_reg_0__2__1_ ( .D(n14102), .CK(clk), .Q(
        weight_queue_0__2__1_), .QN(n1419) );
  DFF_X1 weight_queue_reg_0__2__0_ ( .D(n14097), .CK(clk), .Q(
        weight_queue_0__2__0_), .QN(n1420) );
  DFF_X1 weight_queue_reg_0__3__7_ ( .D(n14092), .CK(clk), .Q(
        weight_queue_0__3__7_), .QN(n1421) );
  DFF_X1 weight_queue_reg_0__3__6_ ( .D(n14087), .CK(clk), .Q(
        weight_queue_0__3__6_), .QN(n1422) );
  DFF_X1 weight_queue_reg_0__3__5_ ( .D(n14082), .CK(clk), .Q(
        weight_queue_0__3__5_), .QN(n1423) );
  DFF_X1 weight_queue_reg_0__3__4_ ( .D(n14077), .CK(clk), .Q(
        weight_queue_0__3__4_), .QN(n1424) );
  DFF_X1 weight_queue_reg_0__3__3_ ( .D(n14072), .CK(clk), .Q(
        weight_queue_0__3__3_), .QN(n1425) );
  DFF_X1 weight_queue_reg_0__3__2_ ( .D(n14067), .CK(clk), .Q(
        weight_queue_0__3__2_), .QN(n1426) );
  DFF_X1 weight_queue_reg_0__3__1_ ( .D(n14062), .CK(clk), .Q(
        weight_queue_0__3__1_), .QN(n1427) );
  DFF_X1 weight_queue_reg_0__3__0_ ( .D(n14057), .CK(clk), .Q(
        weight_queue_0__3__0_), .QN(n1428) );
  DFF_X1 weight_queue_reg_0__4__7_ ( .D(n14052), .CK(clk), .Q(
        weight_queue_0__4__7_), .QN(n1429) );
  DFF_X1 weight_queue_reg_0__4__6_ ( .D(n14047), .CK(clk), .Q(
        weight_queue_0__4__6_), .QN(n1430) );
  DFF_X1 weight_queue_reg_0__4__5_ ( .D(n14042), .CK(clk), .Q(
        weight_queue_0__4__5_), .QN(n1431) );
  DFF_X1 weight_queue_reg_0__4__4_ ( .D(n14037), .CK(clk), .Q(
        weight_queue_0__4__4_), .QN(n1432) );
  DFF_X1 weight_queue_reg_0__4__3_ ( .D(n14032), .CK(clk), .Q(
        weight_queue_0__4__3_), .QN(n1433) );
  DFF_X1 weight_queue_reg_0__4__2_ ( .D(n14027), .CK(clk), .Q(
        weight_queue_0__4__2_), .QN(n1434) );
  DFF_X1 weight_queue_reg_0__4__1_ ( .D(n14022), .CK(clk), .Q(
        weight_queue_0__4__1_), .QN(n1435) );
  DFF_X1 weight_queue_reg_0__4__0_ ( .D(n14017), .CK(clk), .Q(
        weight_queue_0__4__0_), .QN(n1436) );
  DFF_X1 weight_queue_reg_0__5__7_ ( .D(n14012), .CK(clk), .Q(
        weight_queue_0__5__7_), .QN(n1437) );
  DFF_X1 weight_queue_reg_0__5__6_ ( .D(n14007), .CK(clk), .Q(
        weight_queue_0__5__6_), .QN(n1438) );
  DFF_X1 weight_queue_reg_0__5__5_ ( .D(n14002), .CK(clk), .Q(
        weight_queue_0__5__5_), .QN(n1439) );
  DFF_X1 weight_queue_reg_0__5__4_ ( .D(n13997), .CK(clk), .Q(
        weight_queue_0__5__4_), .QN(n1440) );
  DFF_X1 weight_queue_reg_0__5__3_ ( .D(n13992), .CK(clk), .Q(
        weight_queue_0__5__3_), .QN(n1441) );
  DFF_X1 weight_queue_reg_0__5__2_ ( .D(n13987), .CK(clk), .Q(
        weight_queue_0__5__2_), .QN(n1442) );
  DFF_X1 weight_queue_reg_0__5__1_ ( .D(n13982), .CK(clk), .Q(
        weight_queue_0__5__1_), .QN(n1443) );
  DFF_X1 weight_queue_reg_0__5__0_ ( .D(n13977), .CK(clk), .Q(
        weight_queue_0__5__0_), .QN(n1444) );
  DFF_X1 weight_queue_reg_0__6__7_ ( .D(n13972), .CK(clk), .Q(
        weight_queue_0__6__7_), .QN(n1445) );
  DFF_X1 weight_queue_reg_0__6__6_ ( .D(n13967), .CK(clk), .Q(
        weight_queue_0__6__6_), .QN(n1446) );
  DFF_X1 weight_queue_reg_0__6__5_ ( .D(n13962), .CK(clk), .Q(
        weight_queue_0__6__5_), .QN(n1447) );
  DFF_X1 weight_queue_reg_0__6__4_ ( .D(n13957), .CK(clk), .Q(
        weight_queue_0__6__4_), .QN(n1448) );
  DFF_X1 weight_queue_reg_0__6__3_ ( .D(n13952), .CK(clk), .Q(
        weight_queue_0__6__3_), .QN(n1449) );
  DFF_X1 weight_queue_reg_0__6__2_ ( .D(n13947), .CK(clk), .Q(
        weight_queue_0__6__2_), .QN(n1450) );
  DFF_X1 weight_queue_reg_0__6__1_ ( .D(n13942), .CK(clk), .Q(
        weight_queue_0__6__1_), .QN(n1451) );
  DFF_X1 weight_queue_reg_0__6__0_ ( .D(n13937), .CK(clk), .Q(
        weight_queue_0__6__0_), .QN(n1452) );
  DFF_X1 weight_queue_reg_0__7__7_ ( .D(n13932), .CK(clk), .Q(
        weight_queue_0__7__7_), .QN(n1453) );
  DFF_X1 weight_queue_reg_0__7__6_ ( .D(n13927), .CK(clk), .Q(
        weight_queue_0__7__6_), .QN(n1454) );
  DFF_X1 weight_queue_reg_0__7__5_ ( .D(n13922), .CK(clk), .Q(
        weight_queue_0__7__5_), .QN(n1455) );
  DFF_X1 weight_queue_reg_0__7__4_ ( .D(n13917), .CK(clk), .Q(
        weight_queue_0__7__4_), .QN(n1456) );
  DFF_X1 weight_queue_reg_0__7__3_ ( .D(n13912), .CK(clk), .Q(
        weight_queue_0__7__3_), .QN(n1457) );
  DFF_X1 weight_queue_reg_0__7__2_ ( .D(n13907), .CK(clk), .Q(
        weight_queue_0__7__2_), .QN(n1458) );
  DFF_X1 weight_queue_reg_0__7__1_ ( .D(n13902), .CK(clk), .Q(
        weight_queue_0__7__1_), .QN(n1459) );
  DFF_X1 weight_queue_reg_0__7__0_ ( .D(n13897), .CK(clk), .Q(
        weight_queue_0__7__0_), .QN(n1460) );
  DFF_X1 weight_queue_reg_1__0__7_ ( .D(n13892), .CK(clk), .Q(
        weight_queue_1__0__7_), .QN(n1461) );
  DFF_X1 weight_queue_reg_1__0__6_ ( .D(n13887), .CK(clk), .Q(
        weight_queue_1__0__6_), .QN(n1462) );
  DFF_X1 weight_queue_reg_1__0__5_ ( .D(n13882), .CK(clk), .Q(
        weight_queue_1__0__5_), .QN(n1463) );
  DFF_X1 weight_queue_reg_1__0__4_ ( .D(n13877), .CK(clk), .Q(
        weight_queue_1__0__4_), .QN(n1464) );
  DFF_X1 weight_queue_reg_1__0__3_ ( .D(n13872), .CK(clk), .Q(
        weight_queue_1__0__3_), .QN(n1465) );
  DFF_X1 weight_queue_reg_1__0__2_ ( .D(n13867), .CK(clk), .Q(
        weight_queue_1__0__2_), .QN(n1466) );
  DFF_X1 weight_queue_reg_1__0__1_ ( .D(n13862), .CK(clk), .Q(
        weight_queue_1__0__1_), .QN(n1467) );
  DFF_X1 weight_queue_reg_1__0__0_ ( .D(n13857), .CK(clk), .Q(
        weight_queue_1__0__0_), .QN(n1468) );
  DFF_X1 weight_queue_reg_1__1__7_ ( .D(n13852), .CK(clk), .Q(
        weight_queue_1__1__7_), .QN(n1469) );
  DFF_X1 weight_queue_reg_1__1__6_ ( .D(n13847), .CK(clk), .Q(
        weight_queue_1__1__6_), .QN(n1470) );
  DFF_X1 weight_queue_reg_1__1__5_ ( .D(n13842), .CK(clk), .Q(
        weight_queue_1__1__5_), .QN(n1471) );
  DFF_X1 weight_queue_reg_1__1__4_ ( .D(n13837), .CK(clk), .Q(
        weight_queue_1__1__4_), .QN(n1472) );
  DFF_X1 weight_queue_reg_1__1__3_ ( .D(n13832), .CK(clk), .Q(
        weight_queue_1__1__3_), .QN(n1473) );
  DFF_X1 weight_queue_reg_1__1__2_ ( .D(n13827), .CK(clk), .Q(
        weight_queue_1__1__2_), .QN(n1474) );
  DFF_X1 weight_queue_reg_1__1__1_ ( .D(n13822), .CK(clk), .Q(
        weight_queue_1__1__1_), .QN(n1475) );
  DFF_X1 weight_queue_reg_1__1__0_ ( .D(n13817), .CK(clk), .Q(
        weight_queue_1__1__0_), .QN(n1476) );
  DFF_X1 weight_queue_reg_1__2__7_ ( .D(n13812), .CK(clk), .Q(
        weight_queue_1__2__7_), .QN(n1477) );
  DFF_X1 weight_queue_reg_1__2__6_ ( .D(n13807), .CK(clk), .Q(
        weight_queue_1__2__6_), .QN(n1478) );
  DFF_X1 weight_queue_reg_1__2__5_ ( .D(n13802), .CK(clk), .Q(
        weight_queue_1__2__5_), .QN(n1479) );
  DFF_X1 weight_queue_reg_1__2__4_ ( .D(n13797), .CK(clk), .Q(
        weight_queue_1__2__4_), .QN(n1480) );
  DFF_X1 weight_queue_reg_1__2__3_ ( .D(n13792), .CK(clk), .Q(
        weight_queue_1__2__3_), .QN(n1481) );
  DFF_X1 weight_queue_reg_1__2__2_ ( .D(n13787), .CK(clk), .Q(
        weight_queue_1__2__2_), .QN(n1482) );
  DFF_X1 weight_queue_reg_1__2__1_ ( .D(n13782), .CK(clk), .Q(
        weight_queue_1__2__1_), .QN(n1483) );
  DFF_X1 weight_queue_reg_1__2__0_ ( .D(n13777), .CK(clk), .Q(
        weight_queue_1__2__0_), .QN(n1484) );
  DFF_X1 weight_queue_reg_1__3__7_ ( .D(n13772), .CK(clk), .Q(
        weight_queue_1__3__7_), .QN(n1485) );
  DFF_X1 weight_queue_reg_1__3__6_ ( .D(n13767), .CK(clk), .Q(
        weight_queue_1__3__6_), .QN(n1486) );
  DFF_X1 weight_queue_reg_1__3__5_ ( .D(n13762), .CK(clk), .Q(
        weight_queue_1__3__5_), .QN(n1487) );
  DFF_X1 weight_queue_reg_1__3__4_ ( .D(n13757), .CK(clk), .Q(
        weight_queue_1__3__4_), .QN(n1488) );
  DFF_X1 weight_queue_reg_1__3__3_ ( .D(n13752), .CK(clk), .Q(
        weight_queue_1__3__3_), .QN(n1489) );
  DFF_X1 weight_queue_reg_1__3__2_ ( .D(n13747), .CK(clk), .Q(
        weight_queue_1__3__2_), .QN(n1490) );
  DFF_X1 weight_queue_reg_1__3__1_ ( .D(n13742), .CK(clk), .Q(
        weight_queue_1__3__1_), .QN(n1491) );
  DFF_X1 weight_queue_reg_1__3__0_ ( .D(n13737), .CK(clk), .Q(
        weight_queue_1__3__0_), .QN(n1492) );
  DFF_X1 weight_queue_reg_1__4__7_ ( .D(n13732), .CK(clk), .Q(
        weight_queue_1__4__7_), .QN(n1493) );
  DFF_X1 weight_queue_reg_1__4__6_ ( .D(n13727), .CK(clk), .Q(
        weight_queue_1__4__6_), .QN(n1494) );
  DFF_X1 weight_queue_reg_1__4__5_ ( .D(n13722), .CK(clk), .Q(
        weight_queue_1__4__5_), .QN(n1495) );
  DFF_X1 weight_queue_reg_1__4__4_ ( .D(n13717), .CK(clk), .Q(
        weight_queue_1__4__4_), .QN(n1496) );
  DFF_X1 weight_queue_reg_1__4__3_ ( .D(n13712), .CK(clk), .Q(
        weight_queue_1__4__3_), .QN(n1497) );
  DFF_X1 weight_queue_reg_1__4__2_ ( .D(n13707), .CK(clk), .Q(
        weight_queue_1__4__2_), .QN(n1498) );
  DFF_X1 weight_queue_reg_1__4__1_ ( .D(n13702), .CK(clk), .Q(
        weight_queue_1__4__1_), .QN(n1499) );
  DFF_X1 weight_queue_reg_1__4__0_ ( .D(n13697), .CK(clk), .Q(
        weight_queue_1__4__0_), .QN(n1500) );
  DFF_X1 weight_queue_reg_1__5__7_ ( .D(n13692), .CK(clk), .Q(
        weight_queue_1__5__7_), .QN(n1501) );
  DFF_X1 weight_queue_reg_1__5__6_ ( .D(n13687), .CK(clk), .Q(
        weight_queue_1__5__6_), .QN(n1502) );
  DFF_X1 weight_queue_reg_1__5__5_ ( .D(n13682), .CK(clk), .Q(
        weight_queue_1__5__5_), .QN(n1503) );
  DFF_X1 weight_queue_reg_1__5__4_ ( .D(n13677), .CK(clk), .Q(
        weight_queue_1__5__4_), .QN(n1504) );
  DFF_X1 weight_queue_reg_1__5__3_ ( .D(n13672), .CK(clk), .Q(
        weight_queue_1__5__3_), .QN(n1505) );
  DFF_X1 weight_queue_reg_1__5__2_ ( .D(n13667), .CK(clk), .Q(
        weight_queue_1__5__2_), .QN(n1506) );
  DFF_X1 weight_queue_reg_1__5__1_ ( .D(n13662), .CK(clk), .Q(
        weight_queue_1__5__1_), .QN(n1507) );
  DFF_X1 weight_queue_reg_1__5__0_ ( .D(n13657), .CK(clk), .Q(
        weight_queue_1__5__0_), .QN(n1508) );
  DFF_X1 weight_queue_reg_1__6__7_ ( .D(n13652), .CK(clk), .Q(
        weight_queue_1__6__7_), .QN(n1509) );
  DFF_X1 weight_queue_reg_1__6__6_ ( .D(n13647), .CK(clk), .Q(
        weight_queue_1__6__6_), .QN(n1510) );
  DFF_X1 weight_queue_reg_1__6__5_ ( .D(n13642), .CK(clk), .Q(
        weight_queue_1__6__5_), .QN(n1511) );
  DFF_X1 weight_queue_reg_1__6__4_ ( .D(n13637), .CK(clk), .Q(
        weight_queue_1__6__4_), .QN(n1512) );
  DFF_X1 weight_queue_reg_1__6__3_ ( .D(n13632), .CK(clk), .Q(
        weight_queue_1__6__3_), .QN(n1513) );
  DFF_X1 weight_queue_reg_1__6__2_ ( .D(n13627), .CK(clk), .Q(
        weight_queue_1__6__2_), .QN(n1514) );
  DFF_X1 weight_queue_reg_1__6__1_ ( .D(n13622), .CK(clk), .Q(
        weight_queue_1__6__1_), .QN(n1515) );
  DFF_X1 weight_queue_reg_1__6__0_ ( .D(n13617), .CK(clk), .Q(
        weight_queue_1__6__0_), .QN(n1516) );
  DFF_X1 weight_queue_reg_1__7__7_ ( .D(n13612), .CK(clk), .Q(
        weight_queue_1__7__7_), .QN(n1517) );
  DFF_X1 weight_queue_reg_1__7__6_ ( .D(n13607), .CK(clk), .Q(
        weight_queue_1__7__6_), .QN(n1518) );
  DFF_X1 weight_queue_reg_1__7__5_ ( .D(n13602), .CK(clk), .Q(
        weight_queue_1__7__5_), .QN(n1519) );
  DFF_X1 weight_queue_reg_1__7__4_ ( .D(n13597), .CK(clk), .Q(
        weight_queue_1__7__4_), .QN(n1520) );
  DFF_X1 weight_queue_reg_1__7__3_ ( .D(n13592), .CK(clk), .Q(
        weight_queue_1__7__3_), .QN(n1521) );
  DFF_X1 weight_queue_reg_1__7__2_ ( .D(n13587), .CK(clk), .Q(
        weight_queue_1__7__2_), .QN(n1522) );
  DFF_X1 weight_queue_reg_1__7__1_ ( .D(n13582), .CK(clk), .Q(
        weight_queue_1__7__1_), .QN(n1523) );
  DFF_X1 weight_queue_reg_1__7__0_ ( .D(n13577), .CK(clk), .Q(
        weight_queue_1__7__0_), .QN(n1524) );
  DFF_X1 weight_queue_reg_2__0__7_ ( .D(n13572), .CK(clk), .Q(
        weight_queue_2__0__7_), .QN(n1525) );
  DFF_X1 weight_queue_reg_2__0__6_ ( .D(n13567), .CK(clk), .Q(
        weight_queue_2__0__6_), .QN(n1526) );
  DFF_X1 weight_queue_reg_2__0__5_ ( .D(n13562), .CK(clk), .Q(
        weight_queue_2__0__5_), .QN(n1527) );
  DFF_X1 weight_queue_reg_2__0__4_ ( .D(n13557), .CK(clk), .Q(
        weight_queue_2__0__4_), .QN(n1528) );
  DFF_X1 weight_queue_reg_2__0__3_ ( .D(n13552), .CK(clk), .Q(
        weight_queue_2__0__3_), .QN(n1529) );
  DFF_X1 weight_queue_reg_2__0__2_ ( .D(n13547), .CK(clk), .Q(
        weight_queue_2__0__2_), .QN(n1530) );
  DFF_X1 weight_queue_reg_2__0__1_ ( .D(n13542), .CK(clk), .Q(
        weight_queue_2__0__1_), .QN(n1531) );
  DFF_X1 weight_queue_reg_2__0__0_ ( .D(n13537), .CK(clk), .Q(
        weight_queue_2__0__0_), .QN(n1532) );
  DFF_X1 weight_queue_reg_2__1__7_ ( .D(n13532), .CK(clk), .Q(
        weight_queue_2__1__7_), .QN(n1533) );
  DFF_X1 weight_queue_reg_2__1__6_ ( .D(n13527), .CK(clk), .Q(
        weight_queue_2__1__6_), .QN(n1534) );
  DFF_X1 weight_queue_reg_2__1__5_ ( .D(n13522), .CK(clk), .Q(
        weight_queue_2__1__5_), .QN(n1535) );
  DFF_X1 weight_queue_reg_2__1__4_ ( .D(n13517), .CK(clk), .Q(
        weight_queue_2__1__4_), .QN(n1536) );
  DFF_X1 weight_queue_reg_2__1__3_ ( .D(n13512), .CK(clk), .Q(
        weight_queue_2__1__3_), .QN(n1537) );
  DFF_X1 weight_queue_reg_2__1__2_ ( .D(n13507), .CK(clk), .Q(
        weight_queue_2__1__2_), .QN(n1538) );
  DFF_X1 weight_queue_reg_2__1__1_ ( .D(n13502), .CK(clk), .Q(
        weight_queue_2__1__1_), .QN(n1539) );
  DFF_X1 weight_queue_reg_2__1__0_ ( .D(n13497), .CK(clk), .Q(
        weight_queue_2__1__0_), .QN(n1540) );
  DFF_X1 weight_queue_reg_2__2__7_ ( .D(n13492), .CK(clk), .Q(
        weight_queue_2__2__7_), .QN(n1541) );
  DFF_X1 weight_queue_reg_2__2__6_ ( .D(n13487), .CK(clk), .Q(
        weight_queue_2__2__6_), .QN(n1542) );
  DFF_X1 weight_queue_reg_2__2__5_ ( .D(n13482), .CK(clk), .Q(
        weight_queue_2__2__5_), .QN(n1543) );
  DFF_X1 weight_queue_reg_2__2__4_ ( .D(n13477), .CK(clk), .Q(
        weight_queue_2__2__4_), .QN(n1544) );
  DFF_X1 weight_queue_reg_2__2__3_ ( .D(n13472), .CK(clk), .Q(
        weight_queue_2__2__3_), .QN(n1545) );
  DFF_X1 weight_queue_reg_2__2__2_ ( .D(n13467), .CK(clk), .Q(
        weight_queue_2__2__2_), .QN(n1546) );
  DFF_X1 weight_queue_reg_2__2__1_ ( .D(n13462), .CK(clk), .Q(
        weight_queue_2__2__1_), .QN(n1547) );
  DFF_X1 weight_queue_reg_2__2__0_ ( .D(n13457), .CK(clk), .Q(
        weight_queue_2__2__0_), .QN(n1548) );
  DFF_X1 weight_queue_reg_2__3__7_ ( .D(n13452), .CK(clk), .Q(
        weight_queue_2__3__7_), .QN(n1549) );
  DFF_X1 weight_queue_reg_2__3__6_ ( .D(n13447), .CK(clk), .Q(
        weight_queue_2__3__6_), .QN(n1550) );
  DFF_X1 weight_queue_reg_2__3__5_ ( .D(n13442), .CK(clk), .Q(
        weight_queue_2__3__5_), .QN(n1551) );
  DFF_X1 weight_queue_reg_2__3__4_ ( .D(n13437), .CK(clk), .Q(
        weight_queue_2__3__4_), .QN(n1552) );
  DFF_X1 weight_queue_reg_2__3__3_ ( .D(n13432), .CK(clk), .Q(
        weight_queue_2__3__3_), .QN(n1553) );
  DFF_X1 weight_queue_reg_2__3__2_ ( .D(n13427), .CK(clk), .Q(
        weight_queue_2__3__2_), .QN(n1554) );
  DFF_X1 weight_queue_reg_2__3__1_ ( .D(n13422), .CK(clk), .Q(
        weight_queue_2__3__1_), .QN(n1555) );
  DFF_X1 weight_queue_reg_2__3__0_ ( .D(n13417), .CK(clk), .Q(
        weight_queue_2__3__0_), .QN(n1556) );
  DFF_X1 weight_queue_reg_2__4__7_ ( .D(n13412), .CK(clk), .Q(
        weight_queue_2__4__7_), .QN(n1557) );
  DFF_X1 weight_queue_reg_2__4__6_ ( .D(n13407), .CK(clk), .Q(
        weight_queue_2__4__6_), .QN(n1558) );
  DFF_X1 weight_queue_reg_2__4__5_ ( .D(n13402), .CK(clk), .Q(
        weight_queue_2__4__5_), .QN(n1559) );
  DFF_X1 weight_queue_reg_2__4__4_ ( .D(n13397), .CK(clk), .Q(
        weight_queue_2__4__4_), .QN(n1560) );
  DFF_X1 weight_queue_reg_2__4__3_ ( .D(n13392), .CK(clk), .Q(
        weight_queue_2__4__3_), .QN(n1561) );
  DFF_X1 weight_queue_reg_2__4__2_ ( .D(n13387), .CK(clk), .Q(
        weight_queue_2__4__2_), .QN(n1562) );
  DFF_X1 weight_queue_reg_2__4__1_ ( .D(n13382), .CK(clk), .Q(
        weight_queue_2__4__1_), .QN(n1563) );
  DFF_X1 weight_queue_reg_2__4__0_ ( .D(n13377), .CK(clk), .Q(
        weight_queue_2__4__0_), .QN(n1564) );
  DFF_X1 weight_queue_reg_2__5__7_ ( .D(n13372), .CK(clk), .Q(
        weight_queue_2__5__7_), .QN(n1565) );
  DFF_X1 weight_queue_reg_2__5__6_ ( .D(n13367), .CK(clk), .Q(
        weight_queue_2__5__6_), .QN(n1566) );
  DFF_X1 weight_queue_reg_2__5__5_ ( .D(n13362), .CK(clk), .Q(
        weight_queue_2__5__5_), .QN(n1567) );
  DFF_X1 weight_queue_reg_2__5__4_ ( .D(n13357), .CK(clk), .Q(
        weight_queue_2__5__4_), .QN(n1568) );
  DFF_X1 weight_queue_reg_2__5__3_ ( .D(n13352), .CK(clk), .Q(
        weight_queue_2__5__3_), .QN(n1569) );
  DFF_X1 weight_queue_reg_2__5__2_ ( .D(n13347), .CK(clk), .Q(
        weight_queue_2__5__2_), .QN(n1570) );
  DFF_X1 weight_queue_reg_2__5__1_ ( .D(n13342), .CK(clk), .Q(
        weight_queue_2__5__1_), .QN(n1571) );
  DFF_X1 weight_queue_reg_2__5__0_ ( .D(n13337), .CK(clk), .Q(
        weight_queue_2__5__0_), .QN(n1572) );
  DFF_X1 weight_queue_reg_2__6__7_ ( .D(n13332), .CK(clk), .Q(
        weight_queue_2__6__7_), .QN(n1573) );
  DFF_X1 weight_queue_reg_2__6__6_ ( .D(n13327), .CK(clk), .Q(
        weight_queue_2__6__6_), .QN(n1574) );
  DFF_X1 weight_queue_reg_2__6__5_ ( .D(n13322), .CK(clk), .Q(
        weight_queue_2__6__5_), .QN(n1575) );
  DFF_X1 weight_queue_reg_2__6__4_ ( .D(n13317), .CK(clk), .Q(
        weight_queue_2__6__4_), .QN(n1576) );
  DFF_X1 weight_queue_reg_2__6__3_ ( .D(n13312), .CK(clk), .Q(
        weight_queue_2__6__3_), .QN(n1577) );
  DFF_X1 weight_queue_reg_2__6__2_ ( .D(n13307), .CK(clk), .Q(
        weight_queue_2__6__2_), .QN(n1578) );
  DFF_X1 weight_queue_reg_2__6__1_ ( .D(n13302), .CK(clk), .Q(
        weight_queue_2__6__1_), .QN(n1579) );
  DFF_X1 weight_queue_reg_2__6__0_ ( .D(n13297), .CK(clk), .Q(
        weight_queue_2__6__0_), .QN(n1580) );
  DFF_X1 weight_queue_reg_2__7__7_ ( .D(n13292), .CK(clk), .Q(
        weight_queue_2__7__7_), .QN(n1581) );
  DFF_X1 weight_queue_reg_2__7__6_ ( .D(n13287), .CK(clk), .Q(
        weight_queue_2__7__6_), .QN(n1582) );
  DFF_X1 weight_queue_reg_2__7__5_ ( .D(n13282), .CK(clk), .Q(
        weight_queue_2__7__5_), .QN(n1583) );
  DFF_X1 weight_queue_reg_2__7__4_ ( .D(n13277), .CK(clk), .Q(
        weight_queue_2__7__4_), .QN(n1584) );
  DFF_X1 weight_queue_reg_2__7__3_ ( .D(n13272), .CK(clk), .Q(
        weight_queue_2__7__3_), .QN(n1585) );
  DFF_X1 weight_queue_reg_2__7__2_ ( .D(n13267), .CK(clk), .Q(
        weight_queue_2__7__2_), .QN(n1586) );
  DFF_X1 weight_queue_reg_2__7__1_ ( .D(n13262), .CK(clk), .Q(
        weight_queue_2__7__1_), .QN(n1587) );
  DFF_X1 weight_queue_reg_2__7__0_ ( .D(n13257), .CK(clk), .Q(
        weight_queue_2__7__0_), .QN(n1588) );
  DFF_X1 weight_queue_reg_3__0__7_ ( .D(n13252), .CK(clk), .Q(
        weight_queue_3__0__7_), .QN(n1589) );
  DFF_X1 weight_queue_reg_3__0__6_ ( .D(n13247), .CK(clk), .Q(
        weight_queue_3__0__6_), .QN(n1590) );
  DFF_X1 weight_queue_reg_3__0__5_ ( .D(n13242), .CK(clk), .Q(
        weight_queue_3__0__5_), .QN(n1591) );
  DFF_X1 weight_queue_reg_3__0__4_ ( .D(n13237), .CK(clk), .Q(
        weight_queue_3__0__4_), .QN(n1592) );
  DFF_X1 weight_queue_reg_3__0__3_ ( .D(n13232), .CK(clk), .Q(
        weight_queue_3__0__3_), .QN(n1593) );
  DFF_X1 weight_queue_reg_3__0__2_ ( .D(n13227), .CK(clk), .Q(
        weight_queue_3__0__2_), .QN(n1594) );
  DFF_X1 weight_queue_reg_3__0__1_ ( .D(n13222), .CK(clk), .Q(
        weight_queue_3__0__1_), .QN(n1595) );
  DFF_X1 weight_queue_reg_3__0__0_ ( .D(n13217), .CK(clk), .Q(
        weight_queue_3__0__0_), .QN(n1596) );
  DFF_X1 weight_queue_reg_3__1__7_ ( .D(n13212), .CK(clk), .Q(
        weight_queue_3__1__7_), .QN(n1597) );
  DFF_X1 weight_queue_reg_3__1__6_ ( .D(n13207), .CK(clk), .Q(
        weight_queue_3__1__6_), .QN(n1598) );
  DFF_X1 weight_queue_reg_3__1__5_ ( .D(n13202), .CK(clk), .Q(
        weight_queue_3__1__5_), .QN(n1599) );
  DFF_X1 weight_queue_reg_3__1__4_ ( .D(n13197), .CK(clk), .Q(
        weight_queue_3__1__4_), .QN(n1600) );
  DFF_X1 weight_queue_reg_3__1__3_ ( .D(n13192), .CK(clk), .Q(
        weight_queue_3__1__3_), .QN(n1601) );
  DFF_X1 weight_queue_reg_3__1__2_ ( .D(n13187), .CK(clk), .Q(
        weight_queue_3__1__2_), .QN(n1602) );
  DFF_X1 weight_queue_reg_3__1__1_ ( .D(n13182), .CK(clk), .Q(
        weight_queue_3__1__1_), .QN(n1603) );
  DFF_X1 weight_queue_reg_3__1__0_ ( .D(n13177), .CK(clk), .Q(
        weight_queue_3__1__0_), .QN(n1604) );
  DFF_X1 weight_queue_reg_3__2__7_ ( .D(n13172), .CK(clk), .Q(
        weight_queue_3__2__7_), .QN(n1605) );
  DFF_X1 weight_queue_reg_3__2__6_ ( .D(n13167), .CK(clk), .Q(
        weight_queue_3__2__6_), .QN(n1606) );
  DFF_X1 weight_queue_reg_3__2__5_ ( .D(n13162), .CK(clk), .Q(
        weight_queue_3__2__5_), .QN(n1607) );
  DFF_X1 weight_queue_reg_3__2__4_ ( .D(n13157), .CK(clk), .Q(
        weight_queue_3__2__4_), .QN(n1608) );
  DFF_X1 weight_queue_reg_3__2__3_ ( .D(n13152), .CK(clk), .Q(
        weight_queue_3__2__3_), .QN(n1609) );
  DFF_X1 weight_queue_reg_3__2__2_ ( .D(n13147), .CK(clk), .Q(
        weight_queue_3__2__2_), .QN(n1610) );
  DFF_X1 weight_queue_reg_3__2__1_ ( .D(n13142), .CK(clk), .Q(
        weight_queue_3__2__1_), .QN(n1611) );
  DFF_X1 weight_queue_reg_3__2__0_ ( .D(n13137), .CK(clk), .Q(
        weight_queue_3__2__0_), .QN(n1612) );
  DFF_X1 weight_queue_reg_3__3__7_ ( .D(n13132), .CK(clk), .Q(
        weight_queue_3__3__7_), .QN(n1613) );
  DFF_X1 weight_queue_reg_3__3__6_ ( .D(n13127), .CK(clk), .Q(
        weight_queue_3__3__6_), .QN(n1614) );
  DFF_X1 weight_queue_reg_3__3__5_ ( .D(n13122), .CK(clk), .Q(
        weight_queue_3__3__5_), .QN(n1615) );
  DFF_X1 weight_queue_reg_3__3__4_ ( .D(n13117), .CK(clk), .Q(
        weight_queue_3__3__4_), .QN(n1616) );
  DFF_X1 weight_queue_reg_3__3__3_ ( .D(n13112), .CK(clk), .Q(
        weight_queue_3__3__3_), .QN(n1617) );
  DFF_X1 weight_queue_reg_3__3__2_ ( .D(n13107), .CK(clk), .Q(
        weight_queue_3__3__2_), .QN(n1618) );
  DFF_X1 weight_queue_reg_3__3__1_ ( .D(n13102), .CK(clk), .Q(
        weight_queue_3__3__1_), .QN(n1619) );
  DFF_X1 weight_queue_reg_3__3__0_ ( .D(n13097), .CK(clk), .Q(
        weight_queue_3__3__0_), .QN(n1620) );
  DFF_X1 weight_queue_reg_3__4__7_ ( .D(n13092), .CK(clk), .Q(
        weight_queue_3__4__7_), .QN(n1621) );
  DFF_X1 weight_queue_reg_3__4__6_ ( .D(n13087), .CK(clk), .Q(
        weight_queue_3__4__6_), .QN(n1622) );
  DFF_X1 weight_queue_reg_3__4__5_ ( .D(n13082), .CK(clk), .Q(
        weight_queue_3__4__5_), .QN(n1623) );
  DFF_X1 weight_queue_reg_3__4__4_ ( .D(n13077), .CK(clk), .Q(
        weight_queue_3__4__4_), .QN(n1624) );
  DFF_X1 weight_queue_reg_3__4__3_ ( .D(n13072), .CK(clk), .Q(
        weight_queue_3__4__3_), .QN(n1625) );
  DFF_X1 weight_queue_reg_3__4__2_ ( .D(n13067), .CK(clk), .Q(
        weight_queue_3__4__2_), .QN(n1626) );
  DFF_X1 weight_queue_reg_3__4__1_ ( .D(n13062), .CK(clk), .Q(
        weight_queue_3__4__1_), .QN(n1627) );
  DFF_X1 weight_queue_reg_3__4__0_ ( .D(n13057), .CK(clk), .Q(
        weight_queue_3__4__0_), .QN(n1628) );
  DFF_X1 weight_queue_reg_3__5__7_ ( .D(n13052), .CK(clk), .Q(
        weight_queue_3__5__7_), .QN(n1629) );
  DFF_X1 weight_queue_reg_3__5__6_ ( .D(n13047), .CK(clk), .Q(
        weight_queue_3__5__6_), .QN(n1630) );
  DFF_X1 weight_queue_reg_3__5__5_ ( .D(n13042), .CK(clk), .Q(
        weight_queue_3__5__5_), .QN(n1631) );
  DFF_X1 weight_queue_reg_3__5__4_ ( .D(n13037), .CK(clk), .Q(
        weight_queue_3__5__4_), .QN(n1632) );
  DFF_X1 weight_queue_reg_3__5__3_ ( .D(n13032), .CK(clk), .Q(
        weight_queue_3__5__3_), .QN(n1633) );
  DFF_X1 weight_queue_reg_3__5__2_ ( .D(n13027), .CK(clk), .Q(
        weight_queue_3__5__2_), .QN(n1634) );
  DFF_X1 weight_queue_reg_3__5__1_ ( .D(n13022), .CK(clk), .Q(
        weight_queue_3__5__1_), .QN(n1635) );
  DFF_X1 weight_queue_reg_3__5__0_ ( .D(n13017), .CK(clk), .Q(
        weight_queue_3__5__0_), .QN(n1636) );
  DFF_X1 weight_queue_reg_3__6__7_ ( .D(n13012), .CK(clk), .Q(
        weight_queue_3__6__7_), .QN(n1637) );
  DFF_X1 weight_queue_reg_3__6__6_ ( .D(n13007), .CK(clk), .Q(
        weight_queue_3__6__6_), .QN(n1638) );
  DFF_X1 weight_queue_reg_3__6__5_ ( .D(n13002), .CK(clk), .Q(
        weight_queue_3__6__5_), .QN(n1639) );
  DFF_X1 weight_queue_reg_3__6__4_ ( .D(n12997), .CK(clk), .Q(
        weight_queue_3__6__4_), .QN(n1640) );
  DFF_X1 weight_queue_reg_3__6__3_ ( .D(n12992), .CK(clk), .Q(
        weight_queue_3__6__3_), .QN(n1641) );
  DFF_X1 weight_queue_reg_3__6__2_ ( .D(n12987), .CK(clk), .Q(
        weight_queue_3__6__2_), .QN(n1642) );
  DFF_X1 weight_queue_reg_3__6__1_ ( .D(n12982), .CK(clk), .Q(
        weight_queue_3__6__1_), .QN(n1643) );
  DFF_X1 weight_queue_reg_3__6__0_ ( .D(n12977), .CK(clk), .Q(
        weight_queue_3__6__0_), .QN(n1644) );
  DFF_X1 weight_queue_reg_3__7__7_ ( .D(n12972), .CK(clk), .Q(
        weight_queue_3__7__7_), .QN(n1645) );
  DFF_X1 weight_queue_reg_3__7__6_ ( .D(n12967), .CK(clk), .Q(
        weight_queue_3__7__6_), .QN(n1646) );
  DFF_X1 weight_queue_reg_3__7__5_ ( .D(n12962), .CK(clk), .Q(
        weight_queue_3__7__5_), .QN(n1647) );
  DFF_X1 weight_queue_reg_3__7__4_ ( .D(n12957), .CK(clk), .Q(
        weight_queue_3__7__4_), .QN(n1648) );
  DFF_X1 weight_queue_reg_3__7__3_ ( .D(n12952), .CK(clk), .Q(
        weight_queue_3__7__3_), .QN(n1649) );
  DFF_X1 weight_queue_reg_3__7__2_ ( .D(n12947), .CK(clk), .Q(
        weight_queue_3__7__2_), .QN(n1650) );
  DFF_X1 weight_queue_reg_3__7__1_ ( .D(n12942), .CK(clk), .Q(
        weight_queue_3__7__1_), .QN(n1651) );
  DFF_X1 weight_queue_reg_3__7__0_ ( .D(n12937), .CK(clk), .Q(
        weight_queue_3__7__0_), .QN(n1652) );
  DFF_X1 weight_queue_reg_4__0__7_ ( .D(n12932), .CK(clk), .Q(
        weight_queue_4__0__7_), .QN(n1653) );
  DFF_X1 weight_queue_reg_4__0__6_ ( .D(n12927), .CK(clk), .Q(
        weight_queue_4__0__6_), .QN(n1654) );
  DFF_X1 weight_queue_reg_4__0__5_ ( .D(n12922), .CK(clk), .Q(
        weight_queue_4__0__5_), .QN(n1655) );
  DFF_X1 weight_queue_reg_4__0__4_ ( .D(n12917), .CK(clk), .Q(
        weight_queue_4__0__4_), .QN(n1656) );
  DFF_X1 weight_queue_reg_4__0__3_ ( .D(n12912), .CK(clk), .Q(
        weight_queue_4__0__3_), .QN(n1657) );
  DFF_X1 weight_queue_reg_4__0__2_ ( .D(n12907), .CK(clk), .Q(
        weight_queue_4__0__2_), .QN(n1658) );
  DFF_X1 weight_queue_reg_4__0__1_ ( .D(n12902), .CK(clk), .Q(
        weight_queue_4__0__1_), .QN(n1659) );
  DFF_X1 weight_queue_reg_4__0__0_ ( .D(n12897), .CK(clk), .Q(
        weight_queue_4__0__0_), .QN(n1660) );
  DFF_X1 weight_queue_reg_4__1__7_ ( .D(n12892), .CK(clk), .Q(
        weight_queue_4__1__7_), .QN(n1661) );
  DFF_X1 weight_queue_reg_4__1__6_ ( .D(n12887), .CK(clk), .Q(
        weight_queue_4__1__6_), .QN(n1662) );
  DFF_X1 weight_queue_reg_4__1__5_ ( .D(n12882), .CK(clk), .Q(
        weight_queue_4__1__5_), .QN(n1663) );
  DFF_X1 weight_queue_reg_4__1__4_ ( .D(n12877), .CK(clk), .Q(
        weight_queue_4__1__4_), .QN(n1664) );
  DFF_X1 weight_queue_reg_4__1__3_ ( .D(n12872), .CK(clk), .Q(
        weight_queue_4__1__3_), .QN(n1665) );
  DFF_X1 weight_queue_reg_4__1__2_ ( .D(n12867), .CK(clk), .Q(
        weight_queue_4__1__2_), .QN(n1666) );
  DFF_X1 weight_queue_reg_4__1__1_ ( .D(n12862), .CK(clk), .Q(
        weight_queue_4__1__1_), .QN(n1667) );
  DFF_X1 weight_queue_reg_4__1__0_ ( .D(n12857), .CK(clk), .Q(
        weight_queue_4__1__0_), .QN(n1668) );
  DFF_X1 weight_queue_reg_4__2__7_ ( .D(n12852), .CK(clk), .Q(
        weight_queue_4__2__7_), .QN(n1669) );
  DFF_X1 weight_queue_reg_4__2__6_ ( .D(n12847), .CK(clk), .Q(
        weight_queue_4__2__6_), .QN(n1670) );
  DFF_X1 weight_queue_reg_4__2__5_ ( .D(n12842), .CK(clk), .Q(
        weight_queue_4__2__5_), .QN(n1671) );
  DFF_X1 weight_queue_reg_4__2__4_ ( .D(n12837), .CK(clk), .Q(
        weight_queue_4__2__4_), .QN(n1672) );
  DFF_X1 weight_queue_reg_4__2__3_ ( .D(n12832), .CK(clk), .Q(
        weight_queue_4__2__3_), .QN(n1673) );
  DFF_X1 weight_queue_reg_4__2__2_ ( .D(n12827), .CK(clk), .Q(
        weight_queue_4__2__2_), .QN(n1674) );
  DFF_X1 weight_queue_reg_4__2__1_ ( .D(n12822), .CK(clk), .Q(
        weight_queue_4__2__1_), .QN(n1675) );
  DFF_X1 weight_queue_reg_4__2__0_ ( .D(n12817), .CK(clk), .Q(
        weight_queue_4__2__0_), .QN(n1676) );
  DFF_X1 weight_queue_reg_4__3__7_ ( .D(n12812), .CK(clk), .Q(
        weight_queue_4__3__7_), .QN(n1677) );
  DFF_X1 weight_queue_reg_4__3__6_ ( .D(n12807), .CK(clk), .Q(
        weight_queue_4__3__6_), .QN(n1678) );
  DFF_X1 weight_queue_reg_4__3__5_ ( .D(n12802), .CK(clk), .Q(
        weight_queue_4__3__5_), .QN(n1679) );
  DFF_X1 weight_queue_reg_4__3__4_ ( .D(n12797), .CK(clk), .Q(
        weight_queue_4__3__4_), .QN(n1680) );
  DFF_X1 weight_queue_reg_4__3__3_ ( .D(n12792), .CK(clk), .Q(
        weight_queue_4__3__3_), .QN(n1681) );
  DFF_X1 weight_queue_reg_4__3__2_ ( .D(n12787), .CK(clk), .Q(
        weight_queue_4__3__2_), .QN(n1682) );
  DFF_X1 weight_queue_reg_4__3__1_ ( .D(n12782), .CK(clk), .Q(
        weight_queue_4__3__1_), .QN(n1683) );
  DFF_X1 weight_queue_reg_4__3__0_ ( .D(n12777), .CK(clk), .Q(
        weight_queue_4__3__0_), .QN(n1684) );
  DFF_X1 weight_queue_reg_4__4__7_ ( .D(n12772), .CK(clk), .Q(
        weight_queue_4__4__7_), .QN(n1685) );
  DFF_X1 weight_queue_reg_4__4__6_ ( .D(n12767), .CK(clk), .Q(
        weight_queue_4__4__6_), .QN(n1686) );
  DFF_X1 weight_queue_reg_4__4__5_ ( .D(n12762), .CK(clk), .Q(
        weight_queue_4__4__5_), .QN(n1687) );
  DFF_X1 weight_queue_reg_4__4__4_ ( .D(n12757), .CK(clk), .Q(
        weight_queue_4__4__4_), .QN(n1688) );
  DFF_X1 weight_queue_reg_4__4__3_ ( .D(n12752), .CK(clk), .Q(
        weight_queue_4__4__3_), .QN(n1689) );
  DFF_X1 weight_queue_reg_4__4__2_ ( .D(n12747), .CK(clk), .Q(
        weight_queue_4__4__2_), .QN(n1690) );
  DFF_X1 weight_queue_reg_4__4__1_ ( .D(n12742), .CK(clk), .Q(
        weight_queue_4__4__1_), .QN(n1691) );
  DFF_X1 weight_queue_reg_4__4__0_ ( .D(n12737), .CK(clk), .Q(
        weight_queue_4__4__0_), .QN(n1692) );
  DFF_X1 weight_queue_reg_4__5__7_ ( .D(n12732), .CK(clk), .Q(
        weight_queue_4__5__7_), .QN(n1693) );
  DFF_X1 weight_queue_reg_4__5__6_ ( .D(n12727), .CK(clk), .Q(
        weight_queue_4__5__6_), .QN(n1694) );
  DFF_X1 weight_queue_reg_4__5__5_ ( .D(n12722), .CK(clk), .Q(
        weight_queue_4__5__5_), .QN(n1695) );
  DFF_X1 weight_queue_reg_4__5__4_ ( .D(n12717), .CK(clk), .Q(
        weight_queue_4__5__4_), .QN(n1696) );
  DFF_X1 weight_queue_reg_4__5__3_ ( .D(n12712), .CK(clk), .Q(
        weight_queue_4__5__3_), .QN(n1697) );
  DFF_X1 weight_queue_reg_4__5__2_ ( .D(n12707), .CK(clk), .Q(
        weight_queue_4__5__2_), .QN(n1698) );
  DFF_X1 weight_queue_reg_4__5__1_ ( .D(n12702), .CK(clk), .Q(
        weight_queue_4__5__1_), .QN(n1699) );
  DFF_X1 weight_queue_reg_4__5__0_ ( .D(n12697), .CK(clk), .Q(
        weight_queue_4__5__0_), .QN(n1700) );
  DFF_X1 weight_queue_reg_4__6__7_ ( .D(n12692), .CK(clk), .Q(
        weight_queue_4__6__7_), .QN(n1701) );
  DFF_X1 weight_queue_reg_4__6__6_ ( .D(n12687), .CK(clk), .Q(
        weight_queue_4__6__6_), .QN(n1702) );
  DFF_X1 weight_queue_reg_4__6__5_ ( .D(n12682), .CK(clk), .Q(
        weight_queue_4__6__5_), .QN(n1703) );
  DFF_X1 weight_queue_reg_4__6__4_ ( .D(n12677), .CK(clk), .Q(
        weight_queue_4__6__4_), .QN(n1704) );
  DFF_X1 weight_queue_reg_4__6__3_ ( .D(n12672), .CK(clk), .Q(
        weight_queue_4__6__3_), .QN(n1705) );
  DFF_X1 weight_queue_reg_4__6__2_ ( .D(n12667), .CK(clk), .Q(
        weight_queue_4__6__2_), .QN(n1706) );
  DFF_X1 weight_queue_reg_4__6__1_ ( .D(n12662), .CK(clk), .Q(
        weight_queue_4__6__1_), .QN(n1707) );
  DFF_X1 weight_queue_reg_4__6__0_ ( .D(n12657), .CK(clk), .Q(
        weight_queue_4__6__0_), .QN(n1708) );
  DFF_X1 weight_queue_reg_4__7__7_ ( .D(n12652), .CK(clk), .Q(
        weight_queue_4__7__7_), .QN(n1709) );
  DFF_X1 weight_queue_reg_4__7__6_ ( .D(n12647), .CK(clk), .Q(
        weight_queue_4__7__6_), .QN(n1710) );
  DFF_X1 weight_queue_reg_4__7__5_ ( .D(n12642), .CK(clk), .Q(
        weight_queue_4__7__5_), .QN(n1711) );
  DFF_X1 weight_queue_reg_4__7__4_ ( .D(n12637), .CK(clk), .Q(
        weight_queue_4__7__4_), .QN(n1712) );
  DFF_X1 weight_queue_reg_4__7__3_ ( .D(n12632), .CK(clk), .Q(
        weight_queue_4__7__3_), .QN(n1713) );
  DFF_X1 weight_queue_reg_4__7__2_ ( .D(n12627), .CK(clk), .Q(
        weight_queue_4__7__2_), .QN(n1714) );
  DFF_X1 weight_queue_reg_4__7__1_ ( .D(n12622), .CK(clk), .Q(
        weight_queue_4__7__1_), .QN(n1715) );
  DFF_X1 weight_queue_reg_4__7__0_ ( .D(n12617), .CK(clk), .Q(
        weight_queue_4__7__0_), .QN(n1716) );
  DFF_X1 weight_queue_reg_5__0__7_ ( .D(n12612), .CK(clk), .Q(
        weight_queue_5__0__7_), .QN(n1717) );
  DFF_X1 weight_queue_reg_5__0__6_ ( .D(n12607), .CK(clk), .Q(
        weight_queue_5__0__6_), .QN(n1718) );
  DFF_X1 weight_queue_reg_5__0__5_ ( .D(n12602), .CK(clk), .Q(
        weight_queue_5__0__5_), .QN(n1719) );
  DFF_X1 weight_queue_reg_5__0__4_ ( .D(n12597), .CK(clk), .Q(
        weight_queue_5__0__4_), .QN(n1720) );
  DFF_X1 weight_queue_reg_5__0__3_ ( .D(n12592), .CK(clk), .Q(
        weight_queue_5__0__3_), .QN(n1721) );
  DFF_X1 weight_queue_reg_5__0__2_ ( .D(n12587), .CK(clk), .Q(
        weight_queue_5__0__2_), .QN(n1722) );
  DFF_X1 weight_queue_reg_5__0__1_ ( .D(n12582), .CK(clk), .Q(
        weight_queue_5__0__1_), .QN(n1723) );
  DFF_X1 weight_queue_reg_5__0__0_ ( .D(n12577), .CK(clk), .Q(
        weight_queue_5__0__0_), .QN(n1724) );
  DFF_X1 weight_queue_reg_5__1__7_ ( .D(n12572), .CK(clk), .Q(
        weight_queue_5__1__7_), .QN(n1725) );
  DFF_X1 weight_queue_reg_5__1__6_ ( .D(n12567), .CK(clk), .Q(
        weight_queue_5__1__6_), .QN(n1726) );
  DFF_X1 weight_queue_reg_5__1__5_ ( .D(n12562), .CK(clk), .Q(
        weight_queue_5__1__5_), .QN(n1727) );
  DFF_X1 weight_queue_reg_5__1__4_ ( .D(n12557), .CK(clk), .Q(
        weight_queue_5__1__4_), .QN(n1728) );
  DFF_X1 weight_queue_reg_5__1__3_ ( .D(n12552), .CK(clk), .Q(
        weight_queue_5__1__3_), .QN(n1729) );
  DFF_X1 weight_queue_reg_5__1__2_ ( .D(n12547), .CK(clk), .Q(
        weight_queue_5__1__2_), .QN(n1730) );
  DFF_X1 weight_queue_reg_5__1__1_ ( .D(n12542), .CK(clk), .Q(
        weight_queue_5__1__1_), .QN(n1731) );
  DFF_X1 weight_queue_reg_5__1__0_ ( .D(n12537), .CK(clk), .Q(
        weight_queue_5__1__0_), .QN(n1732) );
  DFF_X1 weight_queue_reg_5__2__7_ ( .D(n12532), .CK(clk), .Q(
        weight_queue_5__2__7_), .QN(n1733) );
  DFF_X1 weight_queue_reg_5__2__6_ ( .D(n12527), .CK(clk), .Q(
        weight_queue_5__2__6_), .QN(n1734) );
  DFF_X1 weight_queue_reg_5__2__5_ ( .D(n12522), .CK(clk), .Q(
        weight_queue_5__2__5_), .QN(n1735) );
  DFF_X1 weight_queue_reg_5__2__4_ ( .D(n12517), .CK(clk), .Q(
        weight_queue_5__2__4_), .QN(n1736) );
  DFF_X1 weight_queue_reg_5__2__3_ ( .D(n12512), .CK(clk), .Q(
        weight_queue_5__2__3_), .QN(n1737) );
  DFF_X1 weight_queue_reg_5__2__2_ ( .D(n12507), .CK(clk), .Q(
        weight_queue_5__2__2_), .QN(n1738) );
  DFF_X1 weight_queue_reg_5__2__1_ ( .D(n12502), .CK(clk), .Q(
        weight_queue_5__2__1_), .QN(n1739) );
  DFF_X1 weight_queue_reg_5__2__0_ ( .D(n12497), .CK(clk), .Q(
        weight_queue_5__2__0_), .QN(n1740) );
  DFF_X1 weight_queue_reg_5__3__7_ ( .D(n12492), .CK(clk), .Q(
        weight_queue_5__3__7_), .QN(n1741) );
  DFF_X1 weight_queue_reg_5__3__6_ ( .D(n12487), .CK(clk), .Q(
        weight_queue_5__3__6_), .QN(n1742) );
  DFF_X1 weight_queue_reg_5__3__5_ ( .D(n12482), .CK(clk), .Q(
        weight_queue_5__3__5_), .QN(n1743) );
  DFF_X1 weight_queue_reg_5__3__4_ ( .D(n12477), .CK(clk), .Q(
        weight_queue_5__3__4_), .QN(n1744) );
  DFF_X1 weight_queue_reg_5__3__3_ ( .D(n12472), .CK(clk), .Q(
        weight_queue_5__3__3_), .QN(n1745) );
  DFF_X1 weight_queue_reg_5__3__2_ ( .D(n12467), .CK(clk), .Q(
        weight_queue_5__3__2_), .QN(n1746) );
  DFF_X1 weight_queue_reg_5__3__1_ ( .D(n12462), .CK(clk), .Q(
        weight_queue_5__3__1_), .QN(n1747) );
  DFF_X1 weight_queue_reg_5__3__0_ ( .D(n12457), .CK(clk), .Q(
        weight_queue_5__3__0_), .QN(n1748) );
  DFF_X1 weight_queue_reg_5__4__7_ ( .D(n12452), .CK(clk), .Q(
        weight_queue_5__4__7_), .QN(n1749) );
  DFF_X1 weight_queue_reg_5__4__6_ ( .D(n12447), .CK(clk), .Q(
        weight_queue_5__4__6_), .QN(n1750) );
  DFF_X1 weight_queue_reg_5__4__5_ ( .D(n12442), .CK(clk), .Q(
        weight_queue_5__4__5_), .QN(n1751) );
  DFF_X1 weight_queue_reg_5__4__4_ ( .D(n12437), .CK(clk), .Q(
        weight_queue_5__4__4_), .QN(n1752) );
  DFF_X1 weight_queue_reg_5__4__3_ ( .D(n12432), .CK(clk), .Q(
        weight_queue_5__4__3_), .QN(n1753) );
  DFF_X1 weight_queue_reg_5__4__2_ ( .D(n12427), .CK(clk), .Q(
        weight_queue_5__4__2_), .QN(n1754) );
  DFF_X1 weight_queue_reg_5__4__1_ ( .D(n12422), .CK(clk), .Q(
        weight_queue_5__4__1_), .QN(n1755) );
  DFF_X1 weight_queue_reg_5__4__0_ ( .D(n12417), .CK(clk), .Q(
        weight_queue_5__4__0_), .QN(n1756) );
  DFF_X1 weight_queue_reg_5__5__7_ ( .D(n12412), .CK(clk), .Q(
        weight_queue_5__5__7_), .QN(n1757) );
  DFF_X1 weight_queue_reg_5__5__6_ ( .D(n12407), .CK(clk), .Q(
        weight_queue_5__5__6_), .QN(n1758) );
  DFF_X1 weight_queue_reg_5__5__5_ ( .D(n12402), .CK(clk), .Q(
        weight_queue_5__5__5_), .QN(n1759) );
  DFF_X1 weight_queue_reg_5__5__4_ ( .D(n12397), .CK(clk), .Q(
        weight_queue_5__5__4_), .QN(n1760) );
  DFF_X1 weight_queue_reg_5__5__3_ ( .D(n12392), .CK(clk), .Q(
        weight_queue_5__5__3_), .QN(n1761) );
  DFF_X1 weight_queue_reg_5__5__2_ ( .D(n12387), .CK(clk), .Q(
        weight_queue_5__5__2_), .QN(n1762) );
  DFF_X1 weight_queue_reg_5__5__1_ ( .D(n12382), .CK(clk), .Q(
        weight_queue_5__5__1_), .QN(n1763) );
  DFF_X1 weight_queue_reg_5__5__0_ ( .D(n12377), .CK(clk), .Q(
        weight_queue_5__5__0_), .QN(n1764) );
  DFF_X1 weight_queue_reg_5__6__7_ ( .D(n12372), .CK(clk), .Q(
        weight_queue_5__6__7_), .QN(n1765) );
  DFF_X1 weight_queue_reg_5__6__6_ ( .D(n12367), .CK(clk), .Q(
        weight_queue_5__6__6_), .QN(n1766) );
  DFF_X1 weight_queue_reg_5__6__5_ ( .D(n12362), .CK(clk), .Q(
        weight_queue_5__6__5_), .QN(n1767) );
  DFF_X1 weight_queue_reg_5__6__4_ ( .D(n12357), .CK(clk), .Q(
        weight_queue_5__6__4_), .QN(n1768) );
  DFF_X1 weight_queue_reg_5__6__3_ ( .D(n12352), .CK(clk), .Q(
        weight_queue_5__6__3_), .QN(n1769) );
  DFF_X1 weight_queue_reg_5__6__2_ ( .D(n12347), .CK(clk), .Q(
        weight_queue_5__6__2_), .QN(n1770) );
  DFF_X1 weight_queue_reg_5__6__1_ ( .D(n12342), .CK(clk), .Q(
        weight_queue_5__6__1_), .QN(n1771) );
  DFF_X1 weight_queue_reg_5__6__0_ ( .D(n12337), .CK(clk), .Q(
        weight_queue_5__6__0_), .QN(n1772) );
  DFF_X1 weight_queue_reg_5__7__7_ ( .D(n12332), .CK(clk), .Q(
        weight_queue_5__7__7_), .QN(n1773) );
  DFF_X1 weight_queue_reg_5__7__6_ ( .D(n12327), .CK(clk), .Q(
        weight_queue_5__7__6_), .QN(n1774) );
  DFF_X1 weight_queue_reg_5__7__5_ ( .D(n12322), .CK(clk), .Q(
        weight_queue_5__7__5_), .QN(n1775) );
  DFF_X1 weight_queue_reg_5__7__4_ ( .D(n12317), .CK(clk), .Q(
        weight_queue_5__7__4_), .QN(n1776) );
  DFF_X1 weight_queue_reg_5__7__3_ ( .D(n12312), .CK(clk), .Q(
        weight_queue_5__7__3_), .QN(n1777) );
  DFF_X1 weight_queue_reg_5__7__2_ ( .D(n12307), .CK(clk), .Q(
        weight_queue_5__7__2_), .QN(n1778) );
  DFF_X1 weight_queue_reg_5__7__1_ ( .D(n12302), .CK(clk), .Q(
        weight_queue_5__7__1_), .QN(n1779) );
  DFF_X1 weight_queue_reg_5__7__0_ ( .D(n12297), .CK(clk), .Q(
        weight_queue_5__7__0_), .QN(n1780) );
  DFF_X1 weight_queue_reg_6__0__7_ ( .D(n12290), .CK(clk), .Q(
        weight_queue_6__0__7_), .QN(n1781) );
  DFF_X1 weight_queue_reg_6__0__6_ ( .D(n12283), .CK(clk), .Q(
        weight_queue_6__0__6_), .QN(n1782) );
  DFF_X1 weight_queue_reg_6__0__5_ ( .D(n12276), .CK(clk), .Q(
        weight_queue_6__0__5_), .QN(n1783) );
  DFF_X1 weight_queue_reg_6__0__4_ ( .D(n12269), .CK(clk), .Q(
        weight_queue_6__0__4_), .QN(n1784) );
  DFF_X1 weight_queue_reg_6__0__3_ ( .D(n12262), .CK(clk), .Q(
        weight_queue_6__0__3_), .QN(n1785) );
  DFF_X1 weight_queue_reg_6__0__2_ ( .D(n12255), .CK(clk), .Q(
        weight_queue_6__0__2_), .QN(n1786) );
  DFF_X1 weight_queue_reg_6__0__1_ ( .D(n12248), .CK(clk), .Q(
        weight_queue_6__0__1_), .QN(n1787) );
  DFF_X1 weight_queue_reg_6__0__0_ ( .D(n12241), .CK(clk), .Q(
        weight_queue_6__0__0_), .QN(n1788) );
  DFF_X1 weight_queue_reg_6__1__7_ ( .D(n12234), .CK(clk), .Q(
        weight_queue_6__1__7_), .QN(n1789) );
  DFF_X1 weight_queue_reg_6__1__6_ ( .D(n12227), .CK(clk), .Q(
        weight_queue_6__1__6_), .QN(n1790) );
  DFF_X1 weight_queue_reg_6__1__5_ ( .D(n12220), .CK(clk), .Q(
        weight_queue_6__1__5_), .QN(n1791) );
  DFF_X1 weight_queue_reg_6__1__4_ ( .D(n12213), .CK(clk), .Q(
        weight_queue_6__1__4_), .QN(n1792) );
  DFF_X1 weight_queue_reg_6__1__3_ ( .D(n12206), .CK(clk), .Q(
        weight_queue_6__1__3_), .QN(n1793) );
  DFF_X1 weight_queue_reg_6__1__2_ ( .D(n12199), .CK(clk), .Q(
        weight_queue_6__1__2_), .QN(n1794) );
  DFF_X1 weight_queue_reg_6__1__1_ ( .D(n12192), .CK(clk), .Q(
        weight_queue_6__1__1_), .QN(n1795) );
  DFF_X1 weight_queue_reg_6__1__0_ ( .D(n12185), .CK(clk), .Q(
        weight_queue_6__1__0_), .QN(n1796) );
  DFF_X1 weight_queue_reg_6__2__7_ ( .D(n12178), .CK(clk), .Q(
        weight_queue_6__2__7_), .QN(n1797) );
  DFF_X1 weight_queue_reg_6__2__6_ ( .D(n12171), .CK(clk), .Q(
        weight_queue_6__2__6_), .QN(n1798) );
  DFF_X1 weight_queue_reg_6__2__5_ ( .D(n12164), .CK(clk), .Q(
        weight_queue_6__2__5_), .QN(n1799) );
  DFF_X1 weight_queue_reg_6__2__4_ ( .D(n12157), .CK(clk), .Q(
        weight_queue_6__2__4_), .QN(n1800) );
  DFF_X1 weight_queue_reg_6__2__3_ ( .D(n12150), .CK(clk), .Q(
        weight_queue_6__2__3_), .QN(n1801) );
  DFF_X1 weight_queue_reg_6__2__2_ ( .D(n12143), .CK(clk), .Q(
        weight_queue_6__2__2_), .QN(n1802) );
  DFF_X1 weight_queue_reg_6__2__1_ ( .D(n12136), .CK(clk), .Q(
        weight_queue_6__2__1_), .QN(n1803) );
  DFF_X1 weight_queue_reg_6__2__0_ ( .D(n12129), .CK(clk), .Q(
        weight_queue_6__2__0_), .QN(n1804) );
  DFF_X1 weight_queue_reg_6__3__7_ ( .D(n12122), .CK(clk), .Q(
        weight_queue_6__3__7_), .QN(n1805) );
  DFF_X1 weight_queue_reg_6__3__6_ ( .D(n12115), .CK(clk), .Q(
        weight_queue_6__3__6_), .QN(n1806) );
  DFF_X1 weight_queue_reg_6__3__5_ ( .D(n12108), .CK(clk), .Q(
        weight_queue_6__3__5_), .QN(n1807) );
  DFF_X1 weight_queue_reg_6__3__4_ ( .D(n12101), .CK(clk), .Q(
        weight_queue_6__3__4_), .QN(n1808) );
  DFF_X1 weight_queue_reg_6__3__3_ ( .D(n12094), .CK(clk), .Q(
        weight_queue_6__3__3_), .QN(n1809) );
  DFF_X1 weight_queue_reg_6__3__2_ ( .D(n12087), .CK(clk), .Q(
        weight_queue_6__3__2_), .QN(n1810) );
  DFF_X1 weight_queue_reg_6__3__1_ ( .D(n12080), .CK(clk), .Q(
        weight_queue_6__3__1_), .QN(n1811) );
  DFF_X1 weight_queue_reg_6__3__0_ ( .D(n12073), .CK(clk), .Q(
        weight_queue_6__3__0_), .QN(n1812) );
  DFF_X1 weight_queue_reg_6__4__7_ ( .D(n12066), .CK(clk), .Q(
        weight_queue_6__4__7_), .QN(n1813) );
  DFF_X1 weight_queue_reg_6__4__6_ ( .D(n12059), .CK(clk), .Q(
        weight_queue_6__4__6_), .QN(n1814) );
  DFF_X1 weight_queue_reg_6__4__5_ ( .D(n12052), .CK(clk), .Q(
        weight_queue_6__4__5_), .QN(n1815) );
  DFF_X1 weight_queue_reg_6__4__4_ ( .D(n12045), .CK(clk), .Q(
        weight_queue_6__4__4_), .QN(n1816) );
  DFF_X1 weight_queue_reg_6__4__3_ ( .D(n12038), .CK(clk), .Q(
        weight_queue_6__4__3_), .QN(n1817) );
  DFF_X1 weight_queue_reg_6__4__2_ ( .D(n12031), .CK(clk), .Q(
        weight_queue_6__4__2_), .QN(n1818) );
  DFF_X1 weight_queue_reg_6__4__1_ ( .D(n12024), .CK(clk), .Q(
        weight_queue_6__4__1_), .QN(n1819) );
  DFF_X1 weight_queue_reg_6__4__0_ ( .D(n12017), .CK(clk), .Q(
        weight_queue_6__4__0_), .QN(n1820) );
  DFF_X1 weight_queue_reg_6__5__7_ ( .D(n12010), .CK(clk), .Q(
        weight_queue_6__5__7_), .QN(n1821) );
  DFF_X1 weight_queue_reg_6__5__6_ ( .D(n12003), .CK(clk), .Q(
        weight_queue_6__5__6_), .QN(n1822) );
  DFF_X1 weight_queue_reg_6__5__5_ ( .D(n11996), .CK(clk), .Q(
        weight_queue_6__5__5_), .QN(n1823) );
  DFF_X1 weight_queue_reg_6__5__4_ ( .D(n11989), .CK(clk), .Q(
        weight_queue_6__5__4_), .QN(n1824) );
  DFF_X1 weight_queue_reg_6__5__3_ ( .D(n11982), .CK(clk), .Q(
        weight_queue_6__5__3_), .QN(n1825) );
  DFF_X1 weight_queue_reg_6__5__2_ ( .D(n11975), .CK(clk), .Q(
        weight_queue_6__5__2_), .QN(n1826) );
  DFF_X1 weight_queue_reg_6__5__1_ ( .D(n11968), .CK(clk), .Q(
        weight_queue_6__5__1_), .QN(n1827) );
  DFF_X1 weight_queue_reg_6__5__0_ ( .D(n11961), .CK(clk), .Q(
        weight_queue_6__5__0_), .QN(n1828) );
  DFF_X1 weight_queue_reg_6__6__7_ ( .D(n11954), .CK(clk), .Q(
        weight_queue_6__6__7_), .QN(n1829) );
  DFF_X1 weight_queue_reg_6__6__6_ ( .D(n11947), .CK(clk), .Q(
        weight_queue_6__6__6_), .QN(n1830) );
  DFF_X1 weight_queue_reg_6__6__5_ ( .D(n11940), .CK(clk), .Q(
        weight_queue_6__6__5_), .QN(n1831) );
  DFF_X1 weight_queue_reg_6__6__4_ ( .D(n11933), .CK(clk), .Q(
        weight_queue_6__6__4_), .QN(n1832) );
  DFF_X1 weight_queue_reg_6__6__3_ ( .D(n11926), .CK(clk), .Q(
        weight_queue_6__6__3_), .QN(n1833) );
  DFF_X1 weight_queue_reg_6__6__2_ ( .D(n11919), .CK(clk), .Q(
        weight_queue_6__6__2_), .QN(n1834) );
  DFF_X1 weight_queue_reg_6__6__1_ ( .D(n11912), .CK(clk), .Q(
        weight_queue_6__6__1_), .QN(n1835) );
  DFF_X1 weight_queue_reg_6__6__0_ ( .D(n11905), .CK(clk), .Q(
        weight_queue_6__6__0_), .QN(n1836) );
  DFF_X1 weight_queue_reg_6__7__7_ ( .D(n11898), .CK(clk), .Q(
        weight_queue_6__7__7_), .QN(n1837) );
  DFF_X1 weight_queue_reg_6__7__6_ ( .D(n11891), .CK(clk), .Q(
        weight_queue_6__7__6_), .QN(n1838) );
  DFF_X1 weight_queue_reg_6__7__5_ ( .D(n11884), .CK(clk), .Q(
        weight_queue_6__7__5_), .QN(n1839) );
  DFF_X1 weight_queue_reg_6__7__4_ ( .D(n11877), .CK(clk), .Q(
        weight_queue_6__7__4_), .QN(n1840) );
  DFF_X1 weight_queue_reg_6__7__3_ ( .D(n11870), .CK(clk), .Q(
        weight_queue_6__7__3_), .QN(n1841) );
  DFF_X1 weight_queue_reg_6__7__2_ ( .D(n11863), .CK(clk), .Q(
        weight_queue_6__7__2_), .QN(n1842) );
  DFF_X1 weight_queue_reg_6__7__1_ ( .D(n11856), .CK(clk), .Q(
        weight_queue_6__7__1_), .QN(n1843) );
  DFF_X1 weight_queue_reg_6__7__0_ ( .D(n11849), .CK(clk), .Q(
        weight_queue_6__7__0_), .QN(n1844) );
  DFF_X1 weight_queue_reg_7__0__7_ ( .D(n11848), .CK(clk), .Q(
        weight_queue_7__0__7_), .QN(n17200) );
  DFF_X1 weight_queue_reg_7__0__6_ ( .D(n11845), .CK(clk), .Q(
        weight_queue_7__0__6_), .QN(n17199) );
  DFF_X1 weight_queue_reg_7__0__5_ ( .D(n11842), .CK(clk), .Q(
        weight_queue_7__0__5_), .QN(n17198) );
  DFF_X1 weight_queue_reg_7__0__4_ ( .D(n11839), .CK(clk), .Q(
        weight_queue_7__0__4_), .QN(n17197) );
  DFF_X1 weight_queue_reg_7__0__3_ ( .D(n11836), .CK(clk), .Q(
        weight_queue_7__0__3_), .QN(n17196) );
  DFF_X1 weight_queue_reg_7__0__2_ ( .D(n11833), .CK(clk), .Q(
        weight_queue_7__0__2_), .QN(n17195) );
  DFF_X1 weight_queue_reg_7__0__1_ ( .D(n11830), .CK(clk), .Q(
        weight_queue_7__0__1_), .QN(n17194) );
  DFF_X1 weight_queue_reg_7__0__0_ ( .D(n11827), .CK(clk), .Q(
        weight_queue_7__0__0_), .QN(n17193) );
  DFF_X1 weight_queue_reg_7__1__7_ ( .D(n11824), .CK(clk), .Q(
        weight_queue_7__1__7_), .QN(n17192) );
  DFF_X1 weight_queue_reg_7__1__6_ ( .D(n11821), .CK(clk), .Q(
        weight_queue_7__1__6_), .QN(n17191) );
  DFF_X1 weight_queue_reg_7__1__5_ ( .D(n11818), .CK(clk), .Q(
        weight_queue_7__1__5_), .QN(n17190) );
  DFF_X1 weight_queue_reg_7__1__4_ ( .D(n11815), .CK(clk), .Q(
        weight_queue_7__1__4_), .QN(n17189) );
  DFF_X1 weight_queue_reg_7__1__3_ ( .D(n11812), .CK(clk), .Q(
        weight_queue_7__1__3_), .QN(n17188) );
  DFF_X1 weight_queue_reg_7__1__2_ ( .D(n11809), .CK(clk), .Q(
        weight_queue_7__1__2_), .QN(n17187) );
  DFF_X1 weight_queue_reg_7__1__1_ ( .D(n11806), .CK(clk), .Q(
        weight_queue_7__1__1_), .QN(n17186) );
  DFF_X1 weight_queue_reg_7__1__0_ ( .D(n11803), .CK(clk), .Q(
        weight_queue_7__1__0_), .QN(n17185) );
  DFF_X1 weight_queue_reg_7__2__7_ ( .D(n11800), .CK(clk), .Q(
        weight_queue_7__2__7_), .QN(n17184) );
  DFF_X1 weight_queue_reg_7__2__6_ ( .D(n11797), .CK(clk), .Q(
        weight_queue_7__2__6_), .QN(n17183) );
  DFF_X1 weight_queue_reg_7__2__5_ ( .D(n11794), .CK(clk), .Q(
        weight_queue_7__2__5_), .QN(n17182) );
  DFF_X1 weight_queue_reg_7__2__4_ ( .D(n11791), .CK(clk), .Q(
        weight_queue_7__2__4_), .QN(n17181) );
  DFF_X1 weight_queue_reg_7__2__3_ ( .D(n11788), .CK(clk), .Q(
        weight_queue_7__2__3_), .QN(n17180) );
  DFF_X1 weight_queue_reg_7__2__2_ ( .D(n11785), .CK(clk), .Q(
        weight_queue_7__2__2_), .QN(n17179) );
  DFF_X1 weight_queue_reg_7__2__1_ ( .D(n11782), .CK(clk), .Q(
        weight_queue_7__2__1_), .QN(n17178) );
  DFF_X1 weight_queue_reg_7__2__0_ ( .D(n11779), .CK(clk), .Q(
        weight_queue_7__2__0_), .QN(n17177) );
  DFF_X1 weight_queue_reg_7__3__7_ ( .D(n11776), .CK(clk), .Q(
        weight_queue_7__3__7_), .QN(n17176) );
  DFF_X1 weight_queue_reg_7__3__6_ ( .D(n11773), .CK(clk), .Q(
        weight_queue_7__3__6_), .QN(n17175) );
  DFF_X1 weight_queue_reg_7__3__5_ ( .D(n11770), .CK(clk), .Q(
        weight_queue_7__3__5_), .QN(n17174) );
  DFF_X1 weight_queue_reg_7__3__4_ ( .D(n11767), .CK(clk), .Q(
        weight_queue_7__3__4_), .QN(n17173) );
  DFF_X1 weight_queue_reg_7__3__3_ ( .D(n11764), .CK(clk), .Q(
        weight_queue_7__3__3_), .QN(n17172) );
  DFF_X1 weight_queue_reg_7__3__2_ ( .D(n11761), .CK(clk), .Q(
        weight_queue_7__3__2_), .QN(n17171) );
  DFF_X1 weight_queue_reg_7__3__1_ ( .D(n11758), .CK(clk), .Q(
        weight_queue_7__3__1_), .QN(n17170) );
  DFF_X1 weight_queue_reg_7__3__0_ ( .D(n11755), .CK(clk), .Q(
        weight_queue_7__3__0_), .QN(n17169) );
  DFF_X1 weight_queue_reg_7__4__7_ ( .D(n11752), .CK(clk), .Q(
        weight_queue_7__4__7_), .QN(n17168) );
  DFF_X1 weight_queue_reg_7__4__6_ ( .D(n11749), .CK(clk), .Q(
        weight_queue_7__4__6_), .QN(n17167) );
  DFF_X1 weight_queue_reg_7__4__5_ ( .D(n11746), .CK(clk), .Q(
        weight_queue_7__4__5_), .QN(n17166) );
  DFF_X1 weight_queue_reg_7__4__4_ ( .D(n11743), .CK(clk), .Q(
        weight_queue_7__4__4_), .QN(n17165) );
  DFF_X1 weight_queue_reg_7__4__3_ ( .D(n11740), .CK(clk), .Q(
        weight_queue_7__4__3_), .QN(n17164) );
  DFF_X1 weight_queue_reg_7__4__2_ ( .D(n11737), .CK(clk), .Q(
        weight_queue_7__4__2_), .QN(n17163) );
  DFF_X1 weight_queue_reg_7__4__1_ ( .D(n11734), .CK(clk), .Q(
        weight_queue_7__4__1_), .QN(n17162) );
  DFF_X1 weight_queue_reg_7__4__0_ ( .D(n11731), .CK(clk), .Q(
        weight_queue_7__4__0_), .QN(n17161) );
  DFF_X1 weight_queue_reg_7__5__7_ ( .D(n11728), .CK(clk), .Q(
        weight_queue_7__5__7_), .QN(n17160) );
  DFF_X1 weight_queue_reg_7__5__6_ ( .D(n11725), .CK(clk), .Q(
        weight_queue_7__5__6_), .QN(n17159) );
  DFF_X1 weight_queue_reg_7__5__5_ ( .D(n11722), .CK(clk), .Q(
        weight_queue_7__5__5_), .QN(n17158) );
  DFF_X1 weight_queue_reg_7__5__4_ ( .D(n11719), .CK(clk), .Q(
        weight_queue_7__5__4_), .QN(n17157) );
  DFF_X1 weight_queue_reg_7__5__3_ ( .D(n11716), .CK(clk), .Q(
        weight_queue_7__5__3_), .QN(n17156) );
  DFF_X1 weight_queue_reg_7__5__2_ ( .D(n11713), .CK(clk), .Q(
        weight_queue_7__5__2_), .QN(n17155) );
  DFF_X1 weight_queue_reg_7__5__1_ ( .D(n11710), .CK(clk), .Q(
        weight_queue_7__5__1_), .QN(n17154) );
  DFF_X1 weight_queue_reg_7__5__0_ ( .D(n11707), .CK(clk), .Q(
        weight_queue_7__5__0_), .QN(n17153) );
  DFF_X1 weight_queue_reg_7__6__7_ ( .D(n11704), .CK(clk), .Q(
        weight_queue_7__6__7_), .QN(n17152) );
  DFF_X1 weight_queue_reg_7__6__6_ ( .D(n11701), .CK(clk), .Q(
        weight_queue_7__6__6_), .QN(n17151) );
  DFF_X1 weight_queue_reg_7__6__5_ ( .D(n11698), .CK(clk), .Q(
        weight_queue_7__6__5_), .QN(n17150) );
  DFF_X1 weight_queue_reg_7__6__4_ ( .D(n11695), .CK(clk), .Q(
        weight_queue_7__6__4_), .QN(n17149) );
  DFF_X1 weight_queue_reg_7__6__3_ ( .D(n11692), .CK(clk), .Q(
        weight_queue_7__6__3_), .QN(n17148) );
  DFF_X1 weight_queue_reg_7__6__2_ ( .D(n11689), .CK(clk), .Q(
        weight_queue_7__6__2_), .QN(n17147) );
  DFF_X1 weight_queue_reg_7__6__1_ ( .D(n11686), .CK(clk), .Q(
        weight_queue_7__6__1_), .QN(n17146) );
  DFF_X1 weight_queue_reg_7__6__0_ ( .D(n11683), .CK(clk), .Q(
        weight_queue_7__6__0_), .QN(n17145) );
  DFF_X1 weight_queue_reg_7__7__7_ ( .D(n11680), .CK(clk), .Q(
        weight_queue_7__7__7_), .QN(n17144) );
  DFF_X1 weight_queue_reg_7__7__6_ ( .D(n11677), .CK(clk), .Q(
        weight_queue_7__7__6_), .QN(n17143) );
  DFF_X1 weight_queue_reg_7__7__5_ ( .D(n11674), .CK(clk), .Q(
        weight_queue_7__7__5_), .QN(n17142) );
  DFF_X1 weight_queue_reg_7__7__4_ ( .D(n11671), .CK(clk), .Q(
        weight_queue_7__7__4_), .QN(n17141) );
  DFF_X1 weight_queue_reg_7__7__3_ ( .D(n11668), .CK(clk), .Q(
        weight_queue_7__7__3_), .QN(n17140) );
  DFF_X1 weight_queue_reg_7__7__2_ ( .D(n11665), .CK(clk), .Q(
        weight_queue_7__7__2_), .QN(n17139) );
  DFF_X1 weight_queue_reg_7__7__1_ ( .D(n11662), .CK(clk), .Q(
        weight_queue_7__7__1_), .QN(n17138) );
  DFF_X1 weight_queue_reg_7__7__0_ ( .D(n11659), .CK(clk), .Q(
        weight_queue_7__7__0_), .QN(n17137) );
  DFF_X1 matrix_mul_2D_reg_0__0__15_ ( .D(n11656), .CK(clk), .Q(
        matrix_mul_2D_0__0__15_), .QN(n17988) );
  DFF_X1 matrix_mul_2D_reg_0__0__16_ ( .D(n11655), .CK(clk), .Q(
        matrix_mul_2D_0__0__16_), .QN(n17986) );
  DFF_X1 matrix_mul_2D_reg_0__0__17_ ( .D(n11654), .CK(clk), .Q(
        matrix_mul_2D_0__0__17_), .QN(n17984) );
  DFF_X1 matrix_mul_2D_reg_0__0__18_ ( .D(n11653), .CK(clk), .Q(
        matrix_mul_2D_0__0__18_), .QN(n17982) );
  DFF_X1 matrix_mul_2D_reg_0__0__19_ ( .D(n11652), .CK(clk), .Q(
        matrix_mul_2D_0__0__19_), .QN(n17980) );
  DFF_X1 matrix_mul_2D_reg_0__0__20_ ( .D(n11651), .CK(clk), .Q(
        matrix_mul_2D_0__0__20_), .QN(n17978) );
  DFF_X1 matrix_mul_2D_reg_0__1__0_ ( .D(n11647), .CK(clk), .Q(
        matrix_mul_2D_0__1__0_), .QN(n1874) );
  DFF_X1 matrix_mul_2D_reg_0__1__1_ ( .D(n11642), .CK(clk), .Q(
        matrix_mul_2D_0__1__1_), .QN(n1873) );
  DFF_X1 matrix_mul_2D_reg_0__1__2_ ( .D(n11637), .CK(clk), .Q(
        matrix_mul_2D_0__1__2_), .QN(n1872) );
  DFF_X1 matrix_mul_2D_reg_0__1__3_ ( .D(n11632), .CK(clk), .Q(
        matrix_mul_2D_0__1__3_), .QN(n1871) );
  DFF_X1 matrix_mul_2D_reg_0__1__4_ ( .D(n11627), .CK(clk), .Q(
        matrix_mul_2D_0__1__4_), .QN(n1870) );
  DFF_X1 matrix_mul_2D_reg_0__1__5_ ( .D(n11622), .CK(clk), .Q(
        matrix_mul_2D_0__1__5_), .QN(n1869) );
  DFF_X1 matrix_mul_2D_reg_0__1__6_ ( .D(n11617), .CK(clk), .Q(
        matrix_mul_2D_0__1__6_), .QN(n1868) );
  DFF_X1 matrix_mul_2D_reg_0__1__7_ ( .D(n11612), .CK(clk), .Q(
        matrix_mul_2D_0__1__7_), .QN(n1867) );
  DFF_X1 matrix_mul_2D_reg_0__1__8_ ( .D(n11607), .CK(clk), .Q(
        matrix_mul_2D_0__1__8_), .QN(n1866) );
  DFF_X1 matrix_mul_2D_reg_0__1__9_ ( .D(n11602), .CK(clk), .Q(
        matrix_mul_2D_0__1__9_), .QN(n1865) );
  DFF_X1 matrix_mul_2D_reg_0__1__10_ ( .D(n11597), .CK(clk), .Q(
        matrix_mul_2D_0__1__10_), .QN(n1864) );
  DFF_X1 matrix_mul_2D_reg_0__1__11_ ( .D(n11592), .CK(clk), .Q(
        matrix_mul_2D_0__1__11_), .QN(n1863) );
  DFF_X1 matrix_mul_2D_reg_0__1__12_ ( .D(n11587), .CK(clk), .Q(
        matrix_mul_2D_0__1__12_), .QN(n1862) );
  DFF_X1 matrix_mul_2D_reg_0__1__13_ ( .D(n11582), .CK(clk), .Q(
        matrix_mul_2D_0__1__13_), .QN(n1861) );
  DFF_X1 matrix_mul_2D_reg_0__1__14_ ( .D(n11577), .CK(clk), .Q(
        matrix_mul_2D_0__1__14_), .QN(n1860) );
  DFF_X1 matrix_mul_2D_reg_0__1__15_ ( .D(n11576), .CK(clk), .Q(
        matrix_mul_2D_0__1__15_), .QN(n17976) );
  DFF_X1 matrix_mul_2D_reg_0__1__16_ ( .D(n11575), .CK(clk), .Q(
        matrix_mul_2D_0__1__16_), .QN(n17974) );
  DFF_X1 matrix_mul_2D_reg_0__1__17_ ( .D(n11574), .CK(clk), .Q(
        matrix_mul_2D_0__1__17_), .QN(n17972) );
  DFF_X1 matrix_mul_2D_reg_0__1__18_ ( .D(n11573), .CK(clk), .Q(
        matrix_mul_2D_0__1__18_), .QN(n17970) );
  DFF_X1 matrix_mul_2D_reg_0__1__19_ ( .D(n11572), .CK(clk), .Q(
        matrix_mul_2D_0__1__19_), .QN(n17968) );
  DFF_X1 matrix_mul_2D_reg_0__1__20_ ( .D(n11571), .CK(clk), .Q(
        matrix_mul_2D_0__1__20_), .QN(n17966) );
  DFF_X1 matrix_mul_2D_reg_0__2__0_ ( .D(n11567), .CK(clk), .Q(
        matrix_mul_2D_0__2__0_), .QN(n1889) );
  DFF_X1 matrix_mul_2D_reg_0__2__1_ ( .D(n11562), .CK(clk), .Q(
        matrix_mul_2D_0__2__1_), .QN(n1888) );
  DFF_X1 matrix_mul_2D_reg_0__2__2_ ( .D(n11557), .CK(clk), .Q(
        matrix_mul_2D_0__2__2_), .QN(n1887) );
  DFF_X1 matrix_mul_2D_reg_0__2__3_ ( .D(n11552), .CK(clk), .Q(
        matrix_mul_2D_0__2__3_), .QN(n1886) );
  DFF_X1 matrix_mul_2D_reg_0__2__4_ ( .D(n11547), .CK(clk), .Q(
        matrix_mul_2D_0__2__4_), .QN(n1885) );
  DFF_X1 matrix_mul_2D_reg_0__2__5_ ( .D(n11542), .CK(clk), .Q(
        matrix_mul_2D_0__2__5_), .QN(n1884) );
  DFF_X1 matrix_mul_2D_reg_0__2__6_ ( .D(n11537), .CK(clk), .Q(
        matrix_mul_2D_0__2__6_), .QN(n1883) );
  DFF_X1 matrix_mul_2D_reg_0__2__7_ ( .D(n11532), .CK(clk), .Q(
        matrix_mul_2D_0__2__7_), .QN(n1882) );
  DFF_X1 matrix_mul_2D_reg_0__2__8_ ( .D(n11527), .CK(clk), .Q(
        matrix_mul_2D_0__2__8_), .QN(n1881) );
  DFF_X1 matrix_mul_2D_reg_0__2__9_ ( .D(n11522), .CK(clk), .Q(
        matrix_mul_2D_0__2__9_), .QN(n1880) );
  DFF_X1 matrix_mul_2D_reg_0__2__10_ ( .D(n11517), .CK(clk), .Q(
        matrix_mul_2D_0__2__10_), .QN(n1879) );
  DFF_X1 matrix_mul_2D_reg_0__2__11_ ( .D(n11512), .CK(clk), .Q(
        matrix_mul_2D_0__2__11_), .QN(n1878) );
  DFF_X1 matrix_mul_2D_reg_0__2__12_ ( .D(n11507), .CK(clk), .Q(
        matrix_mul_2D_0__2__12_), .QN(n1877) );
  DFF_X1 matrix_mul_2D_reg_0__2__13_ ( .D(n11502), .CK(clk), .Q(
        matrix_mul_2D_0__2__13_), .QN(n1876) );
  DFF_X1 matrix_mul_2D_reg_0__2__14_ ( .D(n11497), .CK(clk), .Q(
        matrix_mul_2D_0__2__14_), .QN(n1875) );
  DFF_X1 matrix_mul_2D_reg_0__2__15_ ( .D(n11496), .CK(clk), .Q(
        matrix_mul_2D_0__2__15_), .QN(n17964) );
  DFF_X1 matrix_mul_2D_reg_0__2__16_ ( .D(n11495), .CK(clk), .Q(
        matrix_mul_2D_0__2__16_), .QN(n17962) );
  DFF_X1 matrix_mul_2D_reg_0__2__17_ ( .D(n11494), .CK(clk), .Q(
        matrix_mul_2D_0__2__17_), .QN(n17960) );
  DFF_X1 matrix_mul_2D_reg_0__2__18_ ( .D(n11493), .CK(clk), .Q(
        matrix_mul_2D_0__2__18_), .QN(n17958) );
  DFF_X1 matrix_mul_2D_reg_0__2__19_ ( .D(n11492), .CK(clk), .Q(
        matrix_mul_2D_0__2__19_), .QN(n17956) );
  DFF_X1 matrix_mul_2D_reg_0__2__20_ ( .D(n11491), .CK(clk), .Q(
        matrix_mul_2D_0__2__20_), .QN(n17954) );
  DFF_X1 matrix_mul_2D_reg_0__3__0_ ( .D(n11487), .CK(clk), .Q(
        matrix_mul_2D_0__3__0_), .QN(n1904) );
  DFF_X1 matrix_mul_2D_reg_0__3__1_ ( .D(n11482), .CK(clk), .Q(
        matrix_mul_2D_0__3__1_), .QN(n1903) );
  DFF_X1 matrix_mul_2D_reg_0__3__2_ ( .D(n11477), .CK(clk), .Q(
        matrix_mul_2D_0__3__2_), .QN(n1902) );
  DFF_X1 matrix_mul_2D_reg_0__3__3_ ( .D(n11472), .CK(clk), .Q(
        matrix_mul_2D_0__3__3_), .QN(n1901) );
  DFF_X1 matrix_mul_2D_reg_0__3__4_ ( .D(n11467), .CK(clk), .Q(
        matrix_mul_2D_0__3__4_), .QN(n1900) );
  DFF_X1 matrix_mul_2D_reg_0__3__5_ ( .D(n11462), .CK(clk), .Q(
        matrix_mul_2D_0__3__5_), .QN(n1899) );
  DFF_X1 matrix_mul_2D_reg_0__3__6_ ( .D(n11457), .CK(clk), .Q(
        matrix_mul_2D_0__3__6_), .QN(n1898) );
  DFF_X1 matrix_mul_2D_reg_0__3__7_ ( .D(n11452), .CK(clk), .Q(
        matrix_mul_2D_0__3__7_), .QN(n1897) );
  DFF_X1 matrix_mul_2D_reg_0__3__8_ ( .D(n11447), .CK(clk), .Q(
        matrix_mul_2D_0__3__8_), .QN(n1896) );
  DFF_X1 matrix_mul_2D_reg_0__3__9_ ( .D(n11442), .CK(clk), .Q(
        matrix_mul_2D_0__3__9_), .QN(n1895) );
  DFF_X1 matrix_mul_2D_reg_0__3__10_ ( .D(n11437), .CK(clk), .Q(
        matrix_mul_2D_0__3__10_), .QN(n1894) );
  DFF_X1 matrix_mul_2D_reg_0__3__11_ ( .D(n11432), .CK(clk), .Q(
        matrix_mul_2D_0__3__11_), .QN(n1893) );
  DFF_X1 matrix_mul_2D_reg_0__3__12_ ( .D(n11427), .CK(clk), .Q(
        matrix_mul_2D_0__3__12_), .QN(n1892) );
  DFF_X1 matrix_mul_2D_reg_0__3__13_ ( .D(n11422), .CK(clk), .Q(
        matrix_mul_2D_0__3__13_), .QN(n1891) );
  DFF_X1 matrix_mul_2D_reg_0__3__14_ ( .D(n11417), .CK(clk), .Q(
        matrix_mul_2D_0__3__14_), .QN(n1890) );
  DFF_X1 matrix_mul_2D_reg_0__3__15_ ( .D(n11416), .CK(clk), .Q(
        matrix_mul_2D_0__3__15_), .QN(n17952) );
  DFF_X1 matrix_mul_2D_reg_0__3__16_ ( .D(n11415), .CK(clk), .Q(
        matrix_mul_2D_0__3__16_), .QN(n17950) );
  DFF_X1 matrix_mul_2D_reg_0__3__17_ ( .D(n11414), .CK(clk), .Q(
        matrix_mul_2D_0__3__17_), .QN(n17948) );
  DFF_X1 matrix_mul_2D_reg_0__3__18_ ( .D(n11413), .CK(clk), .Q(
        matrix_mul_2D_0__3__18_), .QN(n17946) );
  DFF_X1 matrix_mul_2D_reg_0__3__19_ ( .D(n11412), .CK(clk), .Q(
        matrix_mul_2D_0__3__19_), .QN(n17944) );
  DFF_X1 matrix_mul_2D_reg_0__3__20_ ( .D(n11411), .CK(clk), .Q(
        matrix_mul_2D_0__3__20_), .QN(n17942) );
  DFF_X1 matrix_mul_2D_reg_0__4__0_ ( .D(n11407), .CK(clk), .Q(
        matrix_mul_2D_0__4__0_), .QN(n1919) );
  DFF_X1 matrix_mul_2D_reg_0__4__1_ ( .D(n11402), .CK(clk), .Q(
        matrix_mul_2D_0__4__1_), .QN(n1918) );
  DFF_X1 matrix_mul_2D_reg_0__4__2_ ( .D(n11397), .CK(clk), .Q(
        matrix_mul_2D_0__4__2_), .QN(n1917) );
  DFF_X1 matrix_mul_2D_reg_0__4__3_ ( .D(n11392), .CK(clk), .Q(
        matrix_mul_2D_0__4__3_), .QN(n1916) );
  DFF_X1 matrix_mul_2D_reg_0__4__4_ ( .D(n11387), .CK(clk), .Q(
        matrix_mul_2D_0__4__4_), .QN(n1915) );
  DFF_X1 matrix_mul_2D_reg_0__4__5_ ( .D(n11382), .CK(clk), .Q(
        matrix_mul_2D_0__4__5_), .QN(n1914) );
  DFF_X1 matrix_mul_2D_reg_0__4__6_ ( .D(n11377), .CK(clk), .Q(
        matrix_mul_2D_0__4__6_), .QN(n1913) );
  DFF_X1 matrix_mul_2D_reg_0__4__7_ ( .D(n11372), .CK(clk), .Q(
        matrix_mul_2D_0__4__7_), .QN(n1912) );
  DFF_X1 matrix_mul_2D_reg_0__4__8_ ( .D(n11367), .CK(clk), .Q(
        matrix_mul_2D_0__4__8_), .QN(n1911) );
  DFF_X1 matrix_mul_2D_reg_0__4__9_ ( .D(n11362), .CK(clk), .Q(
        matrix_mul_2D_0__4__9_), .QN(n1910) );
  DFF_X1 matrix_mul_2D_reg_0__4__10_ ( .D(n11357), .CK(clk), .Q(
        matrix_mul_2D_0__4__10_), .QN(n1909) );
  DFF_X1 matrix_mul_2D_reg_0__4__11_ ( .D(n11352), .CK(clk), .Q(
        matrix_mul_2D_0__4__11_), .QN(n1908) );
  DFF_X1 matrix_mul_2D_reg_0__4__12_ ( .D(n11347), .CK(clk), .Q(
        matrix_mul_2D_0__4__12_), .QN(n1907) );
  DFF_X1 matrix_mul_2D_reg_0__4__13_ ( .D(n11342), .CK(clk), .Q(
        matrix_mul_2D_0__4__13_), .QN(n1906) );
  DFF_X1 matrix_mul_2D_reg_0__4__14_ ( .D(n11337), .CK(clk), .Q(
        matrix_mul_2D_0__4__14_), .QN(n1905) );
  DFF_X1 matrix_mul_2D_reg_0__4__15_ ( .D(n11336), .CK(clk), .Q(
        matrix_mul_2D_0__4__15_), .QN(n17940) );
  DFF_X1 matrix_mul_2D_reg_0__4__16_ ( .D(n11335), .CK(clk), .Q(
        matrix_mul_2D_0__4__16_), .QN(n17938) );
  DFF_X1 matrix_mul_2D_reg_0__4__17_ ( .D(n11334), .CK(clk), .Q(
        matrix_mul_2D_0__4__17_), .QN(n17936) );
  DFF_X1 matrix_mul_2D_reg_0__4__18_ ( .D(n11333), .CK(clk), .Q(
        matrix_mul_2D_0__4__18_), .QN(n17934) );
  DFF_X1 matrix_mul_2D_reg_0__4__19_ ( .D(n11332), .CK(clk), .Q(
        matrix_mul_2D_0__4__19_), .QN(n17932) );
  DFF_X1 matrix_mul_2D_reg_0__4__20_ ( .D(n11331), .CK(clk), .Q(
        matrix_mul_2D_0__4__20_), .QN(n17930) );
  DFF_X1 matrix_mul_2D_reg_0__5__0_ ( .D(n11326), .CK(clk), .Q(
        matrix_mul_2D_0__5__0_), .QN(n1940) );
  DFF_X1 matrix_mul_2D_reg_0__5__1_ ( .D(n11322), .CK(clk), .Q(
        matrix_mul_2D_0__5__1_), .QN(n1939) );
  DFF_X1 matrix_mul_2D_reg_0__5__2_ ( .D(n11318), .CK(clk), .Q(
        matrix_mul_2D_0__5__2_), .QN(n1938) );
  DFF_X1 matrix_mul_2D_reg_0__5__3_ ( .D(n11314), .CK(clk), .Q(
        matrix_mul_2D_0__5__3_), .QN(n1937) );
  DFF_X1 matrix_mul_2D_reg_0__5__4_ ( .D(n11310), .CK(clk), .Q(
        matrix_mul_2D_0__5__4_), .QN(n1936) );
  DFF_X1 matrix_mul_2D_reg_0__5__5_ ( .D(n11306), .CK(clk), .Q(
        matrix_mul_2D_0__5__5_), .QN(n1935) );
  DFF_X1 matrix_mul_2D_reg_0__5__6_ ( .D(n11302), .CK(clk), .Q(
        matrix_mul_2D_0__5__6_), .QN(n1934) );
  DFF_X1 matrix_mul_2D_reg_0__5__7_ ( .D(n11298), .CK(clk), .Q(
        matrix_mul_2D_0__5__7_), .QN(n1933) );
  DFF_X1 matrix_mul_2D_reg_0__5__8_ ( .D(n11294), .CK(clk), .Q(
        matrix_mul_2D_0__5__8_), .QN(n1932) );
  DFF_X1 matrix_mul_2D_reg_0__5__9_ ( .D(n11290), .CK(clk), .Q(
        matrix_mul_2D_0__5__9_), .QN(n1931) );
  DFF_X1 matrix_mul_2D_reg_0__5__10_ ( .D(n11286), .CK(clk), .Q(
        matrix_mul_2D_0__5__10_), .QN(n1930) );
  DFF_X1 matrix_mul_2D_reg_0__5__11_ ( .D(n11282), .CK(clk), .Q(
        matrix_mul_2D_0__5__11_), .QN(n1929) );
  DFF_X1 matrix_mul_2D_reg_0__5__12_ ( .D(n11278), .CK(clk), .Q(
        matrix_mul_2D_0__5__12_), .QN(n1928) );
  DFF_X1 matrix_mul_2D_reg_0__5__13_ ( .D(n11274), .CK(clk), .Q(
        matrix_mul_2D_0__5__13_), .QN(n1927) );
  DFF_X1 matrix_mul_2D_reg_0__5__14_ ( .D(n11270), .CK(clk), .Q(
        matrix_mul_2D_0__5__14_), .QN(n1926) );
  DFF_X1 matrix_mul_2D_reg_0__5__15_ ( .D(n11269), .CK(clk), .Q(
        matrix_mul_2D_0__5__15_), .QN(n17928) );
  DFF_X1 matrix_mul_2D_reg_0__5__16_ ( .D(n11268), .CK(clk), .Q(
        matrix_mul_2D_0__5__16_), .QN(n17926) );
  DFF_X1 matrix_mul_2D_reg_0__5__17_ ( .D(n11267), .CK(clk), .Q(
        matrix_mul_2D_0__5__17_), .QN(n17924) );
  DFF_X1 matrix_mul_2D_reg_0__5__18_ ( .D(n11266), .CK(clk), .Q(
        matrix_mul_2D_0__5__18_), .QN(n17922) );
  DFF_X1 matrix_mul_2D_reg_0__5__19_ ( .D(n11265), .CK(clk), .Q(
        matrix_mul_2D_0__5__19_), .QN(n17920) );
  DFF_X1 matrix_mul_2D_reg_0__5__20_ ( .D(n11264), .CK(clk), .Q(
        matrix_mul_2D_0__5__20_), .QN(n17918) );
  DFF_X1 matrix_mul_2D_reg_0__6__0_ ( .D(n11260), .CK(clk), .Q(
        matrix_mul_2D_0__6__0_), .QN(n1955) );
  DFF_X1 matrix_mul_2D_reg_0__6__1_ ( .D(n11255), .CK(clk), .Q(
        matrix_mul_2D_0__6__1_), .QN(n1954) );
  DFF_X1 matrix_mul_2D_reg_0__6__2_ ( .D(n11250), .CK(clk), .Q(
        matrix_mul_2D_0__6__2_), .QN(n1953) );
  DFF_X1 matrix_mul_2D_reg_0__6__3_ ( .D(n11245), .CK(clk), .Q(
        matrix_mul_2D_0__6__3_), .QN(n1952) );
  DFF_X1 matrix_mul_2D_reg_0__6__4_ ( .D(n11240), .CK(clk), .Q(
        matrix_mul_2D_0__6__4_), .QN(n1951) );
  DFF_X1 matrix_mul_2D_reg_0__6__5_ ( .D(n11235), .CK(clk), .Q(
        matrix_mul_2D_0__6__5_), .QN(n1950) );
  DFF_X1 matrix_mul_2D_reg_0__6__6_ ( .D(n11230), .CK(clk), .Q(
        matrix_mul_2D_0__6__6_), .QN(n1949) );
  DFF_X1 matrix_mul_2D_reg_0__6__7_ ( .D(n11225), .CK(clk), .Q(
        matrix_mul_2D_0__6__7_), .QN(n1948) );
  DFF_X1 matrix_mul_2D_reg_0__6__8_ ( .D(n11220), .CK(clk), .Q(
        matrix_mul_2D_0__6__8_), .QN(n1947) );
  DFF_X1 matrix_mul_2D_reg_0__6__9_ ( .D(n11215), .CK(clk), .Q(
        matrix_mul_2D_0__6__9_), .QN(n1946) );
  DFF_X1 matrix_mul_2D_reg_0__6__10_ ( .D(n11210), .CK(clk), .Q(
        matrix_mul_2D_0__6__10_), .QN(n1945) );
  DFF_X1 matrix_mul_2D_reg_0__6__11_ ( .D(n11205), .CK(clk), .Q(
        matrix_mul_2D_0__6__11_), .QN(n1944) );
  DFF_X1 matrix_mul_2D_reg_0__6__12_ ( .D(n11200), .CK(clk), .Q(
        matrix_mul_2D_0__6__12_), .QN(n1943) );
  DFF_X1 matrix_mul_2D_reg_0__6__13_ ( .D(n11195), .CK(clk), .Q(
        matrix_mul_2D_0__6__13_), .QN(n1942) );
  DFF_X1 matrix_mul_2D_reg_0__6__14_ ( .D(n11190), .CK(clk), .Q(
        matrix_mul_2D_0__6__14_), .QN(n1941) );
  DFF_X1 matrix_mul_2D_reg_0__6__15_ ( .D(n11189), .CK(clk), .Q(
        matrix_mul_2D_0__6__15_), .QN(n17916) );
  DFF_X1 matrix_mul_2D_reg_0__6__16_ ( .D(n11188), .CK(clk), .Q(
        matrix_mul_2D_0__6__16_), .QN(n17914) );
  DFF_X1 matrix_mul_2D_reg_0__6__17_ ( .D(n11187), .CK(clk), .Q(
        matrix_mul_2D_0__6__17_), .QN(n17912) );
  DFF_X1 matrix_mul_2D_reg_0__6__18_ ( .D(n11186), .CK(clk), .Q(
        matrix_mul_2D_0__6__18_), .QN(n17910) );
  DFF_X1 matrix_mul_2D_reg_0__6__19_ ( .D(n11185), .CK(clk), .Q(
        matrix_mul_2D_0__6__19_), .QN(n17908) );
  DFF_X1 matrix_mul_2D_reg_0__6__20_ ( .D(n11184), .CK(clk), .Q(
        matrix_mul_2D_0__6__20_), .QN(n17906) );
  DFF_X1 matrix_mul_2D_reg_0__7__0_ ( .D(n11179), .CK(clk), .Q(
        matrix_mul_2D_0__7__0_), .QN(n1970) );
  DFF_X1 matrix_mul_2D_reg_0__7__1_ ( .D(n11175), .CK(clk), .Q(
        matrix_mul_2D_0__7__1_), .QN(n1969) );
  DFF_X1 matrix_mul_2D_reg_0__7__2_ ( .D(n11171), .CK(clk), .Q(
        matrix_mul_2D_0__7__2_), .QN(n1968) );
  DFF_X1 matrix_mul_2D_reg_0__7__3_ ( .D(n11167), .CK(clk), .Q(
        matrix_mul_2D_0__7__3_), .QN(n1967) );
  DFF_X1 matrix_mul_2D_reg_0__7__4_ ( .D(n11163), .CK(clk), .Q(
        matrix_mul_2D_0__7__4_), .QN(n1966) );
  DFF_X1 matrix_mul_2D_reg_0__7__5_ ( .D(n11159), .CK(clk), .Q(
        matrix_mul_2D_0__7__5_), .QN(n1965) );
  DFF_X1 matrix_mul_2D_reg_0__7__6_ ( .D(n11155), .CK(clk), .Q(
        matrix_mul_2D_0__7__6_), .QN(n1964) );
  DFF_X1 matrix_mul_2D_reg_0__7__7_ ( .D(n11151), .CK(clk), .Q(
        matrix_mul_2D_0__7__7_), .QN(n1963) );
  DFF_X1 matrix_mul_2D_reg_0__7__8_ ( .D(n11147), .CK(clk), .Q(
        matrix_mul_2D_0__7__8_), .QN(n1962) );
  DFF_X1 matrix_mul_2D_reg_0__7__9_ ( .D(n11143), .CK(clk), .Q(
        matrix_mul_2D_0__7__9_), .QN(n1961) );
  DFF_X1 matrix_mul_2D_reg_0__7__10_ ( .D(n11139), .CK(clk), .Q(
        matrix_mul_2D_0__7__10_), .QN(n1960) );
  DFF_X1 matrix_mul_2D_reg_0__7__11_ ( .D(n11135), .CK(clk), .Q(
        matrix_mul_2D_0__7__11_), .QN(n1959) );
  DFF_X1 matrix_mul_2D_reg_0__7__12_ ( .D(n11131), .CK(clk), .Q(
        matrix_mul_2D_0__7__12_), .QN(n1958) );
  DFF_X1 matrix_mul_2D_reg_0__7__13_ ( .D(n11127), .CK(clk), .Q(
        matrix_mul_2D_0__7__13_), .QN(n1957) );
  DFF_X1 matrix_mul_2D_reg_0__7__14_ ( .D(n11123), .CK(clk), .Q(
        matrix_mul_2D_0__7__14_), .QN(n1956) );
  DFF_X1 matrix_mul_2D_reg_0__7__15_ ( .D(n11122), .CK(clk), .Q(
        matrix_mul_2D_0__7__15_), .QN(n17904) );
  DFF_X1 matrix_mul_2D_reg_0__7__16_ ( .D(n11121), .CK(clk), .Q(
        matrix_mul_2D_0__7__16_), .QN(n17902) );
  DFF_X1 matrix_mul_2D_reg_0__7__17_ ( .D(n11120), .CK(clk), .Q(
        matrix_mul_2D_0__7__17_), .QN(n17900) );
  DFF_X1 matrix_mul_2D_reg_0__7__18_ ( .D(n11119), .CK(clk), .Q(
        matrix_mul_2D_0__7__18_), .QN(n17898) );
  DFF_X1 matrix_mul_2D_reg_0__7__19_ ( .D(n11118), .CK(clk), .Q(
        matrix_mul_2D_0__7__19_), .QN(n17896) );
  DFF_X1 matrix_mul_2D_reg_0__7__20_ ( .D(n11117), .CK(clk), .Q(
        matrix_mul_2D_0__7__20_), .QN(n17894) );
  DFF_X1 matrix_mul_2D_reg_1__0__0_ ( .D(n11113), .CK(clk), .Q(
        matrix_mul_2D_1__0__0_), .QN(n1985) );
  DFF_X1 matrix_mul_2D_reg_1__0__1_ ( .D(n11108), .CK(clk), .Q(
        matrix_mul_2D_1__0__1_), .QN(n1984) );
  DFF_X1 matrix_mul_2D_reg_1__0__2_ ( .D(n11103), .CK(clk), .Q(
        matrix_mul_2D_1__0__2_), .QN(n1983) );
  DFF_X1 matrix_mul_2D_reg_1__0__3_ ( .D(n11098), .CK(clk), .Q(
        matrix_mul_2D_1__0__3_), .QN(n1982) );
  DFF_X1 matrix_mul_2D_reg_1__0__4_ ( .D(n11093), .CK(clk), .Q(
        matrix_mul_2D_1__0__4_), .QN(n1981) );
  DFF_X1 matrix_mul_2D_reg_1__0__5_ ( .D(n11088), .CK(clk), .Q(
        matrix_mul_2D_1__0__5_), .QN(n1980) );
  DFF_X1 matrix_mul_2D_reg_1__0__6_ ( .D(n11083), .CK(clk), .Q(
        matrix_mul_2D_1__0__6_), .QN(n1979) );
  DFF_X1 matrix_mul_2D_reg_1__0__7_ ( .D(n11078), .CK(clk), .Q(
        matrix_mul_2D_1__0__7_), .QN(n1978) );
  DFF_X1 matrix_mul_2D_reg_1__0__8_ ( .D(n11073), .CK(clk), .Q(
        matrix_mul_2D_1__0__8_), .QN(n1977) );
  DFF_X1 matrix_mul_2D_reg_1__0__9_ ( .D(n11068), .CK(clk), .Q(
        matrix_mul_2D_1__0__9_), .QN(n1976) );
  DFF_X1 matrix_mul_2D_reg_1__0__10_ ( .D(n11063), .CK(clk), .Q(
        matrix_mul_2D_1__0__10_), .QN(n1975) );
  DFF_X1 matrix_mul_2D_reg_1__0__11_ ( .D(n11058), .CK(clk), .Q(
        matrix_mul_2D_1__0__11_), .QN(n1974) );
  DFF_X1 matrix_mul_2D_reg_1__0__12_ ( .D(n11053), .CK(clk), .Q(
        matrix_mul_2D_1__0__12_), .QN(n1973) );
  DFF_X1 matrix_mul_2D_reg_1__0__13_ ( .D(n11048), .CK(clk), .Q(
        matrix_mul_2D_1__0__13_), .QN(n1972) );
  DFF_X1 matrix_mul_2D_reg_1__0__14_ ( .D(n11043), .CK(clk), .Q(
        matrix_mul_2D_1__0__14_), .QN(n1971) );
  DFF_X1 matrix_mul_2D_reg_1__0__15_ ( .D(n11042), .CK(clk), .Q(
        matrix_mul_2D_1__0__15_), .QN(n17892) );
  DFF_X1 matrix_mul_2D_reg_1__0__16_ ( .D(n11041), .CK(clk), .Q(
        matrix_mul_2D_1__0__16_), .QN(n17890) );
  DFF_X1 matrix_mul_2D_reg_1__0__17_ ( .D(n11040), .CK(clk), .Q(
        matrix_mul_2D_1__0__17_), .QN(n17888) );
  DFF_X1 matrix_mul_2D_reg_1__0__18_ ( .D(n11039), .CK(clk), .Q(
        matrix_mul_2D_1__0__18_), .QN(n17886) );
  DFF_X1 matrix_mul_2D_reg_1__0__19_ ( .D(n11038), .CK(clk), .Q(
        matrix_mul_2D_1__0__19_), .QN(n17884) );
  DFF_X1 matrix_mul_2D_reg_1__0__20_ ( .D(n11037), .CK(clk), .Q(
        matrix_mul_2D_1__0__20_), .QN(n17882) );
  DFF_X1 matrix_mul_2D_reg_1__1__0_ ( .D(n11033), .CK(clk), .Q(
        matrix_mul_2D_1__1__0_), .QN(n2000) );
  DFF_X1 matrix_mul_2D_reg_1__1__1_ ( .D(n11028), .CK(clk), .Q(
        matrix_mul_2D_1__1__1_), .QN(n1999) );
  DFF_X1 matrix_mul_2D_reg_1__1__2_ ( .D(n11023), .CK(clk), .Q(
        matrix_mul_2D_1__1__2_), .QN(n1998) );
  DFF_X1 matrix_mul_2D_reg_1__1__3_ ( .D(n11018), .CK(clk), .Q(
        matrix_mul_2D_1__1__3_), .QN(n1997) );
  DFF_X1 matrix_mul_2D_reg_1__1__4_ ( .D(n11013), .CK(clk), .Q(
        matrix_mul_2D_1__1__4_), .QN(n1996) );
  DFF_X1 matrix_mul_2D_reg_1__1__5_ ( .D(n11008), .CK(clk), .Q(
        matrix_mul_2D_1__1__5_), .QN(n1995) );
  DFF_X1 matrix_mul_2D_reg_1__1__6_ ( .D(n11003), .CK(clk), .Q(
        matrix_mul_2D_1__1__6_), .QN(n1994) );
  DFF_X1 matrix_mul_2D_reg_1__1__7_ ( .D(n10998), .CK(clk), .Q(
        matrix_mul_2D_1__1__7_), .QN(n1993) );
  DFF_X1 matrix_mul_2D_reg_1__1__8_ ( .D(n10993), .CK(clk), .Q(
        matrix_mul_2D_1__1__8_), .QN(n1992) );
  DFF_X1 matrix_mul_2D_reg_1__1__9_ ( .D(n10988), .CK(clk), .Q(
        matrix_mul_2D_1__1__9_), .QN(n1991) );
  DFF_X1 matrix_mul_2D_reg_1__1__10_ ( .D(n10983), .CK(clk), .Q(
        matrix_mul_2D_1__1__10_), .QN(n1990) );
  DFF_X1 matrix_mul_2D_reg_1__1__11_ ( .D(n10978), .CK(clk), .Q(
        matrix_mul_2D_1__1__11_), .QN(n1989) );
  DFF_X1 matrix_mul_2D_reg_1__1__12_ ( .D(n10973), .CK(clk), .Q(
        matrix_mul_2D_1__1__12_), .QN(n1988) );
  DFF_X1 matrix_mul_2D_reg_1__1__13_ ( .D(n10968), .CK(clk), .Q(
        matrix_mul_2D_1__1__13_), .QN(n1987) );
  DFF_X1 matrix_mul_2D_reg_1__1__14_ ( .D(n10963), .CK(clk), .Q(
        matrix_mul_2D_1__1__14_), .QN(n1986) );
  DFF_X1 matrix_mul_2D_reg_1__1__15_ ( .D(n10962), .CK(clk), .Q(
        matrix_mul_2D_1__1__15_), .QN(n17880) );
  DFF_X1 matrix_mul_2D_reg_1__1__16_ ( .D(n10961), .CK(clk), .Q(
        matrix_mul_2D_1__1__16_), .QN(n17878) );
  DFF_X1 matrix_mul_2D_reg_1__1__17_ ( .D(n10960), .CK(clk), .Q(
        matrix_mul_2D_1__1__17_), .QN(n17876) );
  DFF_X1 matrix_mul_2D_reg_1__1__18_ ( .D(n10959), .CK(clk), .Q(
        matrix_mul_2D_1__1__18_), .QN(n17874) );
  DFF_X1 matrix_mul_2D_reg_1__1__19_ ( .D(n10958), .CK(clk), .Q(
        matrix_mul_2D_1__1__19_), .QN(n17872) );
  DFF_X1 matrix_mul_2D_reg_1__1__20_ ( .D(n10957), .CK(clk), .Q(
        matrix_mul_2D_1__1__20_), .QN(n17870) );
  DFF_X1 matrix_mul_2D_reg_1__2__0_ ( .D(n10952), .CK(clk), .Q(
        matrix_mul_2D_1__2__0_), .QN(n2021) );
  DFF_X1 matrix_mul_2D_reg_1__2__1_ ( .D(n10948), .CK(clk), .Q(
        matrix_mul_2D_1__2__1_), .QN(n2020) );
  DFF_X1 matrix_mul_2D_reg_1__2__2_ ( .D(n10944), .CK(clk), .Q(
        matrix_mul_2D_1__2__2_), .QN(n2019) );
  DFF_X1 matrix_mul_2D_reg_1__2__3_ ( .D(n10940), .CK(clk), .Q(
        matrix_mul_2D_1__2__3_), .QN(n2018) );
  DFF_X1 matrix_mul_2D_reg_1__2__4_ ( .D(n10936), .CK(clk), .Q(
        matrix_mul_2D_1__2__4_), .QN(n2017) );
  DFF_X1 matrix_mul_2D_reg_1__2__5_ ( .D(n10932), .CK(clk), .Q(
        matrix_mul_2D_1__2__5_), .QN(n2016) );
  DFF_X1 matrix_mul_2D_reg_1__2__6_ ( .D(n10928), .CK(clk), .Q(
        matrix_mul_2D_1__2__6_), .QN(n2015) );
  DFF_X1 matrix_mul_2D_reg_1__2__7_ ( .D(n10924), .CK(clk), .Q(
        matrix_mul_2D_1__2__7_), .QN(n2014) );
  DFF_X1 matrix_mul_2D_reg_1__2__8_ ( .D(n10920), .CK(clk), .Q(
        matrix_mul_2D_1__2__8_), .QN(n2013) );
  DFF_X1 matrix_mul_2D_reg_1__2__9_ ( .D(n10916), .CK(clk), .Q(
        matrix_mul_2D_1__2__9_), .QN(n2012) );
  DFF_X1 matrix_mul_2D_reg_1__2__10_ ( .D(n10912), .CK(clk), .Q(
        matrix_mul_2D_1__2__10_), .QN(n2011) );
  DFF_X1 matrix_mul_2D_reg_1__2__11_ ( .D(n10908), .CK(clk), .Q(
        matrix_mul_2D_1__2__11_), .QN(n2010) );
  DFF_X1 matrix_mul_2D_reg_1__2__12_ ( .D(n10904), .CK(clk), .Q(
        matrix_mul_2D_1__2__12_), .QN(n2009) );
  DFF_X1 matrix_mul_2D_reg_1__2__13_ ( .D(n10900), .CK(clk), .Q(
        matrix_mul_2D_1__2__13_), .QN(n2008) );
  DFF_X1 matrix_mul_2D_reg_1__2__14_ ( .D(n10896), .CK(clk), .Q(
        matrix_mul_2D_1__2__14_), .QN(n2007) );
  DFF_X1 matrix_mul_2D_reg_1__2__15_ ( .D(n10893), .CK(clk), .Q(
        matrix_mul_2D_1__2__15_), .QN(n2006) );
  DFF_X1 matrix_mul_2D_reg_1__2__16_ ( .D(n10890), .CK(clk), .Q(
        matrix_mul_2D_1__2__16_), .QN(n2005) );
  DFF_X1 matrix_mul_2D_reg_1__2__17_ ( .D(n10887), .CK(clk), .Q(
        matrix_mul_2D_1__2__17_), .QN(n2004) );
  DFF_X1 matrix_mul_2D_reg_1__2__18_ ( .D(n10884), .CK(clk), .Q(
        matrix_mul_2D_1__2__18_), .QN(n2003) );
  DFF_X1 matrix_mul_2D_reg_1__2__19_ ( .D(n10881), .CK(clk), .Q(
        matrix_mul_2D_1__2__19_), .QN(n2002) );
  DFF_X1 matrix_mul_2D_reg_1__2__20_ ( .D(n10878), .CK(clk), .Q(
        matrix_mul_2D_1__2__20_), .QN(n2001) );
  DFF_X1 matrix_mul_2D_reg_1__3__0_ ( .D(n10873), .CK(clk), .Q(
        matrix_mul_2D_1__3__0_), .QN(n2042) );
  DFF_X1 matrix_mul_2D_reg_1__3__1_ ( .D(n10869), .CK(clk), .Q(
        matrix_mul_2D_1__3__1_), .QN(n2041) );
  DFF_X1 matrix_mul_2D_reg_1__3__2_ ( .D(n10865), .CK(clk), .Q(
        matrix_mul_2D_1__3__2_), .QN(n2040) );
  DFF_X1 matrix_mul_2D_reg_1__3__3_ ( .D(n10861), .CK(clk), .Q(
        matrix_mul_2D_1__3__3_), .QN(n2039) );
  DFF_X1 matrix_mul_2D_reg_1__3__4_ ( .D(n10857), .CK(clk), .Q(
        matrix_mul_2D_1__3__4_), .QN(n2038) );
  DFF_X1 matrix_mul_2D_reg_1__3__5_ ( .D(n10853), .CK(clk), .Q(
        matrix_mul_2D_1__3__5_), .QN(n2037) );
  DFF_X1 matrix_mul_2D_reg_1__3__6_ ( .D(n10849), .CK(clk), .Q(
        matrix_mul_2D_1__3__6_), .QN(n2036) );
  DFF_X1 matrix_mul_2D_reg_1__3__7_ ( .D(n10845), .CK(clk), .Q(
        matrix_mul_2D_1__3__7_), .QN(n2035) );
  DFF_X1 matrix_mul_2D_reg_1__3__8_ ( .D(n10841), .CK(clk), .Q(
        matrix_mul_2D_1__3__8_), .QN(n2034) );
  DFF_X1 matrix_mul_2D_reg_1__3__9_ ( .D(n10837), .CK(clk), .Q(
        matrix_mul_2D_1__3__9_), .QN(n2033) );
  DFF_X1 matrix_mul_2D_reg_1__3__10_ ( .D(n10833), .CK(clk), .Q(
        matrix_mul_2D_1__3__10_), .QN(n2032) );
  DFF_X1 matrix_mul_2D_reg_1__3__11_ ( .D(n10829), .CK(clk), .Q(
        matrix_mul_2D_1__3__11_), .QN(n2031) );
  DFF_X1 matrix_mul_2D_reg_1__3__12_ ( .D(n10825), .CK(clk), .Q(
        matrix_mul_2D_1__3__12_), .QN(n2030) );
  DFF_X1 matrix_mul_2D_reg_1__3__13_ ( .D(n10821), .CK(clk), .Q(
        matrix_mul_2D_1__3__13_), .QN(n2029) );
  DFF_X1 matrix_mul_2D_reg_1__3__14_ ( .D(n10817), .CK(clk), .Q(
        matrix_mul_2D_1__3__14_), .QN(n2028) );
  DFF_X1 matrix_mul_2D_reg_1__3__15_ ( .D(n10814), .CK(clk), .Q(
        matrix_mul_2D_1__3__15_), .QN(n2027) );
  DFF_X1 matrix_mul_2D_reg_1__3__16_ ( .D(n10811), .CK(clk), .Q(
        matrix_mul_2D_1__3__16_), .QN(n2026) );
  DFF_X1 matrix_mul_2D_reg_1__3__17_ ( .D(n10808), .CK(clk), .Q(
        matrix_mul_2D_1__3__17_), .QN(n2025) );
  DFF_X1 matrix_mul_2D_reg_1__3__18_ ( .D(n10805), .CK(clk), .Q(
        matrix_mul_2D_1__3__18_), .QN(n2024) );
  DFF_X1 matrix_mul_2D_reg_1__3__19_ ( .D(n10802), .CK(clk), .Q(
        matrix_mul_2D_1__3__19_), .QN(n2023) );
  DFF_X1 matrix_mul_2D_reg_1__3__20_ ( .D(n10799), .CK(clk), .Q(
        matrix_mul_2D_1__3__20_), .QN(n2022) );
  DFF_X1 matrix_mul_2D_reg_1__4__0_ ( .D(n10794), .CK(clk), .Q(
        matrix_mul_2D_1__4__0_), .QN(n2063) );
  DFF_X1 matrix_mul_2D_reg_1__4__1_ ( .D(n10790), .CK(clk), .Q(
        matrix_mul_2D_1__4__1_), .QN(n2062) );
  DFF_X1 matrix_mul_2D_reg_1__4__2_ ( .D(n10786), .CK(clk), .Q(
        matrix_mul_2D_1__4__2_), .QN(n2061) );
  DFF_X1 matrix_mul_2D_reg_1__4__3_ ( .D(n10782), .CK(clk), .Q(
        matrix_mul_2D_1__4__3_), .QN(n2060) );
  DFF_X1 matrix_mul_2D_reg_1__4__4_ ( .D(n10778), .CK(clk), .Q(
        matrix_mul_2D_1__4__4_), .QN(n2059) );
  DFF_X1 matrix_mul_2D_reg_1__4__5_ ( .D(n10774), .CK(clk), .Q(
        matrix_mul_2D_1__4__5_), .QN(n2058) );
  DFF_X1 matrix_mul_2D_reg_1__4__6_ ( .D(n10770), .CK(clk), .Q(
        matrix_mul_2D_1__4__6_), .QN(n2057) );
  DFF_X1 matrix_mul_2D_reg_1__4__7_ ( .D(n10766), .CK(clk), .Q(
        matrix_mul_2D_1__4__7_), .QN(n2056) );
  DFF_X1 matrix_mul_2D_reg_1__4__8_ ( .D(n10762), .CK(clk), .Q(
        matrix_mul_2D_1__4__8_), .QN(n2055) );
  DFF_X1 matrix_mul_2D_reg_1__4__9_ ( .D(n10758), .CK(clk), .Q(
        matrix_mul_2D_1__4__9_), .QN(n2054) );
  DFF_X1 matrix_mul_2D_reg_1__4__10_ ( .D(n10754), .CK(clk), .Q(
        matrix_mul_2D_1__4__10_), .QN(n2053) );
  DFF_X1 matrix_mul_2D_reg_1__4__11_ ( .D(n10750), .CK(clk), .Q(
        matrix_mul_2D_1__4__11_), .QN(n2052) );
  DFF_X1 matrix_mul_2D_reg_1__4__12_ ( .D(n10746), .CK(clk), .Q(
        matrix_mul_2D_1__4__12_), .QN(n2051) );
  DFF_X1 matrix_mul_2D_reg_1__4__13_ ( .D(n10742), .CK(clk), .Q(
        matrix_mul_2D_1__4__13_), .QN(n2050) );
  DFF_X1 matrix_mul_2D_reg_1__4__14_ ( .D(n10738), .CK(clk), .Q(
        matrix_mul_2D_1__4__14_), .QN(n2049) );
  DFF_X1 matrix_mul_2D_reg_1__4__15_ ( .D(n10735), .CK(clk), .Q(
        matrix_mul_2D_1__4__15_), .QN(n2048) );
  DFF_X1 matrix_mul_2D_reg_1__4__16_ ( .D(n10732), .CK(clk), .Q(
        matrix_mul_2D_1__4__16_), .QN(n2047) );
  DFF_X1 matrix_mul_2D_reg_1__4__17_ ( .D(n10729), .CK(clk), .Q(
        matrix_mul_2D_1__4__17_), .QN(n2046) );
  DFF_X1 matrix_mul_2D_reg_1__4__18_ ( .D(n10726), .CK(clk), .Q(
        matrix_mul_2D_1__4__18_), .QN(n2045) );
  DFF_X1 matrix_mul_2D_reg_1__4__19_ ( .D(n10723), .CK(clk), .Q(
        matrix_mul_2D_1__4__19_), .QN(n2044) );
  DFF_X1 matrix_mul_2D_reg_1__4__20_ ( .D(n10720), .CK(clk), .Q(
        matrix_mul_2D_1__4__20_), .QN(n2043) );
  DFF_X1 matrix_mul_2D_reg_1__5__0_ ( .D(n10715), .CK(clk), .Q(
        matrix_mul_2D_1__5__0_), .QN(n2084) );
  DFF_X1 matrix_mul_2D_reg_1__5__1_ ( .D(n10711), .CK(clk), .Q(
        matrix_mul_2D_1__5__1_), .QN(n2083) );
  DFF_X1 matrix_mul_2D_reg_1__5__2_ ( .D(n10707), .CK(clk), .Q(
        matrix_mul_2D_1__5__2_), .QN(n2082) );
  DFF_X1 matrix_mul_2D_reg_1__5__3_ ( .D(n10703), .CK(clk), .Q(
        matrix_mul_2D_1__5__3_), .QN(n2081) );
  DFF_X1 matrix_mul_2D_reg_1__5__4_ ( .D(n10699), .CK(clk), .Q(
        matrix_mul_2D_1__5__4_), .QN(n2080) );
  DFF_X1 matrix_mul_2D_reg_1__5__5_ ( .D(n10695), .CK(clk), .Q(
        matrix_mul_2D_1__5__5_), .QN(n2079) );
  DFF_X1 matrix_mul_2D_reg_1__5__6_ ( .D(n10691), .CK(clk), .Q(
        matrix_mul_2D_1__5__6_), .QN(n2078) );
  DFF_X1 matrix_mul_2D_reg_1__5__7_ ( .D(n10687), .CK(clk), .Q(
        matrix_mul_2D_1__5__7_), .QN(n2077) );
  DFF_X1 matrix_mul_2D_reg_1__5__8_ ( .D(n10683), .CK(clk), .Q(
        matrix_mul_2D_1__5__8_), .QN(n2076) );
  DFF_X1 matrix_mul_2D_reg_1__5__9_ ( .D(n10679), .CK(clk), .Q(
        matrix_mul_2D_1__5__9_), .QN(n2075) );
  DFF_X1 matrix_mul_2D_reg_1__5__10_ ( .D(n10675), .CK(clk), .Q(
        matrix_mul_2D_1__5__10_), .QN(n2074) );
  DFF_X1 matrix_mul_2D_reg_1__5__11_ ( .D(n10671), .CK(clk), .Q(
        matrix_mul_2D_1__5__11_), .QN(n2073) );
  DFF_X1 matrix_mul_2D_reg_1__5__12_ ( .D(n10667), .CK(clk), .Q(
        matrix_mul_2D_1__5__12_), .QN(n2072) );
  DFF_X1 matrix_mul_2D_reg_1__5__13_ ( .D(n10663), .CK(clk), .Q(
        matrix_mul_2D_1__5__13_), .QN(n2071) );
  DFF_X1 matrix_mul_2D_reg_1__5__14_ ( .D(n10659), .CK(clk), .Q(
        matrix_mul_2D_1__5__14_), .QN(n2070) );
  DFF_X1 matrix_mul_2D_reg_1__5__15_ ( .D(n10656), .CK(clk), .Q(
        matrix_mul_2D_1__5__15_), .QN(n2069) );
  DFF_X1 matrix_mul_2D_reg_1__5__16_ ( .D(n10653), .CK(clk), .Q(
        matrix_mul_2D_1__5__16_), .QN(n2068) );
  DFF_X1 matrix_mul_2D_reg_1__5__17_ ( .D(n10650), .CK(clk), .Q(
        matrix_mul_2D_1__5__17_), .QN(n2067) );
  DFF_X1 matrix_mul_2D_reg_1__5__18_ ( .D(n10647), .CK(clk), .Q(
        matrix_mul_2D_1__5__18_), .QN(n2066) );
  DFF_X1 matrix_mul_2D_reg_1__5__19_ ( .D(n10644), .CK(clk), .Q(
        matrix_mul_2D_1__5__19_), .QN(n2065) );
  DFF_X1 matrix_mul_2D_reg_1__5__20_ ( .D(n10641), .CK(clk), .Q(
        matrix_mul_2D_1__5__20_), .QN(n2064) );
  DFF_X1 matrix_mul_2D_reg_1__6__0_ ( .D(n10637), .CK(clk), .Q(
        matrix_mul_2D_1__6__0_), .QN(n2099) );
  DFF_X1 matrix_mul_2D_reg_1__6__1_ ( .D(n10632), .CK(clk), .Q(
        matrix_mul_2D_1__6__1_), .QN(n2098) );
  DFF_X1 matrix_mul_2D_reg_1__6__2_ ( .D(n10627), .CK(clk), .Q(
        matrix_mul_2D_1__6__2_), .QN(n2097) );
  DFF_X1 matrix_mul_2D_reg_1__6__3_ ( .D(n10622), .CK(clk), .Q(
        matrix_mul_2D_1__6__3_), .QN(n2096) );
  DFF_X1 matrix_mul_2D_reg_1__6__4_ ( .D(n10617), .CK(clk), .Q(
        matrix_mul_2D_1__6__4_), .QN(n2095) );
  DFF_X1 matrix_mul_2D_reg_1__6__5_ ( .D(n10612), .CK(clk), .Q(
        matrix_mul_2D_1__6__5_), .QN(n2094) );
  DFF_X1 matrix_mul_2D_reg_1__6__6_ ( .D(n10607), .CK(clk), .Q(
        matrix_mul_2D_1__6__6_), .QN(n2093) );
  DFF_X1 matrix_mul_2D_reg_1__6__7_ ( .D(n10602), .CK(clk), .Q(
        matrix_mul_2D_1__6__7_), .QN(n2092) );
  DFF_X1 matrix_mul_2D_reg_1__6__8_ ( .D(n10597), .CK(clk), .Q(
        matrix_mul_2D_1__6__8_), .QN(n2091) );
  DFF_X1 matrix_mul_2D_reg_1__6__9_ ( .D(n10592), .CK(clk), .Q(
        matrix_mul_2D_1__6__9_), .QN(n2090) );
  DFF_X1 matrix_mul_2D_reg_1__6__10_ ( .D(n10587), .CK(clk), .Q(
        matrix_mul_2D_1__6__10_), .QN(n2089) );
  DFF_X1 matrix_mul_2D_reg_1__6__11_ ( .D(n10582), .CK(clk), .Q(
        matrix_mul_2D_1__6__11_), .QN(n2088) );
  DFF_X1 matrix_mul_2D_reg_1__6__12_ ( .D(n10577), .CK(clk), .Q(
        matrix_mul_2D_1__6__12_), .QN(n2087) );
  DFF_X1 matrix_mul_2D_reg_1__6__13_ ( .D(n10572), .CK(clk), .Q(
        matrix_mul_2D_1__6__13_), .QN(n2086) );
  DFF_X1 matrix_mul_2D_reg_1__6__14_ ( .D(n10567), .CK(clk), .Q(
        matrix_mul_2D_1__6__14_), .QN(n2085) );
  DFF_X1 matrix_mul_2D_reg_1__6__15_ ( .D(n10566), .CK(clk), .Q(
        matrix_mul_2D_1__6__15_), .QN(n17868) );
  DFF_X1 matrix_mul_2D_reg_1__6__16_ ( .D(n10565), .CK(clk), .Q(
        matrix_mul_2D_1__6__16_), .QN(n17866) );
  DFF_X1 matrix_mul_2D_reg_1__6__17_ ( .D(n10564), .CK(clk), .Q(
        matrix_mul_2D_1__6__17_), .QN(n17864) );
  DFF_X1 matrix_mul_2D_reg_1__6__18_ ( .D(n10563), .CK(clk), .Q(
        matrix_mul_2D_1__6__18_), .QN(n17862) );
  DFF_X1 matrix_mul_2D_reg_1__6__19_ ( .D(n10562), .CK(clk), .Q(
        matrix_mul_2D_1__6__19_), .QN(n17860) );
  DFF_X1 matrix_mul_2D_reg_1__6__20_ ( .D(n10561), .CK(clk), .Q(
        matrix_mul_2D_1__6__20_), .QN(n17858) );
  DFF_X1 matrix_mul_2D_reg_1__7__0_ ( .D(n10557), .CK(clk), .Q(
        matrix_mul_2D_1__7__0_), .QN(n2114) );
  DFF_X1 matrix_mul_2D_reg_1__7__1_ ( .D(n10552), .CK(clk), .Q(
        matrix_mul_2D_1__7__1_), .QN(n2113) );
  DFF_X1 matrix_mul_2D_reg_1__7__2_ ( .D(n10547), .CK(clk), .Q(
        matrix_mul_2D_1__7__2_), .QN(n2112) );
  DFF_X1 matrix_mul_2D_reg_1__7__3_ ( .D(n10542), .CK(clk), .Q(
        matrix_mul_2D_1__7__3_), .QN(n2111) );
  DFF_X1 matrix_mul_2D_reg_1__7__4_ ( .D(n10537), .CK(clk), .Q(
        matrix_mul_2D_1__7__4_), .QN(n2110) );
  DFF_X1 matrix_mul_2D_reg_1__7__5_ ( .D(n10532), .CK(clk), .Q(
        matrix_mul_2D_1__7__5_), .QN(n2109) );
  DFF_X1 matrix_mul_2D_reg_1__7__6_ ( .D(n10527), .CK(clk), .Q(
        matrix_mul_2D_1__7__6_), .QN(n2108) );
  DFF_X1 matrix_mul_2D_reg_1__7__7_ ( .D(n10522), .CK(clk), .Q(
        matrix_mul_2D_1__7__7_), .QN(n2107) );
  DFF_X1 matrix_mul_2D_reg_1__7__8_ ( .D(n10517), .CK(clk), .Q(
        matrix_mul_2D_1__7__8_), .QN(n2106) );
  DFF_X1 matrix_mul_2D_reg_1__7__9_ ( .D(n10512), .CK(clk), .Q(
        matrix_mul_2D_1__7__9_), .QN(n2105) );
  DFF_X1 matrix_mul_2D_reg_1__7__10_ ( .D(n10507), .CK(clk), .Q(
        matrix_mul_2D_1__7__10_), .QN(n2104) );
  DFF_X1 matrix_mul_2D_reg_1__7__11_ ( .D(n10502), .CK(clk), .Q(
        matrix_mul_2D_1__7__11_), .QN(n2103) );
  DFF_X1 matrix_mul_2D_reg_1__7__12_ ( .D(n10497), .CK(clk), .Q(
        matrix_mul_2D_1__7__12_), .QN(n2102) );
  DFF_X1 matrix_mul_2D_reg_1__7__13_ ( .D(n10492), .CK(clk), .Q(
        matrix_mul_2D_1__7__13_), .QN(n2101) );
  DFF_X1 matrix_mul_2D_reg_1__7__14_ ( .D(n10487), .CK(clk), .Q(
        matrix_mul_2D_1__7__14_), .QN(n2100) );
  DFF_X1 matrix_mul_2D_reg_1__7__15_ ( .D(n10486), .CK(clk), .Q(
        matrix_mul_2D_1__7__15_), .QN(n17856) );
  DFF_X1 matrix_mul_2D_reg_1__7__16_ ( .D(n10485), .CK(clk), .Q(
        matrix_mul_2D_1__7__16_), .QN(n17854) );
  DFF_X1 matrix_mul_2D_reg_1__7__17_ ( .D(n10484), .CK(clk), .Q(
        matrix_mul_2D_1__7__17_), .QN(n17852) );
  DFF_X1 matrix_mul_2D_reg_1__7__18_ ( .D(n10483), .CK(clk), .Q(
        matrix_mul_2D_1__7__18_), .QN(n17850) );
  DFF_X1 matrix_mul_2D_reg_1__7__19_ ( .D(n10482), .CK(clk), .Q(
        matrix_mul_2D_1__7__19_), .QN(n17848) );
  DFF_X1 matrix_mul_2D_reg_1__7__20_ ( .D(n10481), .CK(clk), .Q(
        matrix_mul_2D_1__7__20_), .QN(n17846) );
  DFF_X1 matrix_mul_2D_reg_2__0__0_ ( .D(n10477), .CK(clk), .Q(
        matrix_mul_2D_2__0__0_), .QN(n2129) );
  DFF_X1 matrix_mul_2D_reg_2__0__1_ ( .D(n10472), .CK(clk), .Q(
        matrix_mul_2D_2__0__1_), .QN(n2128) );
  DFF_X1 matrix_mul_2D_reg_2__0__2_ ( .D(n10467), .CK(clk), .Q(
        matrix_mul_2D_2__0__2_), .QN(n2127) );
  DFF_X1 matrix_mul_2D_reg_2__0__3_ ( .D(n10462), .CK(clk), .Q(
        matrix_mul_2D_2__0__3_), .QN(n2126) );
  DFF_X1 matrix_mul_2D_reg_2__0__4_ ( .D(n10457), .CK(clk), .Q(
        matrix_mul_2D_2__0__4_), .QN(n2125) );
  DFF_X1 matrix_mul_2D_reg_2__0__5_ ( .D(n10452), .CK(clk), .Q(
        matrix_mul_2D_2__0__5_), .QN(n2124) );
  DFF_X1 matrix_mul_2D_reg_2__0__6_ ( .D(n10447), .CK(clk), .Q(
        matrix_mul_2D_2__0__6_), .QN(n2123) );
  DFF_X1 matrix_mul_2D_reg_2__0__7_ ( .D(n10442), .CK(clk), .Q(
        matrix_mul_2D_2__0__7_), .QN(n2122) );
  DFF_X1 matrix_mul_2D_reg_2__0__8_ ( .D(n10437), .CK(clk), .Q(
        matrix_mul_2D_2__0__8_), .QN(n2121) );
  DFF_X1 matrix_mul_2D_reg_2__0__9_ ( .D(n10432), .CK(clk), .Q(
        matrix_mul_2D_2__0__9_), .QN(n2120) );
  DFF_X1 matrix_mul_2D_reg_2__0__10_ ( .D(n10427), .CK(clk), .Q(
        matrix_mul_2D_2__0__10_), .QN(n2119) );
  DFF_X1 matrix_mul_2D_reg_2__0__11_ ( .D(n10422), .CK(clk), .Q(
        matrix_mul_2D_2__0__11_), .QN(n2118) );
  DFF_X1 matrix_mul_2D_reg_2__0__12_ ( .D(n10417), .CK(clk), .Q(
        matrix_mul_2D_2__0__12_), .QN(n2117) );
  DFF_X1 matrix_mul_2D_reg_2__0__13_ ( .D(n10412), .CK(clk), .Q(
        matrix_mul_2D_2__0__13_), .QN(n2116) );
  DFF_X1 matrix_mul_2D_reg_2__0__14_ ( .D(n10407), .CK(clk), .Q(
        matrix_mul_2D_2__0__14_), .QN(n2115) );
  DFF_X1 matrix_mul_2D_reg_2__0__15_ ( .D(n10406), .CK(clk), .Q(
        matrix_mul_2D_2__0__15_), .QN(n17844) );
  DFF_X1 matrix_mul_2D_reg_2__0__16_ ( .D(n10405), .CK(clk), .Q(
        matrix_mul_2D_2__0__16_), .QN(n17842) );
  DFF_X1 matrix_mul_2D_reg_2__0__17_ ( .D(n10404), .CK(clk), .Q(
        matrix_mul_2D_2__0__17_), .QN(n17840) );
  DFF_X1 matrix_mul_2D_reg_2__0__18_ ( .D(n10403), .CK(clk), .Q(
        matrix_mul_2D_2__0__18_), .QN(n17838) );
  DFF_X1 matrix_mul_2D_reg_2__0__19_ ( .D(n10402), .CK(clk), .Q(
        matrix_mul_2D_2__0__19_), .QN(n17836) );
  DFF_X1 matrix_mul_2D_reg_2__0__20_ ( .D(n10401), .CK(clk), .Q(
        matrix_mul_2D_2__0__20_), .QN(n17834) );
  DFF_X1 matrix_mul_2D_reg_2__1__0_ ( .D(n10397), .CK(clk), .Q(
        matrix_mul_2D_2__1__0_), .QN(n2144) );
  DFF_X1 matrix_mul_2D_reg_2__1__1_ ( .D(n10392), .CK(clk), .Q(
        matrix_mul_2D_2__1__1_), .QN(n2143) );
  DFF_X1 matrix_mul_2D_reg_2__1__2_ ( .D(n10387), .CK(clk), .Q(
        matrix_mul_2D_2__1__2_), .QN(n2142) );
  DFF_X1 matrix_mul_2D_reg_2__1__3_ ( .D(n10382), .CK(clk), .Q(
        matrix_mul_2D_2__1__3_), .QN(n2141) );
  DFF_X1 matrix_mul_2D_reg_2__1__4_ ( .D(n10377), .CK(clk), .Q(
        matrix_mul_2D_2__1__4_), .QN(n2140) );
  DFF_X1 matrix_mul_2D_reg_2__1__5_ ( .D(n10372), .CK(clk), .Q(
        matrix_mul_2D_2__1__5_), .QN(n2139) );
  DFF_X1 matrix_mul_2D_reg_2__1__6_ ( .D(n10367), .CK(clk), .Q(
        matrix_mul_2D_2__1__6_), .QN(n2138) );
  DFF_X1 matrix_mul_2D_reg_2__1__7_ ( .D(n10362), .CK(clk), .Q(
        matrix_mul_2D_2__1__7_), .QN(n2137) );
  DFF_X1 matrix_mul_2D_reg_2__1__8_ ( .D(n10357), .CK(clk), .Q(
        matrix_mul_2D_2__1__8_), .QN(n2136) );
  DFF_X1 matrix_mul_2D_reg_2__1__9_ ( .D(n10352), .CK(clk), .Q(
        matrix_mul_2D_2__1__9_), .QN(n2135) );
  DFF_X1 matrix_mul_2D_reg_2__1__10_ ( .D(n10347), .CK(clk), .Q(
        matrix_mul_2D_2__1__10_), .QN(n2134) );
  DFF_X1 matrix_mul_2D_reg_2__1__11_ ( .D(n10342), .CK(clk), .Q(
        matrix_mul_2D_2__1__11_), .QN(n2133) );
  DFF_X1 matrix_mul_2D_reg_2__1__12_ ( .D(n10337), .CK(clk), .Q(
        matrix_mul_2D_2__1__12_), .QN(n2132) );
  DFF_X1 matrix_mul_2D_reg_2__1__13_ ( .D(n10332), .CK(clk), .Q(
        matrix_mul_2D_2__1__13_), .QN(n2131) );
  DFF_X1 matrix_mul_2D_reg_2__1__14_ ( .D(n10327), .CK(clk), .Q(
        matrix_mul_2D_2__1__14_), .QN(n2130) );
  DFF_X1 matrix_mul_2D_reg_2__1__15_ ( .D(n10326), .CK(clk), .Q(
        matrix_mul_2D_2__1__15_), .QN(n17832) );
  DFF_X1 matrix_mul_2D_reg_2__1__16_ ( .D(n10325), .CK(clk), .Q(
        matrix_mul_2D_2__1__16_), .QN(n17830) );
  DFF_X1 matrix_mul_2D_reg_2__1__17_ ( .D(n10324), .CK(clk), .Q(
        matrix_mul_2D_2__1__17_), .QN(n17828) );
  DFF_X1 matrix_mul_2D_reg_2__1__18_ ( .D(n10323), .CK(clk), .Q(
        matrix_mul_2D_2__1__18_), .QN(n17826) );
  DFF_X1 matrix_mul_2D_reg_2__1__19_ ( .D(n10322), .CK(clk), .Q(
        matrix_mul_2D_2__1__19_), .QN(n17824) );
  DFF_X1 matrix_mul_2D_reg_2__1__20_ ( .D(n10321), .CK(clk), .Q(
        matrix_mul_2D_2__1__20_), .QN(n17822) );
  DFF_X1 matrix_mul_2D_reg_2__2__0_ ( .D(n10317), .CK(clk), .Q(
        matrix_mul_2D_2__2__0_), .QN(n2159) );
  DFF_X1 matrix_mul_2D_reg_2__2__1_ ( .D(n10312), .CK(clk), .Q(
        matrix_mul_2D_2__2__1_), .QN(n2158) );
  DFF_X1 matrix_mul_2D_reg_2__2__2_ ( .D(n10307), .CK(clk), .Q(
        matrix_mul_2D_2__2__2_), .QN(n2157) );
  DFF_X1 matrix_mul_2D_reg_2__2__3_ ( .D(n10302), .CK(clk), .Q(
        matrix_mul_2D_2__2__3_), .QN(n2156) );
  DFF_X1 matrix_mul_2D_reg_2__2__4_ ( .D(n10297), .CK(clk), .Q(
        matrix_mul_2D_2__2__4_), .QN(n2155) );
  DFF_X1 matrix_mul_2D_reg_2__2__5_ ( .D(n10292), .CK(clk), .Q(
        matrix_mul_2D_2__2__5_), .QN(n2154) );
  DFF_X1 matrix_mul_2D_reg_2__2__6_ ( .D(n10287), .CK(clk), .Q(
        matrix_mul_2D_2__2__6_), .QN(n2153) );
  DFF_X1 matrix_mul_2D_reg_2__2__7_ ( .D(n10282), .CK(clk), .Q(
        matrix_mul_2D_2__2__7_), .QN(n2152) );
  DFF_X1 matrix_mul_2D_reg_2__2__8_ ( .D(n10277), .CK(clk), .Q(
        matrix_mul_2D_2__2__8_), .QN(n2151) );
  DFF_X1 matrix_mul_2D_reg_2__2__9_ ( .D(n10272), .CK(clk), .Q(
        matrix_mul_2D_2__2__9_), .QN(n2150) );
  DFF_X1 matrix_mul_2D_reg_2__2__10_ ( .D(n10267), .CK(clk), .Q(
        matrix_mul_2D_2__2__10_), .QN(n2149) );
  DFF_X1 matrix_mul_2D_reg_2__2__11_ ( .D(n10262), .CK(clk), .Q(
        matrix_mul_2D_2__2__11_), .QN(n2148) );
  DFF_X1 matrix_mul_2D_reg_2__2__12_ ( .D(n10257), .CK(clk), .Q(
        matrix_mul_2D_2__2__12_), .QN(n2147) );
  DFF_X1 matrix_mul_2D_reg_2__2__13_ ( .D(n10252), .CK(clk), .Q(
        matrix_mul_2D_2__2__13_), .QN(n2146) );
  DFF_X1 matrix_mul_2D_reg_2__2__14_ ( .D(n10247), .CK(clk), .Q(
        matrix_mul_2D_2__2__14_), .QN(n2145) );
  DFF_X1 matrix_mul_2D_reg_2__2__15_ ( .D(n10246), .CK(clk), .Q(
        matrix_mul_2D_2__2__15_), .QN(n17820) );
  DFF_X1 matrix_mul_2D_reg_2__2__16_ ( .D(n10245), .CK(clk), .Q(
        matrix_mul_2D_2__2__16_), .QN(n17818) );
  DFF_X1 matrix_mul_2D_reg_2__2__17_ ( .D(n10244), .CK(clk), .Q(
        matrix_mul_2D_2__2__17_), .QN(n17816) );
  DFF_X1 matrix_mul_2D_reg_2__2__18_ ( .D(n10243), .CK(clk), .Q(
        matrix_mul_2D_2__2__18_), .QN(n17814) );
  DFF_X1 matrix_mul_2D_reg_2__2__19_ ( .D(n10242), .CK(clk), .Q(
        matrix_mul_2D_2__2__19_), .QN(n17812) );
  DFF_X1 matrix_mul_2D_reg_2__2__20_ ( .D(n10241), .CK(clk), .Q(
        matrix_mul_2D_2__2__20_), .QN(n17810) );
  DFF_X1 matrix_mul_2D_reg_2__3__0_ ( .D(n10237), .CK(clk), .Q(
        matrix_mul_2D_2__3__0_), .QN(n2174) );
  DFF_X1 matrix_mul_2D_reg_2__3__1_ ( .D(n10232), .CK(clk), .Q(
        matrix_mul_2D_2__3__1_), .QN(n2173) );
  DFF_X1 matrix_mul_2D_reg_2__3__2_ ( .D(n10227), .CK(clk), .Q(
        matrix_mul_2D_2__3__2_), .QN(n2172) );
  DFF_X1 matrix_mul_2D_reg_2__3__3_ ( .D(n10222), .CK(clk), .Q(
        matrix_mul_2D_2__3__3_), .QN(n2171) );
  DFF_X1 matrix_mul_2D_reg_2__3__4_ ( .D(n10217), .CK(clk), .Q(
        matrix_mul_2D_2__3__4_), .QN(n2170) );
  DFF_X1 matrix_mul_2D_reg_2__3__5_ ( .D(n10212), .CK(clk), .Q(
        matrix_mul_2D_2__3__5_), .QN(n2169) );
  DFF_X1 matrix_mul_2D_reg_2__3__6_ ( .D(n10207), .CK(clk), .Q(
        matrix_mul_2D_2__3__6_), .QN(n2168) );
  DFF_X1 matrix_mul_2D_reg_2__3__7_ ( .D(n10202), .CK(clk), .Q(
        matrix_mul_2D_2__3__7_), .QN(n2167) );
  DFF_X1 matrix_mul_2D_reg_2__3__8_ ( .D(n10197), .CK(clk), .Q(
        matrix_mul_2D_2__3__8_), .QN(n2166) );
  DFF_X1 matrix_mul_2D_reg_2__3__9_ ( .D(n10192), .CK(clk), .Q(
        matrix_mul_2D_2__3__9_), .QN(n2165) );
  DFF_X1 matrix_mul_2D_reg_2__3__10_ ( .D(n10187), .CK(clk), .Q(
        matrix_mul_2D_2__3__10_), .QN(n2164) );
  DFF_X1 matrix_mul_2D_reg_2__3__11_ ( .D(n10182), .CK(clk), .Q(
        matrix_mul_2D_2__3__11_), .QN(n2163) );
  DFF_X1 matrix_mul_2D_reg_2__3__12_ ( .D(n10177), .CK(clk), .Q(
        matrix_mul_2D_2__3__12_), .QN(n2162) );
  DFF_X1 matrix_mul_2D_reg_2__3__13_ ( .D(n10172), .CK(clk), .Q(
        matrix_mul_2D_2__3__13_), .QN(n2161) );
  DFF_X1 matrix_mul_2D_reg_2__3__14_ ( .D(n10167), .CK(clk), .Q(
        matrix_mul_2D_2__3__14_), .QN(n2160) );
  DFF_X1 matrix_mul_2D_reg_2__3__15_ ( .D(n10166), .CK(clk), .Q(
        matrix_mul_2D_2__3__15_), .QN(n17808) );
  DFF_X1 matrix_mul_2D_reg_2__3__16_ ( .D(n10165), .CK(clk), .Q(
        matrix_mul_2D_2__3__16_), .QN(n17806) );
  DFF_X1 matrix_mul_2D_reg_2__3__17_ ( .D(n10164), .CK(clk), .Q(
        matrix_mul_2D_2__3__17_), .QN(n17804) );
  DFF_X1 matrix_mul_2D_reg_2__3__18_ ( .D(n10163), .CK(clk), .Q(
        matrix_mul_2D_2__3__18_), .QN(n17802) );
  DFF_X1 matrix_mul_2D_reg_2__3__19_ ( .D(n10162), .CK(clk), .Q(
        matrix_mul_2D_2__3__19_), .QN(n17800) );
  DFF_X1 matrix_mul_2D_reg_2__3__20_ ( .D(n10161), .CK(clk), .Q(
        matrix_mul_2D_2__3__20_), .QN(n17798) );
  DFF_X1 matrix_mul_2D_reg_2__4__0_ ( .D(n10157), .CK(clk), .Q(
        matrix_mul_2D_2__4__0_), .QN(n2189) );
  DFF_X1 matrix_mul_2D_reg_2__4__1_ ( .D(n10152), .CK(clk), .Q(
        matrix_mul_2D_2__4__1_), .QN(n2188) );
  DFF_X1 matrix_mul_2D_reg_2__4__2_ ( .D(n10147), .CK(clk), .Q(
        matrix_mul_2D_2__4__2_), .QN(n2187) );
  DFF_X1 matrix_mul_2D_reg_2__4__3_ ( .D(n10142), .CK(clk), .Q(
        matrix_mul_2D_2__4__3_), .QN(n2186) );
  DFF_X1 matrix_mul_2D_reg_2__4__4_ ( .D(n10137), .CK(clk), .Q(
        matrix_mul_2D_2__4__4_), .QN(n2185) );
  DFF_X1 matrix_mul_2D_reg_2__4__5_ ( .D(n10132), .CK(clk), .Q(
        matrix_mul_2D_2__4__5_), .QN(n2184) );
  DFF_X1 matrix_mul_2D_reg_2__4__6_ ( .D(n10127), .CK(clk), .Q(
        matrix_mul_2D_2__4__6_), .QN(n2183) );
  DFF_X1 matrix_mul_2D_reg_2__4__7_ ( .D(n10122), .CK(clk), .Q(
        matrix_mul_2D_2__4__7_), .QN(n2182) );
  DFF_X1 matrix_mul_2D_reg_2__4__8_ ( .D(n10117), .CK(clk), .Q(
        matrix_mul_2D_2__4__8_), .QN(n2181) );
  DFF_X1 matrix_mul_2D_reg_2__4__9_ ( .D(n10112), .CK(clk), .Q(
        matrix_mul_2D_2__4__9_), .QN(n2180) );
  DFF_X1 matrix_mul_2D_reg_2__4__10_ ( .D(n10107), .CK(clk), .Q(
        matrix_mul_2D_2__4__10_), .QN(n2179) );
  DFF_X1 matrix_mul_2D_reg_2__4__11_ ( .D(n10102), .CK(clk), .Q(
        matrix_mul_2D_2__4__11_), .QN(n2178) );
  DFF_X1 matrix_mul_2D_reg_2__4__12_ ( .D(n10097), .CK(clk), .Q(
        matrix_mul_2D_2__4__12_), .QN(n2177) );
  DFF_X1 matrix_mul_2D_reg_2__4__13_ ( .D(n10092), .CK(clk), .Q(
        matrix_mul_2D_2__4__13_), .QN(n2176) );
  DFF_X1 matrix_mul_2D_reg_2__4__14_ ( .D(n10087), .CK(clk), .Q(
        matrix_mul_2D_2__4__14_), .QN(n2175) );
  DFF_X1 matrix_mul_2D_reg_2__4__15_ ( .D(n10086), .CK(clk), .Q(
        matrix_mul_2D_2__4__15_), .QN(n17796) );
  DFF_X1 matrix_mul_2D_reg_2__4__16_ ( .D(n10085), .CK(clk), .Q(
        matrix_mul_2D_2__4__16_), .QN(n17794) );
  DFF_X1 matrix_mul_2D_reg_2__4__17_ ( .D(n10084), .CK(clk), .Q(
        matrix_mul_2D_2__4__17_), .QN(n17792) );
  DFF_X1 matrix_mul_2D_reg_2__4__18_ ( .D(n10083), .CK(clk), .Q(
        matrix_mul_2D_2__4__18_), .QN(n17790) );
  DFF_X1 matrix_mul_2D_reg_2__4__19_ ( .D(n10082), .CK(clk), .Q(
        matrix_mul_2D_2__4__19_), .QN(n17788) );
  DFF_X1 matrix_mul_2D_reg_2__4__20_ ( .D(n10081), .CK(clk), .Q(
        matrix_mul_2D_2__4__20_), .QN(n17786) );
  DFF_X1 matrix_mul_2D_reg_2__5__0_ ( .D(n10077), .CK(clk), .Q(
        matrix_mul_2D_2__5__0_), .QN(n2204) );
  DFF_X1 matrix_mul_2D_reg_2__5__1_ ( .D(n10072), .CK(clk), .Q(
        matrix_mul_2D_2__5__1_), .QN(n2203) );
  DFF_X1 matrix_mul_2D_reg_2__5__2_ ( .D(n10067), .CK(clk), .Q(
        matrix_mul_2D_2__5__2_), .QN(n2202) );
  DFF_X1 matrix_mul_2D_reg_2__5__3_ ( .D(n10062), .CK(clk), .Q(
        matrix_mul_2D_2__5__3_), .QN(n2201) );
  DFF_X1 matrix_mul_2D_reg_2__5__4_ ( .D(n10057), .CK(clk), .Q(
        matrix_mul_2D_2__5__4_), .QN(n2200) );
  DFF_X1 matrix_mul_2D_reg_2__5__5_ ( .D(n10052), .CK(clk), .Q(
        matrix_mul_2D_2__5__5_), .QN(n2199) );
  DFF_X1 matrix_mul_2D_reg_2__5__6_ ( .D(n10047), .CK(clk), .Q(
        matrix_mul_2D_2__5__6_), .QN(n2198) );
  DFF_X1 matrix_mul_2D_reg_2__5__7_ ( .D(n10042), .CK(clk), .Q(
        matrix_mul_2D_2__5__7_), .QN(n2197) );
  DFF_X1 matrix_mul_2D_reg_2__5__8_ ( .D(n10037), .CK(clk), .Q(
        matrix_mul_2D_2__5__8_), .QN(n2196) );
  DFF_X1 matrix_mul_2D_reg_2__5__9_ ( .D(n10032), .CK(clk), .Q(
        matrix_mul_2D_2__5__9_), .QN(n2195) );
  DFF_X1 matrix_mul_2D_reg_2__5__10_ ( .D(n10027), .CK(clk), .Q(
        matrix_mul_2D_2__5__10_), .QN(n2194) );
  DFF_X1 matrix_mul_2D_reg_2__5__11_ ( .D(n10022), .CK(clk), .Q(
        matrix_mul_2D_2__5__11_), .QN(n2193) );
  DFF_X1 matrix_mul_2D_reg_2__5__12_ ( .D(n10017), .CK(clk), .Q(
        matrix_mul_2D_2__5__12_), .QN(n2192) );
  DFF_X1 matrix_mul_2D_reg_2__5__13_ ( .D(n10012), .CK(clk), .Q(
        matrix_mul_2D_2__5__13_), .QN(n2191) );
  DFF_X1 matrix_mul_2D_reg_2__5__14_ ( .D(n10007), .CK(clk), .Q(
        matrix_mul_2D_2__5__14_), .QN(n2190) );
  DFF_X1 matrix_mul_2D_reg_2__5__15_ ( .D(n10006), .CK(clk), .Q(
        matrix_mul_2D_2__5__15_), .QN(n17784) );
  DFF_X1 matrix_mul_2D_reg_2__5__16_ ( .D(n10005), .CK(clk), .Q(
        matrix_mul_2D_2__5__16_), .QN(n17782) );
  DFF_X1 matrix_mul_2D_reg_2__5__17_ ( .D(n10004), .CK(clk), .Q(
        matrix_mul_2D_2__5__17_), .QN(n17780) );
  DFF_X1 matrix_mul_2D_reg_2__5__18_ ( .D(n10003), .CK(clk), .Q(
        matrix_mul_2D_2__5__18_), .QN(n17778) );
  DFF_X1 matrix_mul_2D_reg_2__5__19_ ( .D(n10002), .CK(clk), .Q(
        matrix_mul_2D_2__5__19_), .QN(n17776) );
  DFF_X1 matrix_mul_2D_reg_2__5__20_ ( .D(n10001), .CK(clk), .Q(
        matrix_mul_2D_2__5__20_), .QN(n17774) );
  DFF_X1 matrix_mul_2D_reg_2__6__0_ ( .D(n9996), .CK(clk), .Q(
        matrix_mul_2D_2__6__0_), .QN(n2225) );
  DFF_X1 matrix_mul_2D_reg_2__6__1_ ( .D(n9992), .CK(clk), .Q(
        matrix_mul_2D_2__6__1_), .QN(n2224) );
  DFF_X1 matrix_mul_2D_reg_2__6__2_ ( .D(n9988), .CK(clk), .Q(
        matrix_mul_2D_2__6__2_), .QN(n2223) );
  DFF_X1 matrix_mul_2D_reg_2__6__3_ ( .D(n9984), .CK(clk), .Q(
        matrix_mul_2D_2__6__3_), .QN(n2222) );
  DFF_X1 matrix_mul_2D_reg_2__6__4_ ( .D(n9980), .CK(clk), .Q(
        matrix_mul_2D_2__6__4_), .QN(n2221) );
  DFF_X1 matrix_mul_2D_reg_2__6__5_ ( .D(n9976), .CK(clk), .Q(
        matrix_mul_2D_2__6__5_), .QN(n2220) );
  DFF_X1 matrix_mul_2D_reg_2__6__6_ ( .D(n9972), .CK(clk), .Q(
        matrix_mul_2D_2__6__6_), .QN(n2219) );
  DFF_X1 matrix_mul_2D_reg_2__6__7_ ( .D(n9968), .CK(clk), .Q(
        matrix_mul_2D_2__6__7_), .QN(n2218) );
  DFF_X1 matrix_mul_2D_reg_2__6__8_ ( .D(n9964), .CK(clk), .Q(
        matrix_mul_2D_2__6__8_), .QN(n2217) );
  DFF_X1 matrix_mul_2D_reg_2__6__9_ ( .D(n9960), .CK(clk), .Q(
        matrix_mul_2D_2__6__9_), .QN(n2216) );
  DFF_X1 matrix_mul_2D_reg_2__6__10_ ( .D(n9956), .CK(clk), .Q(
        matrix_mul_2D_2__6__10_), .QN(n2215) );
  DFF_X1 matrix_mul_2D_reg_2__6__11_ ( .D(n9952), .CK(clk), .Q(
        matrix_mul_2D_2__6__11_), .QN(n2214) );
  DFF_X1 matrix_mul_2D_reg_2__6__12_ ( .D(n9948), .CK(clk), .Q(
        matrix_mul_2D_2__6__12_), .QN(n2213) );
  DFF_X1 matrix_mul_2D_reg_2__6__13_ ( .D(n9944), .CK(clk), .Q(
        matrix_mul_2D_2__6__13_), .QN(n2212) );
  DFF_X1 matrix_mul_2D_reg_2__6__14_ ( .D(n9940), .CK(clk), .Q(
        matrix_mul_2D_2__6__14_), .QN(n2211) );
  DFF_X1 matrix_mul_2D_reg_2__6__15_ ( .D(n9939), .CK(clk), .Q(
        matrix_mul_2D_2__6__15_), .QN(n17772) );
  DFF_X1 matrix_mul_2D_reg_2__6__16_ ( .D(n9938), .CK(clk), .Q(
        matrix_mul_2D_2__6__16_), .QN(n17770) );
  DFF_X1 matrix_mul_2D_reg_2__6__17_ ( .D(n9937), .CK(clk), .Q(
        matrix_mul_2D_2__6__17_), .QN(n17768) );
  DFF_X1 matrix_mul_2D_reg_2__6__18_ ( .D(n9936), .CK(clk), .Q(
        matrix_mul_2D_2__6__18_), .QN(n17766) );
  DFF_X1 matrix_mul_2D_reg_2__6__19_ ( .D(n9935), .CK(clk), .Q(
        matrix_mul_2D_2__6__19_), .QN(n17764) );
  DFF_X1 matrix_mul_2D_reg_2__6__20_ ( .D(n9934), .CK(clk), .Q(
        matrix_mul_2D_2__6__20_), .QN(n17762) );
  DFF_X1 matrix_mul_2D_reg_2__7__0_ ( .D(n9929), .CK(clk), .Q(
        matrix_mul_2D_2__7__0_), .QN(n2240) );
  DFF_X1 matrix_mul_2D_reg_2__7__1_ ( .D(n9925), .CK(clk), .Q(
        matrix_mul_2D_2__7__1_), .QN(n2239) );
  DFF_X1 matrix_mul_2D_reg_2__7__2_ ( .D(n9921), .CK(clk), .Q(
        matrix_mul_2D_2__7__2_), .QN(n2238) );
  DFF_X1 matrix_mul_2D_reg_2__7__3_ ( .D(n9917), .CK(clk), .Q(
        matrix_mul_2D_2__7__3_), .QN(n2237) );
  DFF_X1 matrix_mul_2D_reg_2__7__4_ ( .D(n9913), .CK(clk), .Q(
        matrix_mul_2D_2__7__4_), .QN(n2236) );
  DFF_X1 matrix_mul_2D_reg_2__7__5_ ( .D(n9909), .CK(clk), .Q(
        matrix_mul_2D_2__7__5_), .QN(n2235) );
  DFF_X1 matrix_mul_2D_reg_2__7__6_ ( .D(n9905), .CK(clk), .Q(
        matrix_mul_2D_2__7__6_), .QN(n2234) );
  DFF_X1 matrix_mul_2D_reg_2__7__7_ ( .D(n9901), .CK(clk), .Q(
        matrix_mul_2D_2__7__7_), .QN(n2233) );
  DFF_X1 matrix_mul_2D_reg_2__7__8_ ( .D(n9897), .CK(clk), .Q(
        matrix_mul_2D_2__7__8_), .QN(n2232) );
  DFF_X1 matrix_mul_2D_reg_2__7__9_ ( .D(n9893), .CK(clk), .Q(
        matrix_mul_2D_2__7__9_), .QN(n2231) );
  DFF_X1 matrix_mul_2D_reg_2__7__10_ ( .D(n9889), .CK(clk), .Q(
        matrix_mul_2D_2__7__10_), .QN(n2230) );
  DFF_X1 matrix_mul_2D_reg_2__7__11_ ( .D(n9885), .CK(clk), .Q(
        matrix_mul_2D_2__7__11_), .QN(n2229) );
  DFF_X1 matrix_mul_2D_reg_2__7__12_ ( .D(n9881), .CK(clk), .Q(
        matrix_mul_2D_2__7__12_), .QN(n2228) );
  DFF_X1 matrix_mul_2D_reg_2__7__13_ ( .D(n9877), .CK(clk), .Q(
        matrix_mul_2D_2__7__13_), .QN(n2227) );
  DFF_X1 matrix_mul_2D_reg_2__7__14_ ( .D(n9873), .CK(clk), .Q(
        matrix_mul_2D_2__7__14_), .QN(n2226) );
  DFF_X1 matrix_mul_2D_reg_2__7__15_ ( .D(n9872), .CK(clk), .Q(
        matrix_mul_2D_2__7__15_), .QN(n17760) );
  DFF_X1 matrix_mul_2D_reg_2__7__16_ ( .D(n9871), .CK(clk), .Q(
        matrix_mul_2D_2__7__16_), .QN(n17758) );
  DFF_X1 matrix_mul_2D_reg_2__7__17_ ( .D(n9870), .CK(clk), .Q(
        matrix_mul_2D_2__7__17_), .QN(n17756) );
  DFF_X1 matrix_mul_2D_reg_2__7__18_ ( .D(n9869), .CK(clk), .Q(
        matrix_mul_2D_2__7__18_), .QN(n17754) );
  DFF_X1 matrix_mul_2D_reg_2__7__19_ ( .D(n9868), .CK(clk), .Q(
        matrix_mul_2D_2__7__19_), .QN(n17752) );
  DFF_X1 matrix_mul_2D_reg_2__7__20_ ( .D(n9867), .CK(clk), .Q(
        matrix_mul_2D_2__7__20_), .QN(n17750) );
  DFF_X1 matrix_mul_2D_reg_3__0__0_ ( .D(n9863), .CK(clk), .Q(
        matrix_mul_2D_3__0__0_), .QN(n2255) );
  DFF_X1 matrix_mul_2D_reg_3__0__1_ ( .D(n9858), .CK(clk), .Q(
        matrix_mul_2D_3__0__1_), .QN(n2254) );
  DFF_X1 matrix_mul_2D_reg_3__0__2_ ( .D(n9853), .CK(clk), .Q(
        matrix_mul_2D_3__0__2_), .QN(n2253) );
  DFF_X1 matrix_mul_2D_reg_3__0__3_ ( .D(n9848), .CK(clk), .Q(
        matrix_mul_2D_3__0__3_), .QN(n2252) );
  DFF_X1 matrix_mul_2D_reg_3__0__4_ ( .D(n9843), .CK(clk), .Q(
        matrix_mul_2D_3__0__4_), .QN(n2251) );
  DFF_X1 matrix_mul_2D_reg_3__0__5_ ( .D(n9838), .CK(clk), .Q(
        matrix_mul_2D_3__0__5_), .QN(n2250) );
  DFF_X1 matrix_mul_2D_reg_3__0__6_ ( .D(n9833), .CK(clk), .Q(
        matrix_mul_2D_3__0__6_), .QN(n2249) );
  DFF_X1 matrix_mul_2D_reg_3__0__7_ ( .D(n9828), .CK(clk), .Q(
        matrix_mul_2D_3__0__7_), .QN(n2248) );
  DFF_X1 matrix_mul_2D_reg_3__0__8_ ( .D(n9823), .CK(clk), .Q(
        matrix_mul_2D_3__0__8_), .QN(n2247) );
  DFF_X1 matrix_mul_2D_reg_3__0__9_ ( .D(n9818), .CK(clk), .Q(
        matrix_mul_2D_3__0__9_), .QN(n2246) );
  DFF_X1 matrix_mul_2D_reg_3__0__10_ ( .D(n9813), .CK(clk), .Q(
        matrix_mul_2D_3__0__10_), .QN(n2245) );
  DFF_X1 matrix_mul_2D_reg_3__0__11_ ( .D(n9808), .CK(clk), .Q(
        matrix_mul_2D_3__0__11_), .QN(n2244) );
  DFF_X1 matrix_mul_2D_reg_3__0__12_ ( .D(n9803), .CK(clk), .Q(
        matrix_mul_2D_3__0__12_), .QN(n2243) );
  DFF_X1 matrix_mul_2D_reg_3__0__13_ ( .D(n9798), .CK(clk), .Q(
        matrix_mul_2D_3__0__13_), .QN(n2242) );
  DFF_X1 matrix_mul_2D_reg_3__0__14_ ( .D(n9793), .CK(clk), .Q(
        matrix_mul_2D_3__0__14_), .QN(n2241) );
  DFF_X1 matrix_mul_2D_reg_3__0__15_ ( .D(n9792), .CK(clk), .Q(
        matrix_mul_2D_3__0__15_), .QN(n17748) );
  DFF_X1 matrix_mul_2D_reg_3__0__16_ ( .D(n9791), .CK(clk), .Q(
        matrix_mul_2D_3__0__16_), .QN(n17746) );
  DFF_X1 matrix_mul_2D_reg_3__0__17_ ( .D(n9790), .CK(clk), .Q(
        matrix_mul_2D_3__0__17_), .QN(n17744) );
  DFF_X1 matrix_mul_2D_reg_3__0__18_ ( .D(n9789), .CK(clk), .Q(
        matrix_mul_2D_3__0__18_), .QN(n17742) );
  DFF_X1 matrix_mul_2D_reg_3__0__19_ ( .D(n9788), .CK(clk), .Q(
        matrix_mul_2D_3__0__19_), .QN(n17740) );
  DFF_X1 matrix_mul_2D_reg_3__0__20_ ( .D(n9787), .CK(clk), .Q(
        matrix_mul_2D_3__0__20_), .QN(n17738) );
  DFF_X1 matrix_mul_2D_reg_3__1__0_ ( .D(n9783), .CK(clk), .Q(
        matrix_mul_2D_3__1__0_), .QN(n2270) );
  DFF_X1 matrix_mul_2D_reg_3__1__1_ ( .D(n9778), .CK(clk), .Q(
        matrix_mul_2D_3__1__1_), .QN(n2269) );
  DFF_X1 matrix_mul_2D_reg_3__1__2_ ( .D(n9773), .CK(clk), .Q(
        matrix_mul_2D_3__1__2_), .QN(n2268) );
  DFF_X1 matrix_mul_2D_reg_3__1__3_ ( .D(n9768), .CK(clk), .Q(
        matrix_mul_2D_3__1__3_), .QN(n2267) );
  DFF_X1 matrix_mul_2D_reg_3__1__4_ ( .D(n9763), .CK(clk), .Q(
        matrix_mul_2D_3__1__4_), .QN(n2266) );
  DFF_X1 matrix_mul_2D_reg_3__1__5_ ( .D(n9758), .CK(clk), .Q(
        matrix_mul_2D_3__1__5_), .QN(n2265) );
  DFF_X1 matrix_mul_2D_reg_3__1__6_ ( .D(n9753), .CK(clk), .Q(
        matrix_mul_2D_3__1__6_), .QN(n2264) );
  DFF_X1 matrix_mul_2D_reg_3__1__7_ ( .D(n9748), .CK(clk), .Q(
        matrix_mul_2D_3__1__7_), .QN(n2263) );
  DFF_X1 matrix_mul_2D_reg_3__1__8_ ( .D(n9743), .CK(clk), .Q(
        matrix_mul_2D_3__1__8_), .QN(n2262) );
  DFF_X1 matrix_mul_2D_reg_3__1__9_ ( .D(n9738), .CK(clk), .Q(
        matrix_mul_2D_3__1__9_), .QN(n2261) );
  DFF_X1 matrix_mul_2D_reg_3__1__10_ ( .D(n9733), .CK(clk), .Q(
        matrix_mul_2D_3__1__10_), .QN(n2260) );
  DFF_X1 matrix_mul_2D_reg_3__1__11_ ( .D(n9728), .CK(clk), .Q(
        matrix_mul_2D_3__1__11_), .QN(n2259) );
  DFF_X1 matrix_mul_2D_reg_3__1__12_ ( .D(n9723), .CK(clk), .Q(
        matrix_mul_2D_3__1__12_), .QN(n2258) );
  DFF_X1 matrix_mul_2D_reg_3__1__13_ ( .D(n9718), .CK(clk), .Q(
        matrix_mul_2D_3__1__13_), .QN(n2257) );
  DFF_X1 matrix_mul_2D_reg_3__1__14_ ( .D(n9713), .CK(clk), .Q(
        matrix_mul_2D_3__1__14_), .QN(n2256) );
  DFF_X1 matrix_mul_2D_reg_3__1__15_ ( .D(n9712), .CK(clk), .Q(
        matrix_mul_2D_3__1__15_), .QN(n17736) );
  DFF_X1 matrix_mul_2D_reg_3__1__16_ ( .D(n9711), .CK(clk), .Q(
        matrix_mul_2D_3__1__16_), .QN(n17734) );
  DFF_X1 matrix_mul_2D_reg_3__1__17_ ( .D(n9710), .CK(clk), .Q(
        matrix_mul_2D_3__1__17_), .QN(n17732) );
  DFF_X1 matrix_mul_2D_reg_3__1__18_ ( .D(n9709), .CK(clk), .Q(
        matrix_mul_2D_3__1__18_), .QN(n17730) );
  DFF_X1 matrix_mul_2D_reg_3__1__19_ ( .D(n9708), .CK(clk), .Q(
        matrix_mul_2D_3__1__19_), .QN(n17728) );
  DFF_X1 matrix_mul_2D_reg_3__1__20_ ( .D(n9707), .CK(clk), .Q(
        matrix_mul_2D_3__1__20_), .QN(n17726) );
  DFF_X1 matrix_mul_2D_reg_3__2__0_ ( .D(n9703), .CK(clk), .Q(
        matrix_mul_2D_3__2__0_), .QN(n2285) );
  DFF_X1 matrix_mul_2D_reg_3__2__1_ ( .D(n9698), .CK(clk), .Q(
        matrix_mul_2D_3__2__1_), .QN(n2284) );
  DFF_X1 matrix_mul_2D_reg_3__2__2_ ( .D(n9693), .CK(clk), .Q(
        matrix_mul_2D_3__2__2_), .QN(n2283) );
  DFF_X1 matrix_mul_2D_reg_3__2__3_ ( .D(n9688), .CK(clk), .Q(
        matrix_mul_2D_3__2__3_), .QN(n2282) );
  DFF_X1 matrix_mul_2D_reg_3__2__4_ ( .D(n9683), .CK(clk), .Q(
        matrix_mul_2D_3__2__4_), .QN(n2281) );
  DFF_X1 matrix_mul_2D_reg_3__2__5_ ( .D(n9678), .CK(clk), .Q(
        matrix_mul_2D_3__2__5_), .QN(n2280) );
  DFF_X1 matrix_mul_2D_reg_3__2__6_ ( .D(n9673), .CK(clk), .Q(
        matrix_mul_2D_3__2__6_), .QN(n2279) );
  DFF_X1 matrix_mul_2D_reg_3__2__7_ ( .D(n9668), .CK(clk), .Q(
        matrix_mul_2D_3__2__7_), .QN(n2278) );
  DFF_X1 matrix_mul_2D_reg_3__2__8_ ( .D(n9663), .CK(clk), .Q(
        matrix_mul_2D_3__2__8_), .QN(n2277) );
  DFF_X1 matrix_mul_2D_reg_3__2__9_ ( .D(n9658), .CK(clk), .Q(
        matrix_mul_2D_3__2__9_), .QN(n2276) );
  DFF_X1 matrix_mul_2D_reg_3__2__10_ ( .D(n9653), .CK(clk), .Q(
        matrix_mul_2D_3__2__10_), .QN(n2275) );
  DFF_X1 matrix_mul_2D_reg_3__2__11_ ( .D(n9648), .CK(clk), .Q(
        matrix_mul_2D_3__2__11_), .QN(n2274) );
  DFF_X1 matrix_mul_2D_reg_3__2__12_ ( .D(n9643), .CK(clk), .Q(
        matrix_mul_2D_3__2__12_), .QN(n2273) );
  DFF_X1 matrix_mul_2D_reg_3__2__13_ ( .D(n9638), .CK(clk), .Q(
        matrix_mul_2D_3__2__13_), .QN(n2272) );
  DFF_X1 matrix_mul_2D_reg_3__2__14_ ( .D(n9633), .CK(clk), .Q(
        matrix_mul_2D_3__2__14_), .QN(n2271) );
  DFF_X1 matrix_mul_2D_reg_3__2__15_ ( .D(n9632), .CK(clk), .Q(
        matrix_mul_2D_3__2__15_), .QN(n17724) );
  DFF_X1 matrix_mul_2D_reg_3__2__16_ ( .D(n9631), .CK(clk), .Q(
        matrix_mul_2D_3__2__16_), .QN(n17722) );
  DFF_X1 matrix_mul_2D_reg_3__2__17_ ( .D(n9630), .CK(clk), .Q(
        matrix_mul_2D_3__2__17_), .QN(n17720) );
  DFF_X1 matrix_mul_2D_reg_3__2__18_ ( .D(n9629), .CK(clk), .Q(
        matrix_mul_2D_3__2__18_), .QN(n17718) );
  DFF_X1 matrix_mul_2D_reg_3__2__19_ ( .D(n9628), .CK(clk), .Q(
        matrix_mul_2D_3__2__19_), .QN(n17716) );
  DFF_X1 matrix_mul_2D_reg_3__2__20_ ( .D(n9627), .CK(clk), .Q(
        matrix_mul_2D_3__2__20_), .QN(n17714) );
  DFF_X1 matrix_mul_2D_reg_3__3__0_ ( .D(n9622), .CK(clk), .Q(
        matrix_mul_2D_3__3__0_), .QN(n2306) );
  DFF_X1 matrix_mul_2D_reg_3__3__1_ ( .D(n9618), .CK(clk), .Q(
        matrix_mul_2D_3__3__1_), .QN(n2305) );
  DFF_X1 matrix_mul_2D_reg_3__3__2_ ( .D(n9614), .CK(clk), .Q(
        matrix_mul_2D_3__3__2_), .QN(n2304) );
  DFF_X1 matrix_mul_2D_reg_3__3__3_ ( .D(n9610), .CK(clk), .Q(
        matrix_mul_2D_3__3__3_), .QN(n2303) );
  DFF_X1 matrix_mul_2D_reg_3__3__4_ ( .D(n9606), .CK(clk), .Q(
        matrix_mul_2D_3__3__4_), .QN(n2302) );
  DFF_X1 matrix_mul_2D_reg_3__3__5_ ( .D(n9602), .CK(clk), .Q(
        matrix_mul_2D_3__3__5_), .QN(n2301) );
  DFF_X1 matrix_mul_2D_reg_3__3__6_ ( .D(n9598), .CK(clk), .Q(
        matrix_mul_2D_3__3__6_), .QN(n2300) );
  DFF_X1 matrix_mul_2D_reg_3__3__7_ ( .D(n9594), .CK(clk), .Q(
        matrix_mul_2D_3__3__7_), .QN(n2299) );
  DFF_X1 matrix_mul_2D_reg_3__3__8_ ( .D(n9590), .CK(clk), .Q(
        matrix_mul_2D_3__3__8_), .QN(n2298) );
  DFF_X1 matrix_mul_2D_reg_3__3__9_ ( .D(n9586), .CK(clk), .Q(
        matrix_mul_2D_3__3__9_), .QN(n2297) );
  DFF_X1 matrix_mul_2D_reg_3__3__10_ ( .D(n9582), .CK(clk), .Q(
        matrix_mul_2D_3__3__10_), .QN(n2296) );
  DFF_X1 matrix_mul_2D_reg_3__3__11_ ( .D(n9578), .CK(clk), .Q(
        matrix_mul_2D_3__3__11_), .QN(n2295) );
  DFF_X1 matrix_mul_2D_reg_3__3__12_ ( .D(n9574), .CK(clk), .Q(
        matrix_mul_2D_3__3__12_), .QN(n2294) );
  DFF_X1 matrix_mul_2D_reg_3__3__13_ ( .D(n9570), .CK(clk), .Q(
        matrix_mul_2D_3__3__13_), .QN(n2293) );
  DFF_X1 matrix_mul_2D_reg_3__3__14_ ( .D(n9566), .CK(clk), .Q(
        matrix_mul_2D_3__3__14_), .QN(n2292) );
  DFF_X1 matrix_mul_2D_reg_3__3__15_ ( .D(n9565), .CK(clk), .Q(
        matrix_mul_2D_3__3__15_), .QN(n17712) );
  DFF_X1 matrix_mul_2D_reg_3__3__16_ ( .D(n9564), .CK(clk), .Q(
        matrix_mul_2D_3__3__16_), .QN(n17710) );
  DFF_X1 matrix_mul_2D_reg_3__3__17_ ( .D(n9563), .CK(clk), .Q(
        matrix_mul_2D_3__3__17_), .QN(n17708) );
  DFF_X1 matrix_mul_2D_reg_3__3__18_ ( .D(n9562), .CK(clk), .Q(
        matrix_mul_2D_3__3__18_), .QN(n17706) );
  DFF_X1 matrix_mul_2D_reg_3__3__19_ ( .D(n9561), .CK(clk), .Q(
        matrix_mul_2D_3__3__19_), .QN(n17704) );
  DFF_X1 matrix_mul_2D_reg_3__3__20_ ( .D(n9560), .CK(clk), .Q(
        matrix_mul_2D_3__3__20_), .QN(n17702) );
  DFF_X1 matrix_mul_2D_reg_3__4__0_ ( .D(n9555), .CK(clk), .Q(
        matrix_mul_2D_3__4__0_), .QN(n2321) );
  DFF_X1 matrix_mul_2D_reg_3__4__1_ ( .D(n9551), .CK(clk), .Q(
        matrix_mul_2D_3__4__1_), .QN(n2320) );
  DFF_X1 matrix_mul_2D_reg_3__4__2_ ( .D(n9547), .CK(clk), .Q(
        matrix_mul_2D_3__4__2_), .QN(n2319) );
  DFF_X1 matrix_mul_2D_reg_3__4__3_ ( .D(n9543), .CK(clk), .Q(
        matrix_mul_2D_3__4__3_), .QN(n2318) );
  DFF_X1 matrix_mul_2D_reg_3__4__4_ ( .D(n9539), .CK(clk), .Q(
        matrix_mul_2D_3__4__4_), .QN(n2317) );
  DFF_X1 matrix_mul_2D_reg_3__4__5_ ( .D(n9535), .CK(clk), .Q(
        matrix_mul_2D_3__4__5_), .QN(n2316) );
  DFF_X1 matrix_mul_2D_reg_3__4__6_ ( .D(n9531), .CK(clk), .Q(
        matrix_mul_2D_3__4__6_), .QN(n2315) );
  DFF_X1 matrix_mul_2D_reg_3__4__7_ ( .D(n9527), .CK(clk), .Q(
        matrix_mul_2D_3__4__7_), .QN(n2314) );
  DFF_X1 matrix_mul_2D_reg_3__4__8_ ( .D(n9523), .CK(clk), .Q(
        matrix_mul_2D_3__4__8_), .QN(n2313) );
  DFF_X1 matrix_mul_2D_reg_3__4__9_ ( .D(n9519), .CK(clk), .Q(
        matrix_mul_2D_3__4__9_), .QN(n2312) );
  DFF_X1 matrix_mul_2D_reg_3__4__10_ ( .D(n9515), .CK(clk), .Q(
        matrix_mul_2D_3__4__10_), .QN(n2311) );
  DFF_X1 matrix_mul_2D_reg_3__4__11_ ( .D(n9511), .CK(clk), .Q(
        matrix_mul_2D_3__4__11_), .QN(n2310) );
  DFF_X1 matrix_mul_2D_reg_3__4__12_ ( .D(n9507), .CK(clk), .Q(
        matrix_mul_2D_3__4__12_), .QN(n2309) );
  DFF_X1 matrix_mul_2D_reg_3__4__13_ ( .D(n9503), .CK(clk), .Q(
        matrix_mul_2D_3__4__13_), .QN(n2308) );
  DFF_X1 matrix_mul_2D_reg_3__4__14_ ( .D(n9499), .CK(clk), .Q(
        matrix_mul_2D_3__4__14_), .QN(n2307) );
  DFF_X1 matrix_mul_2D_reg_3__4__15_ ( .D(n9498), .CK(clk), .Q(
        matrix_mul_2D_3__4__15_), .QN(n17700) );
  DFF_X1 matrix_mul_2D_reg_3__4__16_ ( .D(n9497), .CK(clk), .Q(
        matrix_mul_2D_3__4__16_), .QN(n17698) );
  DFF_X1 matrix_mul_2D_reg_3__4__17_ ( .D(n9496), .CK(clk), .Q(
        matrix_mul_2D_3__4__17_), .QN(n17696) );
  DFF_X1 matrix_mul_2D_reg_3__4__18_ ( .D(n9495), .CK(clk), .Q(
        matrix_mul_2D_3__4__18_), .QN(n17694) );
  DFF_X1 matrix_mul_2D_reg_3__4__19_ ( .D(n9494), .CK(clk), .Q(
        matrix_mul_2D_3__4__19_), .QN(n17692) );
  DFF_X1 matrix_mul_2D_reg_3__4__20_ ( .D(n9493), .CK(clk), .Q(
        matrix_mul_2D_3__4__20_), .QN(n17690) );
  DFF_X1 matrix_mul_2D_reg_3__5__0_ ( .D(n9489), .CK(clk), .Q(
        matrix_mul_2D_3__5__0_), .QN(n2336) );
  DFF_X1 matrix_mul_2D_reg_3__5__1_ ( .D(n9484), .CK(clk), .Q(
        matrix_mul_2D_3__5__1_), .QN(n2335) );
  DFF_X1 matrix_mul_2D_reg_3__5__2_ ( .D(n9479), .CK(clk), .Q(
        matrix_mul_2D_3__5__2_), .QN(n2334) );
  DFF_X1 matrix_mul_2D_reg_3__5__3_ ( .D(n9474), .CK(clk), .Q(
        matrix_mul_2D_3__5__3_), .QN(n2333) );
  DFF_X1 matrix_mul_2D_reg_3__5__4_ ( .D(n9469), .CK(clk), .Q(
        matrix_mul_2D_3__5__4_), .QN(n2332) );
  DFF_X1 matrix_mul_2D_reg_3__5__5_ ( .D(n9464), .CK(clk), .Q(
        matrix_mul_2D_3__5__5_), .QN(n2331) );
  DFF_X1 matrix_mul_2D_reg_3__5__6_ ( .D(n9459), .CK(clk), .Q(
        matrix_mul_2D_3__5__6_), .QN(n2330) );
  DFF_X1 matrix_mul_2D_reg_3__5__7_ ( .D(n9454), .CK(clk), .Q(
        matrix_mul_2D_3__5__7_), .QN(n2329) );
  DFF_X1 matrix_mul_2D_reg_3__5__8_ ( .D(n9449), .CK(clk), .Q(
        matrix_mul_2D_3__5__8_), .QN(n2328) );
  DFF_X1 matrix_mul_2D_reg_3__5__9_ ( .D(n9444), .CK(clk), .Q(
        matrix_mul_2D_3__5__9_), .QN(n2327) );
  DFF_X1 matrix_mul_2D_reg_3__5__10_ ( .D(n9439), .CK(clk), .Q(
        matrix_mul_2D_3__5__10_), .QN(n2326) );
  DFF_X1 matrix_mul_2D_reg_3__5__11_ ( .D(n9434), .CK(clk), .Q(
        matrix_mul_2D_3__5__11_), .QN(n2325) );
  DFF_X1 matrix_mul_2D_reg_3__5__12_ ( .D(n9429), .CK(clk), .Q(
        matrix_mul_2D_3__5__12_), .QN(n2324) );
  DFF_X1 matrix_mul_2D_reg_3__5__13_ ( .D(n9424), .CK(clk), .Q(
        matrix_mul_2D_3__5__13_), .QN(n2323) );
  DFF_X1 matrix_mul_2D_reg_3__5__14_ ( .D(n9419), .CK(clk), .Q(
        matrix_mul_2D_3__5__14_), .QN(n2322) );
  DFF_X1 matrix_mul_2D_reg_3__5__15_ ( .D(n9418), .CK(clk), .Q(
        matrix_mul_2D_3__5__15_), .QN(n17688) );
  DFF_X1 matrix_mul_2D_reg_3__5__16_ ( .D(n9417), .CK(clk), .Q(
        matrix_mul_2D_3__5__16_), .QN(n17686) );
  DFF_X1 matrix_mul_2D_reg_3__5__17_ ( .D(n9416), .CK(clk), .Q(
        matrix_mul_2D_3__5__17_), .QN(n17684) );
  DFF_X1 matrix_mul_2D_reg_3__5__18_ ( .D(n9415), .CK(clk), .Q(
        matrix_mul_2D_3__5__18_), .QN(n17682) );
  DFF_X1 matrix_mul_2D_reg_3__5__19_ ( .D(n9414), .CK(clk), .Q(
        matrix_mul_2D_3__5__19_), .QN(n17680) );
  DFF_X1 matrix_mul_2D_reg_3__5__20_ ( .D(n9413), .CK(clk), .Q(
        matrix_mul_2D_3__5__20_), .QN(n17678) );
  DFF_X1 matrix_mul_2D_reg_3__6__0_ ( .D(n9409), .CK(clk), .Q(
        matrix_mul_2D_3__6__0_), .QN(n2351) );
  DFF_X1 matrix_mul_2D_reg_3__6__1_ ( .D(n9404), .CK(clk), .Q(
        matrix_mul_2D_3__6__1_), .QN(n2350) );
  DFF_X1 matrix_mul_2D_reg_3__6__2_ ( .D(n9399), .CK(clk), .Q(
        matrix_mul_2D_3__6__2_), .QN(n2349) );
  DFF_X1 matrix_mul_2D_reg_3__6__3_ ( .D(n9394), .CK(clk), .Q(
        matrix_mul_2D_3__6__3_), .QN(n2348) );
  DFF_X1 matrix_mul_2D_reg_3__6__4_ ( .D(n9389), .CK(clk), .Q(
        matrix_mul_2D_3__6__4_), .QN(n2347) );
  DFF_X1 matrix_mul_2D_reg_3__6__5_ ( .D(n9384), .CK(clk), .Q(
        matrix_mul_2D_3__6__5_), .QN(n2346) );
  DFF_X1 matrix_mul_2D_reg_3__6__6_ ( .D(n9379), .CK(clk), .Q(
        matrix_mul_2D_3__6__6_), .QN(n2345) );
  DFF_X1 matrix_mul_2D_reg_3__6__7_ ( .D(n9374), .CK(clk), .Q(
        matrix_mul_2D_3__6__7_), .QN(n2344) );
  DFF_X1 matrix_mul_2D_reg_3__6__8_ ( .D(n9369), .CK(clk), .Q(
        matrix_mul_2D_3__6__8_), .QN(n2343) );
  DFF_X1 matrix_mul_2D_reg_3__6__9_ ( .D(n9364), .CK(clk), .Q(
        matrix_mul_2D_3__6__9_), .QN(n2342) );
  DFF_X1 matrix_mul_2D_reg_3__6__10_ ( .D(n9359), .CK(clk), .Q(
        matrix_mul_2D_3__6__10_), .QN(n2341) );
  DFF_X1 matrix_mul_2D_reg_3__6__11_ ( .D(n9354), .CK(clk), .Q(
        matrix_mul_2D_3__6__11_), .QN(n2340) );
  DFF_X1 matrix_mul_2D_reg_3__6__12_ ( .D(n9349), .CK(clk), .Q(
        matrix_mul_2D_3__6__12_), .QN(n2339) );
  DFF_X1 matrix_mul_2D_reg_3__6__13_ ( .D(n9344), .CK(clk), .Q(
        matrix_mul_2D_3__6__13_), .QN(n2338) );
  DFF_X1 matrix_mul_2D_reg_3__6__14_ ( .D(n9339), .CK(clk), .Q(
        matrix_mul_2D_3__6__14_), .QN(n2337) );
  DFF_X1 matrix_mul_2D_reg_3__6__15_ ( .D(n9338), .CK(clk), .Q(
        matrix_mul_2D_3__6__15_), .QN(n17676) );
  DFF_X1 matrix_mul_2D_reg_3__6__16_ ( .D(n9337), .CK(clk), .Q(
        matrix_mul_2D_3__6__16_), .QN(n17674) );
  DFF_X1 matrix_mul_2D_reg_3__6__17_ ( .D(n9336), .CK(clk), .Q(
        matrix_mul_2D_3__6__17_), .QN(n17672) );
  DFF_X1 matrix_mul_2D_reg_3__6__18_ ( .D(n9335), .CK(clk), .Q(
        matrix_mul_2D_3__6__18_), .QN(n17670) );
  DFF_X1 matrix_mul_2D_reg_3__6__19_ ( .D(n9334), .CK(clk), .Q(
        matrix_mul_2D_3__6__19_), .QN(n17668) );
  DFF_X1 matrix_mul_2D_reg_3__6__20_ ( .D(n9333), .CK(clk), .Q(
        matrix_mul_2D_3__6__20_), .QN(n17666) );
  DFF_X1 matrix_mul_2D_reg_3__7__0_ ( .D(n9329), .CK(clk), .Q(
        matrix_mul_2D_3__7__0_), .QN(n2366) );
  DFF_X1 matrix_mul_2D_reg_3__7__1_ ( .D(n9324), .CK(clk), .Q(
        matrix_mul_2D_3__7__1_), .QN(n2365) );
  DFF_X1 matrix_mul_2D_reg_3__7__2_ ( .D(n9319), .CK(clk), .Q(
        matrix_mul_2D_3__7__2_), .QN(n2364) );
  DFF_X1 matrix_mul_2D_reg_3__7__3_ ( .D(n9314), .CK(clk), .Q(
        matrix_mul_2D_3__7__3_), .QN(n2363) );
  DFF_X1 matrix_mul_2D_reg_3__7__4_ ( .D(n9309), .CK(clk), .Q(
        matrix_mul_2D_3__7__4_), .QN(n2362) );
  DFF_X1 matrix_mul_2D_reg_3__7__5_ ( .D(n9304), .CK(clk), .Q(
        matrix_mul_2D_3__7__5_), .QN(n2361) );
  DFF_X1 matrix_mul_2D_reg_3__7__6_ ( .D(n9299), .CK(clk), .Q(
        matrix_mul_2D_3__7__6_), .QN(n2360) );
  DFF_X1 matrix_mul_2D_reg_3__7__7_ ( .D(n9294), .CK(clk), .Q(
        matrix_mul_2D_3__7__7_), .QN(n2359) );
  DFF_X1 matrix_mul_2D_reg_3__7__8_ ( .D(n9289), .CK(clk), .Q(
        matrix_mul_2D_3__7__8_), .QN(n2358) );
  DFF_X1 matrix_mul_2D_reg_3__7__9_ ( .D(n9284), .CK(clk), .Q(
        matrix_mul_2D_3__7__9_), .QN(n2357) );
  DFF_X1 matrix_mul_2D_reg_3__7__10_ ( .D(n9279), .CK(clk), .Q(
        matrix_mul_2D_3__7__10_), .QN(n2356) );
  DFF_X1 matrix_mul_2D_reg_3__7__11_ ( .D(n9274), .CK(clk), .Q(
        matrix_mul_2D_3__7__11_), .QN(n2355) );
  DFF_X1 matrix_mul_2D_reg_3__7__12_ ( .D(n9269), .CK(clk), .Q(
        matrix_mul_2D_3__7__12_), .QN(n2354) );
  DFF_X1 matrix_mul_2D_reg_3__7__13_ ( .D(n9264), .CK(clk), .Q(
        matrix_mul_2D_3__7__13_), .QN(n2353) );
  DFF_X1 matrix_mul_2D_reg_3__7__14_ ( .D(n9259), .CK(clk), .Q(
        matrix_mul_2D_3__7__14_), .QN(n2352) );
  DFF_X1 matrix_mul_2D_reg_3__7__15_ ( .D(n9258), .CK(clk), .Q(
        matrix_mul_2D_3__7__15_), .QN(n17664) );
  DFF_X1 matrix_mul_2D_reg_3__7__16_ ( .D(n9257), .CK(clk), .Q(
        matrix_mul_2D_3__7__16_), .QN(n17662) );
  DFF_X1 matrix_mul_2D_reg_3__7__17_ ( .D(n9256), .CK(clk), .Q(
        matrix_mul_2D_3__7__17_), .QN(n17660) );
  DFF_X1 matrix_mul_2D_reg_3__7__18_ ( .D(n9255), .CK(clk), .Q(
        matrix_mul_2D_3__7__18_), .QN(n17658) );
  DFF_X1 matrix_mul_2D_reg_3__7__19_ ( .D(n9254), .CK(clk), .Q(
        matrix_mul_2D_3__7__19_), .QN(n17656) );
  DFF_X1 matrix_mul_2D_reg_3__7__20_ ( .D(n9253), .CK(clk), .Q(
        matrix_mul_2D_3__7__20_), .QN(n17654) );
  DFF_X1 matrix_mul_2D_reg_4__0__0_ ( .D(n9249), .CK(clk), .Q(
        matrix_mul_2D_4__0__0_), .QN(n2381) );
  DFF_X1 matrix_mul_2D_reg_4__0__1_ ( .D(n9244), .CK(clk), .Q(
        matrix_mul_2D_4__0__1_), .QN(n2380) );
  DFF_X1 matrix_mul_2D_reg_4__0__2_ ( .D(n9239), .CK(clk), .Q(
        matrix_mul_2D_4__0__2_), .QN(n2379) );
  DFF_X1 matrix_mul_2D_reg_4__0__3_ ( .D(n9234), .CK(clk), .Q(
        matrix_mul_2D_4__0__3_), .QN(n2378) );
  DFF_X1 matrix_mul_2D_reg_4__0__4_ ( .D(n9229), .CK(clk), .Q(
        matrix_mul_2D_4__0__4_), .QN(n2377) );
  DFF_X1 matrix_mul_2D_reg_4__0__5_ ( .D(n9224), .CK(clk), .Q(
        matrix_mul_2D_4__0__5_), .QN(n2376) );
  DFF_X1 matrix_mul_2D_reg_4__0__6_ ( .D(n9219), .CK(clk), .Q(
        matrix_mul_2D_4__0__6_), .QN(n2375) );
  DFF_X1 matrix_mul_2D_reg_4__0__7_ ( .D(n9214), .CK(clk), .Q(
        matrix_mul_2D_4__0__7_), .QN(n2374) );
  DFF_X1 matrix_mul_2D_reg_4__0__8_ ( .D(n9209), .CK(clk), .Q(
        matrix_mul_2D_4__0__8_), .QN(n2373) );
  DFF_X1 matrix_mul_2D_reg_4__0__9_ ( .D(n9204), .CK(clk), .Q(
        matrix_mul_2D_4__0__9_), .QN(n2372) );
  DFF_X1 matrix_mul_2D_reg_4__0__10_ ( .D(n9199), .CK(clk), .Q(
        matrix_mul_2D_4__0__10_), .QN(n2371) );
  DFF_X1 matrix_mul_2D_reg_4__0__11_ ( .D(n9194), .CK(clk), .Q(
        matrix_mul_2D_4__0__11_), .QN(n2370) );
  DFF_X1 matrix_mul_2D_reg_4__0__12_ ( .D(n9189), .CK(clk), .Q(
        matrix_mul_2D_4__0__12_), .QN(n2369) );
  DFF_X1 matrix_mul_2D_reg_4__0__13_ ( .D(n9184), .CK(clk), .Q(
        matrix_mul_2D_4__0__13_), .QN(n2368) );
  DFF_X1 matrix_mul_2D_reg_4__0__14_ ( .D(n9179), .CK(clk), .Q(
        matrix_mul_2D_4__0__14_), .QN(n2367) );
  DFF_X1 matrix_mul_2D_reg_4__0__15_ ( .D(n9178), .CK(clk), .Q(
        matrix_mul_2D_4__0__15_), .QN(n17652) );
  DFF_X1 matrix_mul_2D_reg_4__0__16_ ( .D(n9177), .CK(clk), .Q(
        matrix_mul_2D_4__0__16_), .QN(n17650) );
  DFF_X1 matrix_mul_2D_reg_4__0__17_ ( .D(n9176), .CK(clk), .Q(
        matrix_mul_2D_4__0__17_), .QN(n17648) );
  DFF_X1 matrix_mul_2D_reg_4__0__18_ ( .D(n9175), .CK(clk), .Q(
        matrix_mul_2D_4__0__18_), .QN(n17646) );
  DFF_X1 matrix_mul_2D_reg_4__0__19_ ( .D(n9174), .CK(clk), .Q(
        matrix_mul_2D_4__0__19_), .QN(n17644) );
  DFF_X1 matrix_mul_2D_reg_4__0__20_ ( .D(n9173), .CK(clk), .Q(
        matrix_mul_2D_4__0__20_), .QN(n17642) );
  DFF_X1 matrix_mul_2D_reg_4__1__0_ ( .D(n9169), .CK(clk), .Q(
        matrix_mul_2D_4__1__0_), .QN(n2396) );
  DFF_X1 matrix_mul_2D_reg_4__1__1_ ( .D(n9164), .CK(clk), .Q(
        matrix_mul_2D_4__1__1_), .QN(n2395) );
  DFF_X1 matrix_mul_2D_reg_4__1__2_ ( .D(n9159), .CK(clk), .Q(
        matrix_mul_2D_4__1__2_), .QN(n2394) );
  DFF_X1 matrix_mul_2D_reg_4__1__3_ ( .D(n9154), .CK(clk), .Q(
        matrix_mul_2D_4__1__3_), .QN(n2393) );
  DFF_X1 matrix_mul_2D_reg_4__1__4_ ( .D(n9149), .CK(clk), .Q(
        matrix_mul_2D_4__1__4_), .QN(n2392) );
  DFF_X1 matrix_mul_2D_reg_4__1__5_ ( .D(n9144), .CK(clk), .Q(
        matrix_mul_2D_4__1__5_), .QN(n2391) );
  DFF_X1 matrix_mul_2D_reg_4__1__6_ ( .D(n9139), .CK(clk), .Q(
        matrix_mul_2D_4__1__6_), .QN(n2390) );
  DFF_X1 matrix_mul_2D_reg_4__1__7_ ( .D(n9134), .CK(clk), .Q(
        matrix_mul_2D_4__1__7_), .QN(n2389) );
  DFF_X1 matrix_mul_2D_reg_4__1__8_ ( .D(n9129), .CK(clk), .Q(
        matrix_mul_2D_4__1__8_), .QN(n2388) );
  DFF_X1 matrix_mul_2D_reg_4__1__9_ ( .D(n9124), .CK(clk), .Q(
        matrix_mul_2D_4__1__9_), .QN(n2387) );
  DFF_X1 matrix_mul_2D_reg_4__1__10_ ( .D(n9119), .CK(clk), .Q(
        matrix_mul_2D_4__1__10_), .QN(n2386) );
  DFF_X1 matrix_mul_2D_reg_4__1__11_ ( .D(n9114), .CK(clk), .Q(
        matrix_mul_2D_4__1__11_), .QN(n2385) );
  DFF_X1 matrix_mul_2D_reg_4__1__12_ ( .D(n9109), .CK(clk), .Q(
        matrix_mul_2D_4__1__12_), .QN(n2384) );
  DFF_X1 matrix_mul_2D_reg_4__1__13_ ( .D(n9104), .CK(clk), .Q(
        matrix_mul_2D_4__1__13_), .QN(n2383) );
  DFF_X1 matrix_mul_2D_reg_4__1__14_ ( .D(n9099), .CK(clk), .Q(
        matrix_mul_2D_4__1__14_), .QN(n2382) );
  DFF_X1 matrix_mul_2D_reg_4__1__15_ ( .D(n9098), .CK(clk), .Q(
        matrix_mul_2D_4__1__15_), .QN(n17640) );
  DFF_X1 matrix_mul_2D_reg_4__1__16_ ( .D(n9097), .CK(clk), .Q(
        matrix_mul_2D_4__1__16_), .QN(n17638) );
  DFF_X1 matrix_mul_2D_reg_4__1__17_ ( .D(n9096), .CK(clk), .Q(
        matrix_mul_2D_4__1__17_), .QN(n17636) );
  DFF_X1 matrix_mul_2D_reg_4__1__18_ ( .D(n9095), .CK(clk), .Q(
        matrix_mul_2D_4__1__18_), .QN(n17634) );
  DFF_X1 matrix_mul_2D_reg_4__1__19_ ( .D(n9094), .CK(clk), .Q(
        matrix_mul_2D_4__1__19_), .QN(n17632) );
  DFF_X1 matrix_mul_2D_reg_4__1__20_ ( .D(n9093), .CK(clk), .Q(
        matrix_mul_2D_4__1__20_), .QN(n17630) );
  DFF_X1 matrix_mul_2D_reg_4__2__0_ ( .D(n9089), .CK(clk), .Q(
        matrix_mul_2D_4__2__0_), .QN(n2411) );
  DFF_X1 matrix_mul_2D_reg_4__2__1_ ( .D(n9084), .CK(clk), .Q(
        matrix_mul_2D_4__2__1_), .QN(n2410) );
  DFF_X1 matrix_mul_2D_reg_4__2__2_ ( .D(n9079), .CK(clk), .Q(
        matrix_mul_2D_4__2__2_), .QN(n2409) );
  DFF_X1 matrix_mul_2D_reg_4__2__3_ ( .D(n9074), .CK(clk), .Q(
        matrix_mul_2D_4__2__3_), .QN(n2408) );
  DFF_X1 matrix_mul_2D_reg_4__2__4_ ( .D(n9069), .CK(clk), .Q(
        matrix_mul_2D_4__2__4_), .QN(n2407) );
  DFF_X1 matrix_mul_2D_reg_4__2__5_ ( .D(n9064), .CK(clk), .Q(
        matrix_mul_2D_4__2__5_), .QN(n2406) );
  DFF_X1 matrix_mul_2D_reg_4__2__6_ ( .D(n9059), .CK(clk), .Q(
        matrix_mul_2D_4__2__6_), .QN(n2405) );
  DFF_X1 matrix_mul_2D_reg_4__2__7_ ( .D(n9054), .CK(clk), .Q(
        matrix_mul_2D_4__2__7_), .QN(n2404) );
  DFF_X1 matrix_mul_2D_reg_4__2__8_ ( .D(n9049), .CK(clk), .Q(
        matrix_mul_2D_4__2__8_), .QN(n2403) );
  DFF_X1 matrix_mul_2D_reg_4__2__9_ ( .D(n9044), .CK(clk), .Q(
        matrix_mul_2D_4__2__9_), .QN(n2402) );
  DFF_X1 matrix_mul_2D_reg_4__2__10_ ( .D(n9039), .CK(clk), .Q(
        matrix_mul_2D_4__2__10_), .QN(n2401) );
  DFF_X1 matrix_mul_2D_reg_4__2__11_ ( .D(n9034), .CK(clk), .Q(
        matrix_mul_2D_4__2__11_), .QN(n2400) );
  DFF_X1 matrix_mul_2D_reg_4__2__12_ ( .D(n9029), .CK(clk), .Q(
        matrix_mul_2D_4__2__12_), .QN(n2399) );
  DFF_X1 matrix_mul_2D_reg_4__2__13_ ( .D(n9024), .CK(clk), .Q(
        matrix_mul_2D_4__2__13_), .QN(n2398) );
  DFF_X1 matrix_mul_2D_reg_4__2__14_ ( .D(n9019), .CK(clk), .Q(
        matrix_mul_2D_4__2__14_), .QN(n2397) );
  DFF_X1 matrix_mul_2D_reg_4__2__15_ ( .D(n9018), .CK(clk), .Q(
        matrix_mul_2D_4__2__15_), .QN(n17628) );
  DFF_X1 matrix_mul_2D_reg_4__2__16_ ( .D(n9017), .CK(clk), .Q(
        matrix_mul_2D_4__2__16_), .QN(n17626) );
  DFF_X1 matrix_mul_2D_reg_4__2__17_ ( .D(n9016), .CK(clk), .Q(
        matrix_mul_2D_4__2__17_), .QN(n17624) );
  DFF_X1 matrix_mul_2D_reg_4__2__18_ ( .D(n9015), .CK(clk), .Q(
        matrix_mul_2D_4__2__18_), .QN(n17622) );
  DFF_X1 matrix_mul_2D_reg_4__2__19_ ( .D(n9014), .CK(clk), .Q(
        matrix_mul_2D_4__2__19_), .QN(n17620) );
  DFF_X1 matrix_mul_2D_reg_4__2__20_ ( .D(n9013), .CK(clk), .Q(
        matrix_mul_2D_4__2__20_), .QN(n17618) );
  DFF_X1 matrix_mul_2D_reg_4__3__0_ ( .D(n9009), .CK(clk), .Q(
        matrix_mul_2D_4__3__0_), .QN(n2426) );
  DFF_X1 matrix_mul_2D_reg_4__3__1_ ( .D(n9004), .CK(clk), .Q(
        matrix_mul_2D_4__3__1_), .QN(n2425) );
  DFF_X1 matrix_mul_2D_reg_4__3__2_ ( .D(n8999), .CK(clk), .Q(
        matrix_mul_2D_4__3__2_), .QN(n2424) );
  DFF_X1 matrix_mul_2D_reg_4__3__3_ ( .D(n8994), .CK(clk), .Q(
        matrix_mul_2D_4__3__3_), .QN(n2423) );
  DFF_X1 matrix_mul_2D_reg_4__3__4_ ( .D(n8989), .CK(clk), .Q(
        matrix_mul_2D_4__3__4_), .QN(n2422) );
  DFF_X1 matrix_mul_2D_reg_4__3__5_ ( .D(n8984), .CK(clk), .Q(
        matrix_mul_2D_4__3__5_), .QN(n2421) );
  DFF_X1 matrix_mul_2D_reg_4__3__6_ ( .D(n8979), .CK(clk), .Q(
        matrix_mul_2D_4__3__6_), .QN(n2420) );
  DFF_X1 matrix_mul_2D_reg_4__3__7_ ( .D(n8974), .CK(clk), .Q(
        matrix_mul_2D_4__3__7_), .QN(n2419) );
  DFF_X1 matrix_mul_2D_reg_4__3__8_ ( .D(n8969), .CK(clk), .Q(
        matrix_mul_2D_4__3__8_), .QN(n2418) );
  DFF_X1 matrix_mul_2D_reg_4__3__9_ ( .D(n8964), .CK(clk), .Q(
        matrix_mul_2D_4__3__9_), .QN(n2417) );
  DFF_X1 matrix_mul_2D_reg_4__3__10_ ( .D(n8959), .CK(clk), .Q(
        matrix_mul_2D_4__3__10_), .QN(n2416) );
  DFF_X1 matrix_mul_2D_reg_4__3__11_ ( .D(n8954), .CK(clk), .Q(
        matrix_mul_2D_4__3__11_), .QN(n2415) );
  DFF_X1 matrix_mul_2D_reg_4__3__12_ ( .D(n8949), .CK(clk), .Q(
        matrix_mul_2D_4__3__12_), .QN(n2414) );
  DFF_X1 matrix_mul_2D_reg_4__3__13_ ( .D(n8944), .CK(clk), .Q(
        matrix_mul_2D_4__3__13_), .QN(n2413) );
  DFF_X1 matrix_mul_2D_reg_4__3__14_ ( .D(n8939), .CK(clk), .Q(
        matrix_mul_2D_4__3__14_), .QN(n2412) );
  DFF_X1 matrix_mul_2D_reg_4__3__15_ ( .D(n8938), .CK(clk), .Q(
        matrix_mul_2D_4__3__15_), .QN(n17616) );
  DFF_X1 matrix_mul_2D_reg_4__3__16_ ( .D(n8937), .CK(clk), .Q(
        matrix_mul_2D_4__3__16_), .QN(n17614) );
  DFF_X1 matrix_mul_2D_reg_4__3__17_ ( .D(n8936), .CK(clk), .Q(
        matrix_mul_2D_4__3__17_), .QN(n17612) );
  DFF_X1 matrix_mul_2D_reg_4__3__18_ ( .D(n8935), .CK(clk), .Q(
        matrix_mul_2D_4__3__18_), .QN(n17610) );
  DFF_X1 matrix_mul_2D_reg_4__3__19_ ( .D(n8934), .CK(clk), .Q(
        matrix_mul_2D_4__3__19_), .QN(n17608) );
  DFF_X1 matrix_mul_2D_reg_4__3__20_ ( .D(n8933), .CK(clk), .Q(
        matrix_mul_2D_4__3__20_), .QN(n17606) );
  DFF_X1 matrix_mul_2D_reg_4__4__0_ ( .D(n8928), .CK(clk), .Q(
        matrix_mul_2D_4__4__0_), .QN(n2447) );
  DFF_X1 matrix_mul_2D_reg_4__4__1_ ( .D(n8924), .CK(clk), .Q(
        matrix_mul_2D_4__4__1_), .QN(n2446) );
  DFF_X1 matrix_mul_2D_reg_4__4__2_ ( .D(n8920), .CK(clk), .Q(
        matrix_mul_2D_4__4__2_), .QN(n2445) );
  DFF_X1 matrix_mul_2D_reg_4__4__3_ ( .D(n8916), .CK(clk), .Q(
        matrix_mul_2D_4__4__3_), .QN(n2444) );
  DFF_X1 matrix_mul_2D_reg_4__4__4_ ( .D(n8912), .CK(clk), .Q(
        matrix_mul_2D_4__4__4_), .QN(n2443) );
  DFF_X1 matrix_mul_2D_reg_4__4__5_ ( .D(n8908), .CK(clk), .Q(
        matrix_mul_2D_4__4__5_), .QN(n2442) );
  DFF_X1 matrix_mul_2D_reg_4__4__6_ ( .D(n8904), .CK(clk), .Q(
        matrix_mul_2D_4__4__6_), .QN(n2441) );
  DFF_X1 matrix_mul_2D_reg_4__4__7_ ( .D(n8900), .CK(clk), .Q(
        matrix_mul_2D_4__4__7_), .QN(n2440) );
  DFF_X1 matrix_mul_2D_reg_4__4__8_ ( .D(n8896), .CK(clk), .Q(
        matrix_mul_2D_4__4__8_), .QN(n2439) );
  DFF_X1 matrix_mul_2D_reg_4__4__9_ ( .D(n8892), .CK(clk), .Q(
        matrix_mul_2D_4__4__9_), .QN(n2438) );
  DFF_X1 matrix_mul_2D_reg_4__4__10_ ( .D(n8888), .CK(clk), .Q(
        matrix_mul_2D_4__4__10_), .QN(n2437) );
  DFF_X1 matrix_mul_2D_reg_4__4__11_ ( .D(n8884), .CK(clk), .Q(
        matrix_mul_2D_4__4__11_), .QN(n2436) );
  DFF_X1 matrix_mul_2D_reg_4__4__12_ ( .D(n8880), .CK(clk), .Q(
        matrix_mul_2D_4__4__12_), .QN(n2435) );
  DFF_X1 matrix_mul_2D_reg_4__4__13_ ( .D(n8876), .CK(clk), .Q(
        matrix_mul_2D_4__4__13_), .QN(n2434) );
  DFF_X1 matrix_mul_2D_reg_4__4__14_ ( .D(n8872), .CK(clk), .Q(
        matrix_mul_2D_4__4__14_), .QN(n2433) );
  DFF_X1 matrix_mul_2D_reg_4__4__15_ ( .D(n8871), .CK(clk), .Q(
        matrix_mul_2D_4__4__15_), .QN(n17604) );
  DFF_X1 matrix_mul_2D_reg_4__4__16_ ( .D(n8870), .CK(clk), .Q(
        matrix_mul_2D_4__4__16_), .QN(n17602) );
  DFF_X1 matrix_mul_2D_reg_4__4__17_ ( .D(n8869), .CK(clk), .Q(
        matrix_mul_2D_4__4__17_), .QN(n17600) );
  DFF_X1 matrix_mul_2D_reg_4__4__18_ ( .D(n8868), .CK(clk), .Q(
        matrix_mul_2D_4__4__18_), .QN(n17598) );
  DFF_X1 matrix_mul_2D_reg_4__4__19_ ( .D(n8867), .CK(clk), .Q(
        matrix_mul_2D_4__4__19_), .QN(n17596) );
  DFF_X1 matrix_mul_2D_reg_4__4__20_ ( .D(n8866), .CK(clk), .Q(
        matrix_mul_2D_4__4__20_), .QN(n17594) );
  DFF_X1 matrix_mul_2D_reg_4__5__0_ ( .D(n8861), .CK(clk), .Q(
        matrix_mul_2D_4__5__0_), .QN(n2462) );
  DFF_X1 matrix_mul_2D_reg_4__5__1_ ( .D(n8857), .CK(clk), .Q(
        matrix_mul_2D_4__5__1_), .QN(n2461) );
  DFF_X1 matrix_mul_2D_reg_4__5__2_ ( .D(n8853), .CK(clk), .Q(
        matrix_mul_2D_4__5__2_), .QN(n2460) );
  DFF_X1 matrix_mul_2D_reg_4__5__3_ ( .D(n8849), .CK(clk), .Q(
        matrix_mul_2D_4__5__3_), .QN(n2459) );
  DFF_X1 matrix_mul_2D_reg_4__5__4_ ( .D(n8845), .CK(clk), .Q(
        matrix_mul_2D_4__5__4_), .QN(n2458) );
  DFF_X1 matrix_mul_2D_reg_4__5__5_ ( .D(n8841), .CK(clk), .Q(
        matrix_mul_2D_4__5__5_), .QN(n2457) );
  DFF_X1 matrix_mul_2D_reg_4__5__6_ ( .D(n8837), .CK(clk), .Q(
        matrix_mul_2D_4__5__6_), .QN(n2456) );
  DFF_X1 matrix_mul_2D_reg_4__5__7_ ( .D(n8833), .CK(clk), .Q(
        matrix_mul_2D_4__5__7_), .QN(n2455) );
  DFF_X1 matrix_mul_2D_reg_4__5__8_ ( .D(n8829), .CK(clk), .Q(
        matrix_mul_2D_4__5__8_), .QN(n2454) );
  DFF_X1 matrix_mul_2D_reg_4__5__9_ ( .D(n8825), .CK(clk), .Q(
        matrix_mul_2D_4__5__9_), .QN(n2453) );
  DFF_X1 matrix_mul_2D_reg_4__5__10_ ( .D(n8821), .CK(clk), .Q(
        matrix_mul_2D_4__5__10_), .QN(n2452) );
  DFF_X1 matrix_mul_2D_reg_4__5__11_ ( .D(n8817), .CK(clk), .Q(
        matrix_mul_2D_4__5__11_), .QN(n2451) );
  DFF_X1 matrix_mul_2D_reg_4__5__12_ ( .D(n8813), .CK(clk), .Q(
        matrix_mul_2D_4__5__12_), .QN(n2450) );
  DFF_X1 matrix_mul_2D_reg_4__5__13_ ( .D(n8809), .CK(clk), .Q(
        matrix_mul_2D_4__5__13_), .QN(n2449) );
  DFF_X1 matrix_mul_2D_reg_4__5__14_ ( .D(n8805), .CK(clk), .Q(
        matrix_mul_2D_4__5__14_), .QN(n2448) );
  DFF_X1 matrix_mul_2D_reg_4__5__15_ ( .D(n8804), .CK(clk), .Q(
        matrix_mul_2D_4__5__15_), .QN(n17592) );
  DFF_X1 matrix_mul_2D_reg_4__5__16_ ( .D(n8803), .CK(clk), .Q(
        matrix_mul_2D_4__5__16_), .QN(n17590) );
  DFF_X1 matrix_mul_2D_reg_4__5__17_ ( .D(n8802), .CK(clk), .Q(
        matrix_mul_2D_4__5__17_), .QN(n17588) );
  DFF_X1 matrix_mul_2D_reg_4__5__18_ ( .D(n8801), .CK(clk), .Q(
        matrix_mul_2D_4__5__18_), .QN(n17586) );
  DFF_X1 matrix_mul_2D_reg_4__5__19_ ( .D(n8800), .CK(clk), .Q(
        matrix_mul_2D_4__5__19_), .QN(n17584) );
  DFF_X1 matrix_mul_2D_reg_4__5__20_ ( .D(n8799), .CK(clk), .Q(
        matrix_mul_2D_4__5__20_), .QN(n17582) );
  DFF_X1 matrix_mul_2D_reg_4__6__0_ ( .D(n8795), .CK(clk), .Q(
        matrix_mul_2D_4__6__0_), .QN(n2477) );
  DFF_X1 matrix_mul_2D_reg_4__6__1_ ( .D(n8790), .CK(clk), .Q(
        matrix_mul_2D_4__6__1_), .QN(n2476) );
  DFF_X1 matrix_mul_2D_reg_4__6__2_ ( .D(n8785), .CK(clk), .Q(
        matrix_mul_2D_4__6__2_), .QN(n2475) );
  DFF_X1 matrix_mul_2D_reg_4__6__3_ ( .D(n8780), .CK(clk), .Q(
        matrix_mul_2D_4__6__3_), .QN(n2474) );
  DFF_X1 matrix_mul_2D_reg_4__6__4_ ( .D(n8775), .CK(clk), .Q(
        matrix_mul_2D_4__6__4_), .QN(n2473) );
  DFF_X1 matrix_mul_2D_reg_4__6__5_ ( .D(n8770), .CK(clk), .Q(
        matrix_mul_2D_4__6__5_), .QN(n2472) );
  DFF_X1 matrix_mul_2D_reg_4__6__6_ ( .D(n8765), .CK(clk), .Q(
        matrix_mul_2D_4__6__6_), .QN(n2471) );
  DFF_X1 matrix_mul_2D_reg_4__6__7_ ( .D(n8760), .CK(clk), .Q(
        matrix_mul_2D_4__6__7_), .QN(n2470) );
  DFF_X1 matrix_mul_2D_reg_4__6__8_ ( .D(n8755), .CK(clk), .Q(
        matrix_mul_2D_4__6__8_), .QN(n2469) );
  DFF_X1 matrix_mul_2D_reg_4__6__9_ ( .D(n8750), .CK(clk), .Q(
        matrix_mul_2D_4__6__9_), .QN(n2468) );
  DFF_X1 matrix_mul_2D_reg_4__6__10_ ( .D(n8745), .CK(clk), .Q(
        matrix_mul_2D_4__6__10_), .QN(n2467) );
  DFF_X1 matrix_mul_2D_reg_4__6__11_ ( .D(n8740), .CK(clk), .Q(
        matrix_mul_2D_4__6__11_), .QN(n2466) );
  DFF_X1 matrix_mul_2D_reg_4__6__12_ ( .D(n8735), .CK(clk), .Q(
        matrix_mul_2D_4__6__12_), .QN(n2465) );
  DFF_X1 matrix_mul_2D_reg_4__6__13_ ( .D(n8730), .CK(clk), .Q(
        matrix_mul_2D_4__6__13_), .QN(n2464) );
  DFF_X1 matrix_mul_2D_reg_4__6__14_ ( .D(n8725), .CK(clk), .Q(
        matrix_mul_2D_4__6__14_), .QN(n2463) );
  DFF_X1 matrix_mul_2D_reg_4__6__15_ ( .D(n8724), .CK(clk), .Q(
        matrix_mul_2D_4__6__15_), .QN(n17580) );
  DFF_X1 matrix_mul_2D_reg_4__6__16_ ( .D(n8723), .CK(clk), .Q(
        matrix_mul_2D_4__6__16_), .QN(n17578) );
  DFF_X1 matrix_mul_2D_reg_4__6__17_ ( .D(n8722), .CK(clk), .Q(
        matrix_mul_2D_4__6__17_), .QN(n17576) );
  DFF_X1 matrix_mul_2D_reg_4__6__18_ ( .D(n8721), .CK(clk), .Q(
        matrix_mul_2D_4__6__18_), .QN(n17574) );
  DFF_X1 matrix_mul_2D_reg_4__6__19_ ( .D(n8720), .CK(clk), .Q(
        matrix_mul_2D_4__6__19_), .QN(n17572) );
  DFF_X1 matrix_mul_2D_reg_4__6__20_ ( .D(n8719), .CK(clk), .Q(
        matrix_mul_2D_4__6__20_), .QN(n17570) );
  DFF_X1 matrix_mul_2D_reg_4__7__0_ ( .D(n8715), .CK(clk), .Q(
        matrix_mul_2D_4__7__0_), .QN(n2492) );
  DFF_X1 matrix_mul_2D_reg_4__7__1_ ( .D(n8710), .CK(clk), .Q(
        matrix_mul_2D_4__7__1_), .QN(n2491) );
  DFF_X1 matrix_mul_2D_reg_4__7__2_ ( .D(n8705), .CK(clk), .Q(
        matrix_mul_2D_4__7__2_), .QN(n2490) );
  DFF_X1 matrix_mul_2D_reg_4__7__3_ ( .D(n8700), .CK(clk), .Q(
        matrix_mul_2D_4__7__3_), .QN(n2489) );
  DFF_X1 matrix_mul_2D_reg_4__7__4_ ( .D(n8695), .CK(clk), .Q(
        matrix_mul_2D_4__7__4_), .QN(n2488) );
  DFF_X1 matrix_mul_2D_reg_4__7__5_ ( .D(n8690), .CK(clk), .Q(
        matrix_mul_2D_4__7__5_), .QN(n2487) );
  DFF_X1 matrix_mul_2D_reg_4__7__6_ ( .D(n8685), .CK(clk), .Q(
        matrix_mul_2D_4__7__6_), .QN(n2486) );
  DFF_X1 matrix_mul_2D_reg_4__7__7_ ( .D(n8680), .CK(clk), .Q(
        matrix_mul_2D_4__7__7_), .QN(n2485) );
  DFF_X1 matrix_mul_2D_reg_4__7__8_ ( .D(n8675), .CK(clk), .Q(
        matrix_mul_2D_4__7__8_), .QN(n2484) );
  DFF_X1 matrix_mul_2D_reg_4__7__9_ ( .D(n8670), .CK(clk), .Q(
        matrix_mul_2D_4__7__9_), .QN(n2483) );
  DFF_X1 matrix_mul_2D_reg_4__7__10_ ( .D(n8665), .CK(clk), .Q(
        matrix_mul_2D_4__7__10_), .QN(n2482) );
  DFF_X1 matrix_mul_2D_reg_4__7__11_ ( .D(n8660), .CK(clk), .Q(
        matrix_mul_2D_4__7__11_), .QN(n2481) );
  DFF_X1 matrix_mul_2D_reg_4__7__12_ ( .D(n8655), .CK(clk), .Q(
        matrix_mul_2D_4__7__12_), .QN(n2480) );
  DFF_X1 matrix_mul_2D_reg_4__7__13_ ( .D(n8650), .CK(clk), .Q(
        matrix_mul_2D_4__7__13_), .QN(n2479) );
  DFF_X1 matrix_mul_2D_reg_4__7__14_ ( .D(n8645), .CK(clk), .Q(
        matrix_mul_2D_4__7__14_), .QN(n2478) );
  DFF_X1 matrix_mul_2D_reg_4__7__15_ ( .D(n8644), .CK(clk), .Q(
        matrix_mul_2D_4__7__15_), .QN(n17568) );
  DFF_X1 matrix_mul_2D_reg_4__7__16_ ( .D(n8643), .CK(clk), .Q(
        matrix_mul_2D_4__7__16_), .QN(n17566) );
  DFF_X1 matrix_mul_2D_reg_4__7__17_ ( .D(n8642), .CK(clk), .Q(
        matrix_mul_2D_4__7__17_), .QN(n17564) );
  DFF_X1 matrix_mul_2D_reg_4__7__18_ ( .D(n8641), .CK(clk), .Q(
        matrix_mul_2D_4__7__18_), .QN(n17562) );
  DFF_X1 matrix_mul_2D_reg_4__7__19_ ( .D(n8640), .CK(clk), .Q(
        matrix_mul_2D_4__7__19_), .QN(n17560) );
  DFF_X1 matrix_mul_2D_reg_4__7__20_ ( .D(n8639), .CK(clk), .Q(
        matrix_mul_2D_4__7__20_), .QN(n17558) );
  DFF_X1 matrix_mul_2D_reg_5__0__0_ ( .D(n8635), .CK(clk), .Q(
        matrix_mul_2D_5__0__0_), .QN(n2507) );
  DFF_X1 matrix_mul_2D_reg_5__0__1_ ( .D(n8630), .CK(clk), .Q(
        matrix_mul_2D_5__0__1_), .QN(n2506) );
  DFF_X1 matrix_mul_2D_reg_5__0__2_ ( .D(n8625), .CK(clk), .Q(
        matrix_mul_2D_5__0__2_), .QN(n2505) );
  DFF_X1 matrix_mul_2D_reg_5__0__3_ ( .D(n8620), .CK(clk), .Q(
        matrix_mul_2D_5__0__3_), .QN(n2504) );
  DFF_X1 matrix_mul_2D_reg_5__0__4_ ( .D(n8615), .CK(clk), .Q(
        matrix_mul_2D_5__0__4_), .QN(n2503) );
  DFF_X1 matrix_mul_2D_reg_5__0__5_ ( .D(n8610), .CK(clk), .Q(
        matrix_mul_2D_5__0__5_), .QN(n2502) );
  DFF_X1 matrix_mul_2D_reg_5__0__6_ ( .D(n8605), .CK(clk), .Q(
        matrix_mul_2D_5__0__6_), .QN(n2501) );
  DFF_X1 matrix_mul_2D_reg_5__0__7_ ( .D(n8600), .CK(clk), .Q(
        matrix_mul_2D_5__0__7_), .QN(n2500) );
  DFF_X1 matrix_mul_2D_reg_5__0__8_ ( .D(n8595), .CK(clk), .Q(
        matrix_mul_2D_5__0__8_), .QN(n2499) );
  DFF_X1 matrix_mul_2D_reg_5__0__9_ ( .D(n8590), .CK(clk), .Q(
        matrix_mul_2D_5__0__9_), .QN(n2498) );
  DFF_X1 matrix_mul_2D_reg_5__0__10_ ( .D(n8585), .CK(clk), .Q(
        matrix_mul_2D_5__0__10_), .QN(n2497) );
  DFF_X1 matrix_mul_2D_reg_5__0__11_ ( .D(n8580), .CK(clk), .Q(
        matrix_mul_2D_5__0__11_), .QN(n2496) );
  DFF_X1 matrix_mul_2D_reg_5__0__12_ ( .D(n8575), .CK(clk), .Q(
        matrix_mul_2D_5__0__12_), .QN(n2495) );
  DFF_X1 matrix_mul_2D_reg_5__0__13_ ( .D(n8570), .CK(clk), .Q(
        matrix_mul_2D_5__0__13_), .QN(n2494) );
  DFF_X1 matrix_mul_2D_reg_5__0__14_ ( .D(n8565), .CK(clk), .Q(
        matrix_mul_2D_5__0__14_), .QN(n2493) );
  DFF_X1 matrix_mul_2D_reg_5__0__15_ ( .D(n8564), .CK(clk), .Q(
        matrix_mul_2D_5__0__15_), .QN(n17556) );
  DFF_X1 matrix_mul_2D_reg_5__0__16_ ( .D(n8563), .CK(clk), .Q(
        matrix_mul_2D_5__0__16_), .QN(n17554) );
  DFF_X1 matrix_mul_2D_reg_5__0__17_ ( .D(n8562), .CK(clk), .Q(
        matrix_mul_2D_5__0__17_), .QN(n17552) );
  DFF_X1 matrix_mul_2D_reg_5__0__18_ ( .D(n8561), .CK(clk), .Q(
        matrix_mul_2D_5__0__18_), .QN(n17550) );
  DFF_X1 matrix_mul_2D_reg_5__0__19_ ( .D(n8560), .CK(clk), .Q(
        matrix_mul_2D_5__0__19_), .QN(n17548) );
  DFF_X1 matrix_mul_2D_reg_5__0__20_ ( .D(n8559), .CK(clk), .Q(
        matrix_mul_2D_5__0__20_), .QN(n17546) );
  DFF_X1 matrix_mul_2D_reg_5__1__0_ ( .D(n8555), .CK(clk), .Q(
        matrix_mul_2D_5__1__0_), .QN(n2522) );
  DFF_X1 matrix_mul_2D_reg_5__1__1_ ( .D(n8550), .CK(clk), .Q(
        matrix_mul_2D_5__1__1_), .QN(n2521) );
  DFF_X1 matrix_mul_2D_reg_5__1__2_ ( .D(n8545), .CK(clk), .Q(
        matrix_mul_2D_5__1__2_), .QN(n2520) );
  DFF_X1 matrix_mul_2D_reg_5__1__3_ ( .D(n8540), .CK(clk), .Q(
        matrix_mul_2D_5__1__3_), .QN(n2519) );
  DFF_X1 matrix_mul_2D_reg_5__1__4_ ( .D(n8535), .CK(clk), .Q(
        matrix_mul_2D_5__1__4_), .QN(n2518) );
  DFF_X1 matrix_mul_2D_reg_5__1__5_ ( .D(n8530), .CK(clk), .Q(
        matrix_mul_2D_5__1__5_), .QN(n2517) );
  DFF_X1 matrix_mul_2D_reg_5__1__6_ ( .D(n8525), .CK(clk), .Q(
        matrix_mul_2D_5__1__6_), .QN(n2516) );
  DFF_X1 matrix_mul_2D_reg_5__1__7_ ( .D(n8520), .CK(clk), .Q(
        matrix_mul_2D_5__1__7_), .QN(n2515) );
  DFF_X1 matrix_mul_2D_reg_5__1__8_ ( .D(n8515), .CK(clk), .Q(
        matrix_mul_2D_5__1__8_), .QN(n2514) );
  DFF_X1 matrix_mul_2D_reg_5__1__9_ ( .D(n8510), .CK(clk), .Q(
        matrix_mul_2D_5__1__9_), .QN(n2513) );
  DFF_X1 matrix_mul_2D_reg_5__1__10_ ( .D(n8505), .CK(clk), .Q(
        matrix_mul_2D_5__1__10_), .QN(n2512) );
  DFF_X1 matrix_mul_2D_reg_5__1__11_ ( .D(n8500), .CK(clk), .Q(
        matrix_mul_2D_5__1__11_), .QN(n2511) );
  DFF_X1 matrix_mul_2D_reg_5__1__12_ ( .D(n8495), .CK(clk), .Q(
        matrix_mul_2D_5__1__12_), .QN(n2510) );
  DFF_X1 matrix_mul_2D_reg_5__1__13_ ( .D(n8490), .CK(clk), .Q(
        matrix_mul_2D_5__1__13_), .QN(n2509) );
  DFF_X1 matrix_mul_2D_reg_5__1__14_ ( .D(n8485), .CK(clk), .Q(
        matrix_mul_2D_5__1__14_), .QN(n2508) );
  DFF_X1 matrix_mul_2D_reg_5__1__15_ ( .D(n8484), .CK(clk), .Q(
        matrix_mul_2D_5__1__15_), .QN(n17544) );
  DFF_X1 matrix_mul_2D_reg_5__1__16_ ( .D(n8483), .CK(clk), .Q(
        matrix_mul_2D_5__1__16_), .QN(n17542) );
  DFF_X1 matrix_mul_2D_reg_5__1__17_ ( .D(n8482), .CK(clk), .Q(
        matrix_mul_2D_5__1__17_), .QN(n17540) );
  DFF_X1 matrix_mul_2D_reg_5__1__18_ ( .D(n8481), .CK(clk), .Q(
        matrix_mul_2D_5__1__18_), .QN(n17538) );
  DFF_X1 matrix_mul_2D_reg_5__1__19_ ( .D(n8480), .CK(clk), .Q(
        matrix_mul_2D_5__1__19_), .QN(n17536) );
  DFF_X1 matrix_mul_2D_reg_5__1__20_ ( .D(n8479), .CK(clk), .Q(
        matrix_mul_2D_5__1__20_), .QN(n17534) );
  DFF_X1 matrix_mul_2D_reg_5__2__0_ ( .D(n8475), .CK(clk), .Q(
        matrix_mul_2D_5__2__0_), .QN(n2537) );
  DFF_X1 matrix_mul_2D_reg_5__2__1_ ( .D(n8470), .CK(clk), .Q(
        matrix_mul_2D_5__2__1_), .QN(n2536) );
  DFF_X1 matrix_mul_2D_reg_5__2__2_ ( .D(n8465), .CK(clk), .Q(
        matrix_mul_2D_5__2__2_), .QN(n2535) );
  DFF_X1 matrix_mul_2D_reg_5__2__3_ ( .D(n8460), .CK(clk), .Q(
        matrix_mul_2D_5__2__3_), .QN(n2534) );
  DFF_X1 matrix_mul_2D_reg_5__2__4_ ( .D(n8455), .CK(clk), .Q(
        matrix_mul_2D_5__2__4_), .QN(n2533) );
  DFF_X1 matrix_mul_2D_reg_5__2__5_ ( .D(n8450), .CK(clk), .Q(
        matrix_mul_2D_5__2__5_), .QN(n2532) );
  DFF_X1 matrix_mul_2D_reg_5__2__6_ ( .D(n8445), .CK(clk), .Q(
        matrix_mul_2D_5__2__6_), .QN(n2531) );
  DFF_X1 matrix_mul_2D_reg_5__2__7_ ( .D(n8440), .CK(clk), .Q(
        matrix_mul_2D_5__2__7_), .QN(n2530) );
  DFF_X1 matrix_mul_2D_reg_5__2__8_ ( .D(n8435), .CK(clk), .Q(
        matrix_mul_2D_5__2__8_), .QN(n2529) );
  DFF_X1 matrix_mul_2D_reg_5__2__9_ ( .D(n8430), .CK(clk), .Q(
        matrix_mul_2D_5__2__9_), .QN(n2528) );
  DFF_X1 matrix_mul_2D_reg_5__2__10_ ( .D(n8425), .CK(clk), .Q(
        matrix_mul_2D_5__2__10_), .QN(n2527) );
  DFF_X1 matrix_mul_2D_reg_5__2__11_ ( .D(n8420), .CK(clk), .Q(
        matrix_mul_2D_5__2__11_), .QN(n2526) );
  DFF_X1 matrix_mul_2D_reg_5__2__12_ ( .D(n8415), .CK(clk), .Q(
        matrix_mul_2D_5__2__12_), .QN(n2525) );
  DFF_X1 matrix_mul_2D_reg_5__2__13_ ( .D(n8410), .CK(clk), .Q(
        matrix_mul_2D_5__2__13_), .QN(n2524) );
  DFF_X1 matrix_mul_2D_reg_5__2__14_ ( .D(n8405), .CK(clk), .Q(
        matrix_mul_2D_5__2__14_), .QN(n2523) );
  DFF_X1 matrix_mul_2D_reg_5__2__15_ ( .D(n8404), .CK(clk), .Q(
        matrix_mul_2D_5__2__15_), .QN(n17532) );
  DFF_X1 matrix_mul_2D_reg_5__2__16_ ( .D(n8403), .CK(clk), .Q(
        matrix_mul_2D_5__2__16_), .QN(n17530) );
  DFF_X1 matrix_mul_2D_reg_5__2__17_ ( .D(n8402), .CK(clk), .Q(
        matrix_mul_2D_5__2__17_), .QN(n17528) );
  DFF_X1 matrix_mul_2D_reg_5__2__18_ ( .D(n8401), .CK(clk), .Q(
        matrix_mul_2D_5__2__18_), .QN(n17526) );
  DFF_X1 matrix_mul_2D_reg_5__2__19_ ( .D(n8400), .CK(clk), .Q(
        matrix_mul_2D_5__2__19_), .QN(n17524) );
  DFF_X1 matrix_mul_2D_reg_5__2__20_ ( .D(n8399), .CK(clk), .Q(
        matrix_mul_2D_5__2__20_), .QN(n17522) );
  DFF_X1 matrix_mul_2D_reg_5__3__0_ ( .D(n8395), .CK(clk), .Q(
        matrix_mul_2D_5__3__0_), .QN(n2552) );
  DFF_X1 matrix_mul_2D_reg_5__3__1_ ( .D(n8390), .CK(clk), .Q(
        matrix_mul_2D_5__3__1_), .QN(n2551) );
  DFF_X1 matrix_mul_2D_reg_5__3__2_ ( .D(n8385), .CK(clk), .Q(
        matrix_mul_2D_5__3__2_), .QN(n2550) );
  DFF_X1 matrix_mul_2D_reg_5__3__3_ ( .D(n8380), .CK(clk), .Q(
        matrix_mul_2D_5__3__3_), .QN(n2549) );
  DFF_X1 matrix_mul_2D_reg_5__3__4_ ( .D(n8375), .CK(clk), .Q(
        matrix_mul_2D_5__3__4_), .QN(n2548) );
  DFF_X1 matrix_mul_2D_reg_5__3__5_ ( .D(n8370), .CK(clk), .Q(
        matrix_mul_2D_5__3__5_), .QN(n2547) );
  DFF_X1 matrix_mul_2D_reg_5__3__6_ ( .D(n8365), .CK(clk), .Q(
        matrix_mul_2D_5__3__6_), .QN(n2546) );
  DFF_X1 matrix_mul_2D_reg_5__3__7_ ( .D(n8360), .CK(clk), .Q(
        matrix_mul_2D_5__3__7_), .QN(n2545) );
  DFF_X1 matrix_mul_2D_reg_5__3__8_ ( .D(n8355), .CK(clk), .Q(
        matrix_mul_2D_5__3__8_), .QN(n2544) );
  DFF_X1 matrix_mul_2D_reg_5__3__9_ ( .D(n8350), .CK(clk), .Q(
        matrix_mul_2D_5__3__9_), .QN(n2543) );
  DFF_X1 matrix_mul_2D_reg_5__3__10_ ( .D(n8345), .CK(clk), .Q(
        matrix_mul_2D_5__3__10_), .QN(n2542) );
  DFF_X1 matrix_mul_2D_reg_5__3__11_ ( .D(n8340), .CK(clk), .Q(
        matrix_mul_2D_5__3__11_), .QN(n2541) );
  DFF_X1 matrix_mul_2D_reg_5__3__12_ ( .D(n8335), .CK(clk), .Q(
        matrix_mul_2D_5__3__12_), .QN(n2540) );
  DFF_X1 matrix_mul_2D_reg_5__3__13_ ( .D(n8330), .CK(clk), .Q(
        matrix_mul_2D_5__3__13_), .QN(n2539) );
  DFF_X1 matrix_mul_2D_reg_5__3__14_ ( .D(n8325), .CK(clk), .Q(
        matrix_mul_2D_5__3__14_), .QN(n2538) );
  DFF_X1 matrix_mul_2D_reg_5__3__15_ ( .D(n8324), .CK(clk), .Q(
        matrix_mul_2D_5__3__15_), .QN(n17520) );
  DFF_X1 matrix_mul_2D_reg_5__3__16_ ( .D(n8323), .CK(clk), .Q(
        matrix_mul_2D_5__3__16_), .QN(n17518) );
  DFF_X1 matrix_mul_2D_reg_5__3__17_ ( .D(n8322), .CK(clk), .Q(
        matrix_mul_2D_5__3__17_), .QN(n17516) );
  DFF_X1 matrix_mul_2D_reg_5__3__18_ ( .D(n8321), .CK(clk), .Q(
        matrix_mul_2D_5__3__18_), .QN(n17514) );
  DFF_X1 matrix_mul_2D_reg_5__3__19_ ( .D(n8320), .CK(clk), .Q(
        matrix_mul_2D_5__3__19_), .QN(n17512) );
  DFF_X1 matrix_mul_2D_reg_5__3__20_ ( .D(n8319), .CK(clk), .Q(
        matrix_mul_2D_5__3__20_), .QN(n17510) );
  DFF_X1 matrix_mul_2D_reg_5__4__0_ ( .D(n8314), .CK(clk), .Q(
        matrix_mul_2D_5__4__0_), .QN(n257300) );
  DFF_X1 matrix_mul_2D_reg_5__4__1_ ( .D(n8310), .CK(clk), .Q(
        matrix_mul_2D_5__4__1_), .QN(n257200) );
  DFF_X1 matrix_mul_2D_reg_5__4__2_ ( .D(n8306), .CK(clk), .Q(
        matrix_mul_2D_5__4__2_), .QN(n257100) );
  DFF_X1 matrix_mul_2D_reg_5__4__3_ ( .D(n8302), .CK(clk), .Q(
        matrix_mul_2D_5__4__3_), .QN(n257000) );
  DFF_X1 matrix_mul_2D_reg_5__4__4_ ( .D(n8298), .CK(clk), .Q(
        matrix_mul_2D_5__4__4_), .QN(n256900) );
  DFF_X1 matrix_mul_2D_reg_5__4__5_ ( .D(n8294), .CK(clk), .Q(
        matrix_mul_2D_5__4__5_), .QN(n256800) );
  DFF_X1 matrix_mul_2D_reg_5__4__6_ ( .D(n8290), .CK(clk), .Q(
        matrix_mul_2D_5__4__6_), .QN(n256700) );
  DFF_X1 matrix_mul_2D_reg_5__4__7_ ( .D(n8286), .CK(clk), .Q(
        matrix_mul_2D_5__4__7_), .QN(n256600) );
  DFF_X1 matrix_mul_2D_reg_5__4__8_ ( .D(n8282), .CK(clk), .Q(
        matrix_mul_2D_5__4__8_), .QN(n256500) );
  DFF_X1 matrix_mul_2D_reg_5__4__9_ ( .D(n8278), .CK(clk), .Q(
        matrix_mul_2D_5__4__9_), .QN(n256400) );
  DFF_X1 matrix_mul_2D_reg_5__4__10_ ( .D(n8274), .CK(clk), .Q(
        matrix_mul_2D_5__4__10_), .QN(n256300) );
  DFF_X1 matrix_mul_2D_reg_5__4__11_ ( .D(n8270), .CK(clk), .Q(
        matrix_mul_2D_5__4__11_), .QN(n256200) );
  DFF_X1 matrix_mul_2D_reg_5__4__12_ ( .D(n8266), .CK(clk), .Q(
        matrix_mul_2D_5__4__12_), .QN(n256100) );
  DFF_X1 matrix_mul_2D_reg_5__4__13_ ( .D(n8262), .CK(clk), .Q(
        matrix_mul_2D_5__4__13_), .QN(n256000) );
  DFF_X1 matrix_mul_2D_reg_5__4__14_ ( .D(n8258), .CK(clk), .Q(
        matrix_mul_2D_5__4__14_), .QN(n255900) );
  DFF_X1 matrix_mul_2D_reg_5__4__15_ ( .D(n8257), .CK(clk), .Q(
        matrix_mul_2D_5__4__15_), .QN(n17508) );
  DFF_X1 matrix_mul_2D_reg_5__4__16_ ( .D(n8256), .CK(clk), .Q(
        matrix_mul_2D_5__4__16_), .QN(n17506) );
  DFF_X1 matrix_mul_2D_reg_5__4__17_ ( .D(n8255), .CK(clk), .Q(
        matrix_mul_2D_5__4__17_), .QN(n17504) );
  DFF_X1 matrix_mul_2D_reg_5__4__18_ ( .D(n8254), .CK(clk), .Q(
        matrix_mul_2D_5__4__18_), .QN(n17502) );
  DFF_X1 matrix_mul_2D_reg_5__4__19_ ( .D(n8253), .CK(clk), .Q(
        matrix_mul_2D_5__4__19_), .QN(n17500) );
  DFF_X1 matrix_mul_2D_reg_5__4__20_ ( .D(n8252), .CK(clk), .Q(
        matrix_mul_2D_5__4__20_), .QN(n17498) );
  DFF_X1 matrix_mul_2D_reg_5__5__0_ ( .D(n8247), .CK(clk), .Q(
        matrix_mul_2D_5__5__0_), .QN(n2588) );
  DFF_X1 matrix_mul_2D_reg_5__5__1_ ( .D(n8243), .CK(clk), .Q(
        matrix_mul_2D_5__5__1_), .QN(n2587) );
  DFF_X1 matrix_mul_2D_reg_5__5__2_ ( .D(n8239), .CK(clk), .Q(
        matrix_mul_2D_5__5__2_), .QN(n2586) );
  DFF_X1 matrix_mul_2D_reg_5__5__3_ ( .D(n8235), .CK(clk), .Q(
        matrix_mul_2D_5__5__3_), .QN(n2585) );
  DFF_X1 matrix_mul_2D_reg_5__5__4_ ( .D(n8231), .CK(clk), .Q(
        matrix_mul_2D_5__5__4_), .QN(n2584) );
  DFF_X1 matrix_mul_2D_reg_5__5__5_ ( .D(n8227), .CK(clk), .Q(
        matrix_mul_2D_5__5__5_), .QN(n2583) );
  DFF_X1 matrix_mul_2D_reg_5__5__6_ ( .D(n8223), .CK(clk), .Q(
        matrix_mul_2D_5__5__6_), .QN(n2582) );
  DFF_X1 matrix_mul_2D_reg_5__5__7_ ( .D(n8219), .CK(clk), .Q(
        matrix_mul_2D_5__5__7_), .QN(n2581) );
  DFF_X1 matrix_mul_2D_reg_5__5__8_ ( .D(n8215), .CK(clk), .Q(
        matrix_mul_2D_5__5__8_), .QN(n2580) );
  DFF_X1 matrix_mul_2D_reg_5__5__9_ ( .D(n8211), .CK(clk), .Q(
        matrix_mul_2D_5__5__9_), .QN(n2579) );
  DFF_X1 matrix_mul_2D_reg_5__5__10_ ( .D(n8207), .CK(clk), .Q(
        matrix_mul_2D_5__5__10_), .QN(n2578) );
  DFF_X1 matrix_mul_2D_reg_5__5__11_ ( .D(n8203), .CK(clk), .Q(
        matrix_mul_2D_5__5__11_), .QN(n2577) );
  DFF_X1 matrix_mul_2D_reg_5__5__12_ ( .D(n8199), .CK(clk), .Q(
        matrix_mul_2D_5__5__12_), .QN(n2576) );
  DFF_X1 matrix_mul_2D_reg_5__5__13_ ( .D(n8195), .CK(clk), .Q(
        matrix_mul_2D_5__5__13_), .QN(n2575) );
  DFF_X1 matrix_mul_2D_reg_5__5__14_ ( .D(n8191), .CK(clk), .Q(
        matrix_mul_2D_5__5__14_), .QN(n257400) );
  DFF_X1 matrix_mul_2D_reg_5__5__15_ ( .D(n8190), .CK(clk), .Q(
        matrix_mul_2D_5__5__15_), .QN(n17496) );
  DFF_X1 matrix_mul_2D_reg_5__5__16_ ( .D(n8189), .CK(clk), .Q(
        matrix_mul_2D_5__5__16_), .QN(n17494) );
  DFF_X1 matrix_mul_2D_reg_5__5__17_ ( .D(n8188), .CK(clk), .Q(
        matrix_mul_2D_5__5__17_), .QN(n17492) );
  DFF_X1 matrix_mul_2D_reg_5__5__18_ ( .D(n8187), .CK(clk), .Q(
        matrix_mul_2D_5__5__18_), .QN(n17490) );
  DFF_X1 matrix_mul_2D_reg_5__5__19_ ( .D(n8186), .CK(clk), .Q(
        matrix_mul_2D_5__5__19_), .QN(n17488) );
  DFF_X1 matrix_mul_2D_reg_5__5__20_ ( .D(n8185), .CK(clk), .Q(
        matrix_mul_2D_5__5__20_), .QN(n17486) );
  DFF_X1 matrix_mul_2D_reg_5__6__0_ ( .D(n8181), .CK(clk), .Q(
        matrix_mul_2D_5__6__0_), .QN(n260300) );
  DFF_X1 matrix_mul_2D_reg_5__6__1_ ( .D(n8176), .CK(clk), .Q(
        matrix_mul_2D_5__6__1_), .QN(n260200) );
  DFF_X1 matrix_mul_2D_reg_5__6__2_ ( .D(n8171), .CK(clk), .Q(
        matrix_mul_2D_5__6__2_), .QN(n260100) );
  DFF_X1 matrix_mul_2D_reg_5__6__3_ ( .D(n8166), .CK(clk), .Q(
        matrix_mul_2D_5__6__3_), .QN(n260000) );
  DFF_X1 matrix_mul_2D_reg_5__6__4_ ( .D(n8161), .CK(clk), .Q(
        matrix_mul_2D_5__6__4_), .QN(n259900) );
  DFF_X1 matrix_mul_2D_reg_5__6__5_ ( .D(n8156), .CK(clk), .Q(
        matrix_mul_2D_5__6__5_), .QN(n259800) );
  DFF_X1 matrix_mul_2D_reg_5__6__6_ ( .D(n8151), .CK(clk), .Q(
        matrix_mul_2D_5__6__6_), .QN(n259700) );
  DFF_X1 matrix_mul_2D_reg_5__6__7_ ( .D(n8146), .CK(clk), .Q(
        matrix_mul_2D_5__6__7_), .QN(n259600) );
  DFF_X1 matrix_mul_2D_reg_5__6__8_ ( .D(n8141), .CK(clk), .Q(
        matrix_mul_2D_5__6__8_), .QN(n259500) );
  DFF_X1 matrix_mul_2D_reg_5__6__9_ ( .D(n8136), .CK(clk), .Q(
        matrix_mul_2D_5__6__9_), .QN(n259400) );
  DFF_X1 matrix_mul_2D_reg_5__6__10_ ( .D(n8131), .CK(clk), .Q(
        matrix_mul_2D_5__6__10_), .QN(n259300) );
  DFF_X1 matrix_mul_2D_reg_5__6__11_ ( .D(n8126), .CK(clk), .Q(
        matrix_mul_2D_5__6__11_), .QN(n259200) );
  DFF_X1 matrix_mul_2D_reg_5__6__12_ ( .D(n8121), .CK(clk), .Q(
        matrix_mul_2D_5__6__12_), .QN(n2591) );
  DFF_X1 matrix_mul_2D_reg_5__6__13_ ( .D(n8116), .CK(clk), .Q(
        matrix_mul_2D_5__6__13_), .QN(n2590) );
  DFF_X1 matrix_mul_2D_reg_5__6__14_ ( .D(n8111), .CK(clk), .Q(
        matrix_mul_2D_5__6__14_), .QN(n2589) );
  DFF_X1 matrix_mul_2D_reg_5__6__15_ ( .D(n8110), .CK(clk), .Q(
        matrix_mul_2D_5__6__15_), .QN(n17484) );
  DFF_X1 matrix_mul_2D_reg_5__6__16_ ( .D(n8109), .CK(clk), .Q(
        matrix_mul_2D_5__6__16_), .QN(n17482) );
  DFF_X1 matrix_mul_2D_reg_5__6__17_ ( .D(n8108), .CK(clk), .Q(
        matrix_mul_2D_5__6__17_), .QN(n17480) );
  DFF_X1 matrix_mul_2D_reg_5__6__18_ ( .D(n8107), .CK(clk), .Q(
        matrix_mul_2D_5__6__18_), .QN(n17478) );
  DFF_X1 matrix_mul_2D_reg_5__6__19_ ( .D(n8106), .CK(clk), .Q(
        matrix_mul_2D_5__6__19_), .QN(n17476) );
  DFF_X1 matrix_mul_2D_reg_5__6__20_ ( .D(n8105), .CK(clk), .Q(
        matrix_mul_2D_5__6__20_), .QN(n17474) );
  DFF_X1 matrix_mul_2D_reg_5__7__0_ ( .D(n8101), .CK(clk), .Q(
        matrix_mul_2D_5__7__0_), .QN(n2618) );
  DFF_X1 matrix_mul_2D_reg_5__7__1_ ( .D(n8096), .CK(clk), .Q(
        matrix_mul_2D_5__7__1_), .QN(n2617) );
  DFF_X1 matrix_mul_2D_reg_5__7__2_ ( .D(n8091), .CK(clk), .Q(
        matrix_mul_2D_5__7__2_), .QN(n2616) );
  DFF_X1 matrix_mul_2D_reg_5__7__3_ ( .D(n8086), .CK(clk), .Q(
        matrix_mul_2D_5__7__3_), .QN(n2615) );
  DFF_X1 matrix_mul_2D_reg_5__7__4_ ( .D(n8081), .CK(clk), .Q(
        matrix_mul_2D_5__7__4_), .QN(n2614) );
  DFF_X1 matrix_mul_2D_reg_5__7__5_ ( .D(n8076), .CK(clk), .Q(
        matrix_mul_2D_5__7__5_), .QN(n2613) );
  DFF_X1 matrix_mul_2D_reg_5__7__6_ ( .D(n8071), .CK(clk), .Q(
        matrix_mul_2D_5__7__6_), .QN(n261200) );
  DFF_X1 matrix_mul_2D_reg_5__7__7_ ( .D(n8066), .CK(clk), .Q(
        matrix_mul_2D_5__7__7_), .QN(n261100) );
  DFF_X1 matrix_mul_2D_reg_5__7__8_ ( .D(n8061), .CK(clk), .Q(
        matrix_mul_2D_5__7__8_), .QN(n261000) );
  DFF_X1 matrix_mul_2D_reg_5__7__9_ ( .D(n8056), .CK(clk), .Q(
        matrix_mul_2D_5__7__9_), .QN(n260900) );
  DFF_X1 matrix_mul_2D_reg_5__7__10_ ( .D(n8051), .CK(clk), .Q(
        matrix_mul_2D_5__7__10_), .QN(n260800) );
  DFF_X1 matrix_mul_2D_reg_5__7__11_ ( .D(n8046), .CK(clk), .Q(
        matrix_mul_2D_5__7__11_), .QN(n260700) );
  DFF_X1 matrix_mul_2D_reg_5__7__12_ ( .D(n8041), .CK(clk), .Q(
        matrix_mul_2D_5__7__12_), .QN(n260600) );
  DFF_X1 matrix_mul_2D_reg_5__7__13_ ( .D(n8036), .CK(clk), .Q(
        matrix_mul_2D_5__7__13_), .QN(n260500) );
  DFF_X1 matrix_mul_2D_reg_5__7__14_ ( .D(n8031), .CK(clk), .Q(
        matrix_mul_2D_5__7__14_), .QN(n260400) );
  DFF_X1 matrix_mul_2D_reg_5__7__15_ ( .D(n8030), .CK(clk), .Q(
        matrix_mul_2D_5__7__15_), .QN(n17472) );
  DFF_X1 matrix_mul_2D_reg_5__7__16_ ( .D(n8029), .CK(clk), .Q(
        matrix_mul_2D_5__7__16_), .QN(n17470) );
  DFF_X1 matrix_mul_2D_reg_5__7__17_ ( .D(n8028), .CK(clk), .Q(
        matrix_mul_2D_5__7__17_), .QN(n17468) );
  DFF_X1 matrix_mul_2D_reg_5__7__18_ ( .D(n8027), .CK(clk), .Q(
        matrix_mul_2D_5__7__18_), .QN(n17466) );
  DFF_X1 matrix_mul_2D_reg_5__7__19_ ( .D(n8026), .CK(clk), .Q(
        matrix_mul_2D_5__7__19_), .QN(n17464) );
  DFF_X1 matrix_mul_2D_reg_5__7__20_ ( .D(n8025), .CK(clk), .Q(
        matrix_mul_2D_5__7__20_), .QN(n17462) );
  DFF_X1 matrix_mul_2D_reg_6__0__0_ ( .D(n8021), .CK(clk), .Q(
        matrix_mul_2D_6__0__0_), .QN(n2633) );
  DFF_X1 matrix_mul_2D_reg_6__0__1_ ( .D(n8016), .CK(clk), .Q(
        matrix_mul_2D_6__0__1_), .QN(n2632) );
  DFF_X1 matrix_mul_2D_reg_6__0__2_ ( .D(n8011), .CK(clk), .Q(
        matrix_mul_2D_6__0__2_), .QN(n2631) );
  DFF_X1 matrix_mul_2D_reg_6__0__3_ ( .D(n8006), .CK(clk), .Q(
        matrix_mul_2D_6__0__3_), .QN(n2630) );
  DFF_X1 matrix_mul_2D_reg_6__0__4_ ( .D(n8001), .CK(clk), .Q(
        matrix_mul_2D_6__0__4_), .QN(n2629) );
  DFF_X1 matrix_mul_2D_reg_6__0__5_ ( .D(n79960), .CK(clk), .Q(
        matrix_mul_2D_6__0__5_), .QN(n2628) );
  DFF_X1 matrix_mul_2D_reg_6__0__6_ ( .D(n79910), .CK(clk), .Q(
        matrix_mul_2D_6__0__6_), .QN(n2627) );
  DFF_X1 matrix_mul_2D_reg_6__0__7_ ( .D(n79860), .CK(clk), .Q(
        matrix_mul_2D_6__0__7_), .QN(n2626) );
  DFF_X1 matrix_mul_2D_reg_6__0__8_ ( .D(n79810), .CK(clk), .Q(
        matrix_mul_2D_6__0__8_), .QN(n2625) );
  DFF_X1 matrix_mul_2D_reg_6__0__9_ ( .D(n7976), .CK(clk), .Q(
        matrix_mul_2D_6__0__9_), .QN(n2624) );
  DFF_X1 matrix_mul_2D_reg_6__0__10_ ( .D(n7971), .CK(clk), .Q(
        matrix_mul_2D_6__0__10_), .QN(n2623) );
  DFF_X1 matrix_mul_2D_reg_6__0__11_ ( .D(n7966), .CK(clk), .Q(
        matrix_mul_2D_6__0__11_), .QN(n2622) );
  DFF_X1 matrix_mul_2D_reg_6__0__12_ ( .D(n79610), .CK(clk), .Q(
        matrix_mul_2D_6__0__12_), .QN(n2621) );
  DFF_X1 matrix_mul_2D_reg_6__0__13_ ( .D(n79560), .CK(clk), .Q(
        matrix_mul_2D_6__0__13_), .QN(n2620) );
  DFF_X1 matrix_mul_2D_reg_6__0__14_ ( .D(n79510), .CK(clk), .Q(
        matrix_mul_2D_6__0__14_), .QN(n2619) );
  DFF_X1 matrix_mul_2D_reg_6__0__15_ ( .D(n79500), .CK(clk), .Q(
        matrix_mul_2D_6__0__15_), .QN(n17460) );
  DFF_X1 matrix_mul_2D_reg_6__0__16_ ( .D(n79490), .CK(clk), .Q(
        matrix_mul_2D_6__0__16_), .QN(n17458) );
  DFF_X1 matrix_mul_2D_reg_6__0__17_ ( .D(n79480), .CK(clk), .Q(
        matrix_mul_2D_6__0__17_), .QN(n17456) );
  DFF_X1 matrix_mul_2D_reg_6__0__18_ ( .D(n79470), .CK(clk), .Q(
        matrix_mul_2D_6__0__18_), .QN(n17454) );
  DFF_X1 matrix_mul_2D_reg_6__0__19_ ( .D(n79460), .CK(clk), .Q(
        matrix_mul_2D_6__0__19_), .QN(n17452) );
  DFF_X1 matrix_mul_2D_reg_6__0__20_ ( .D(n7945), .CK(clk), .Q(
        matrix_mul_2D_6__0__20_), .QN(n17450) );
  DFF_X1 matrix_mul_2D_reg_6__1__0_ ( .D(n7941), .CK(clk), .Q(
        matrix_mul_2D_6__1__0_), .QN(n264800) );
  DFF_X1 matrix_mul_2D_reg_6__1__1_ ( .D(n7936), .CK(clk), .Q(
        matrix_mul_2D_6__1__1_), .QN(n264700) );
  DFF_X1 matrix_mul_2D_reg_6__1__2_ ( .D(n7931), .CK(clk), .Q(
        matrix_mul_2D_6__1__2_), .QN(n264600) );
  DFF_X1 matrix_mul_2D_reg_6__1__3_ ( .D(n7926), .CK(clk), .Q(
        matrix_mul_2D_6__1__3_), .QN(n264500) );
  DFF_X1 matrix_mul_2D_reg_6__1__4_ ( .D(n7921), .CK(clk), .Q(
        matrix_mul_2D_6__1__4_), .QN(n264400) );
  DFF_X1 matrix_mul_2D_reg_6__1__5_ ( .D(n79160), .CK(clk), .Q(
        matrix_mul_2D_6__1__5_), .QN(n264300) );
  DFF_X1 matrix_mul_2D_reg_6__1__6_ ( .D(n79110), .CK(clk), .Q(
        matrix_mul_2D_6__1__6_), .QN(n264200) );
  DFF_X1 matrix_mul_2D_reg_6__1__7_ ( .D(n79060), .CK(clk), .Q(
        matrix_mul_2D_6__1__7_), .QN(n264100) );
  DFF_X1 matrix_mul_2D_reg_6__1__8_ ( .D(n79010), .CK(clk), .Q(
        matrix_mul_2D_6__1__8_), .QN(n2640) );
  DFF_X1 matrix_mul_2D_reg_6__1__9_ ( .D(n7896), .CK(clk), .Q(
        matrix_mul_2D_6__1__9_), .QN(n2639) );
  DFF_X1 matrix_mul_2D_reg_6__1__10_ ( .D(n7891), .CK(clk), .Q(
        matrix_mul_2D_6__1__10_), .QN(n2638) );
  DFF_X1 matrix_mul_2D_reg_6__1__11_ ( .D(n7886), .CK(clk), .Q(
        matrix_mul_2D_6__1__11_), .QN(n263700) );
  DFF_X1 matrix_mul_2D_reg_6__1__12_ ( .D(n7881), .CK(clk), .Q(
        matrix_mul_2D_6__1__12_), .QN(n2636) );
  DFF_X1 matrix_mul_2D_reg_6__1__13_ ( .D(n78760), .CK(clk), .Q(
        matrix_mul_2D_6__1__13_), .QN(n2635) );
  DFF_X1 matrix_mul_2D_reg_6__1__14_ ( .D(n78710), .CK(clk), .Q(
        matrix_mul_2D_6__1__14_), .QN(n2634) );
  DFF_X1 matrix_mul_2D_reg_6__1__15_ ( .D(n78700), .CK(clk), .Q(
        matrix_mul_2D_6__1__15_), .QN(n17448) );
  DFF_X1 matrix_mul_2D_reg_6__1__16_ ( .D(n78690), .CK(clk), .Q(
        matrix_mul_2D_6__1__16_), .QN(n17446) );
  DFF_X1 matrix_mul_2D_reg_6__1__17_ ( .D(n78680), .CK(clk), .Q(
        matrix_mul_2D_6__1__17_), .QN(n17444) );
  DFF_X1 matrix_mul_2D_reg_6__1__18_ ( .D(n78670), .CK(clk), .Q(
        matrix_mul_2D_6__1__18_), .QN(n17442) );
  DFF_X1 matrix_mul_2D_reg_6__1__19_ ( .D(n78660), .CK(clk), .Q(
        matrix_mul_2D_6__1__19_), .QN(n17440) );
  DFF_X1 matrix_mul_2D_reg_6__1__20_ ( .D(n78650), .CK(clk), .Q(
        matrix_mul_2D_6__1__20_), .QN(n17438) );
  DFF_X1 matrix_mul_2D_reg_6__2__0_ ( .D(n7860), .CK(clk), .Q(
        matrix_mul_2D_6__2__0_), .QN(n2669) );
  DFF_X1 matrix_mul_2D_reg_6__2__1_ ( .D(n7856), .CK(clk), .Q(
        matrix_mul_2D_6__2__1_), .QN(n2668) );
  DFF_X1 matrix_mul_2D_reg_6__2__2_ ( .D(n7852), .CK(clk), .Q(
        matrix_mul_2D_6__2__2_), .QN(n2667) );
  DFF_X1 matrix_mul_2D_reg_6__2__3_ ( .D(n7848), .CK(clk), .Q(
        matrix_mul_2D_6__2__3_), .QN(n2666) );
  DFF_X1 matrix_mul_2D_reg_6__2__4_ ( .D(n7844), .CK(clk), .Q(
        matrix_mul_2D_6__2__4_), .QN(n2665) );
  DFF_X1 matrix_mul_2D_reg_6__2__5_ ( .D(n7840), .CK(clk), .Q(
        matrix_mul_2D_6__2__5_), .QN(n2664) );
  DFF_X1 matrix_mul_2D_reg_6__2__6_ ( .D(n7836), .CK(clk), .Q(
        matrix_mul_2D_6__2__6_), .QN(n2663) );
  DFF_X1 matrix_mul_2D_reg_6__2__7_ ( .D(n7832), .CK(clk), .Q(
        matrix_mul_2D_6__2__7_), .QN(n2662) );
  DFF_X1 matrix_mul_2D_reg_6__2__8_ ( .D(n78280), .CK(clk), .Q(
        matrix_mul_2D_6__2__8_), .QN(n2661) );
  DFF_X1 matrix_mul_2D_reg_6__2__9_ ( .D(n78240), .CK(clk), .Q(
        matrix_mul_2D_6__2__9_), .QN(n2660) );
  DFF_X1 matrix_mul_2D_reg_6__2__10_ ( .D(n78200), .CK(clk), .Q(
        matrix_mul_2D_6__2__10_), .QN(n2659) );
  DFF_X1 matrix_mul_2D_reg_6__2__11_ ( .D(n78160), .CK(clk), .Q(
        matrix_mul_2D_6__2__11_), .QN(n2658) );
  DFF_X1 matrix_mul_2D_reg_6__2__12_ ( .D(n78120), .CK(clk), .Q(
        matrix_mul_2D_6__2__12_), .QN(n2657) );
  DFF_X1 matrix_mul_2D_reg_6__2__13_ ( .D(n78080), .CK(clk), .Q(
        matrix_mul_2D_6__2__13_), .QN(n265600) );
  DFF_X1 matrix_mul_2D_reg_6__2__14_ ( .D(n7804), .CK(clk), .Q(
        matrix_mul_2D_6__2__14_), .QN(n265500) );
  DFF_X1 matrix_mul_2D_reg_6__2__15_ ( .D(n7803), .CK(clk), .Q(
        matrix_mul_2D_6__2__15_), .QN(n17436) );
  DFF_X1 matrix_mul_2D_reg_6__2__16_ ( .D(n7802), .CK(clk), .Q(
        matrix_mul_2D_6__2__16_), .QN(n17434) );
  DFF_X1 matrix_mul_2D_reg_6__2__17_ ( .D(n7801), .CK(clk), .Q(
        matrix_mul_2D_6__2__17_), .QN(n17432) );
  DFF_X1 matrix_mul_2D_reg_6__2__18_ ( .D(n7800), .CK(clk), .Q(
        matrix_mul_2D_6__2__18_), .QN(n17430) );
  DFF_X1 matrix_mul_2D_reg_6__2__19_ ( .D(n7799), .CK(clk), .Q(
        matrix_mul_2D_6__2__19_), .QN(n17428) );
  DFF_X1 matrix_mul_2D_reg_6__2__20_ ( .D(n7798), .CK(clk), .Q(
        matrix_mul_2D_6__2__20_), .QN(n17426) );
  DFF_X1 matrix_mul_2D_reg_6__3__0_ ( .D(n7793), .CK(clk), .Q(
        matrix_mul_2D_6__3__0_), .QN(n268400) );
  DFF_X1 matrix_mul_2D_reg_6__3__1_ ( .D(n77890), .CK(clk), .Q(
        matrix_mul_2D_6__3__1_), .QN(n268300) );
  DFF_X1 matrix_mul_2D_reg_6__3__2_ ( .D(n77850), .CK(clk), .Q(
        matrix_mul_2D_6__3__2_), .QN(n268200) );
  DFF_X1 matrix_mul_2D_reg_6__3__3_ ( .D(n77810), .CK(clk), .Q(
        matrix_mul_2D_6__3__3_), .QN(n268100) );
  DFF_X1 matrix_mul_2D_reg_6__3__4_ ( .D(n77770), .CK(clk), .Q(
        matrix_mul_2D_6__3__4_), .QN(n268000) );
  DFF_X1 matrix_mul_2D_reg_6__3__5_ ( .D(n7773), .CK(clk), .Q(
        matrix_mul_2D_6__3__5_), .QN(n267900) );
  DFF_X1 matrix_mul_2D_reg_6__3__6_ ( .D(n7769), .CK(clk), .Q(
        matrix_mul_2D_6__3__6_), .QN(n267800) );
  DFF_X1 matrix_mul_2D_reg_6__3__7_ ( .D(n7765), .CK(clk), .Q(
        matrix_mul_2D_6__3__7_), .QN(n267700) );
  DFF_X1 matrix_mul_2D_reg_6__3__8_ ( .D(n7761), .CK(clk), .Q(
        matrix_mul_2D_6__3__8_), .QN(n267600) );
  DFF_X1 matrix_mul_2D_reg_6__3__9_ ( .D(n7757), .CK(clk), .Q(
        matrix_mul_2D_6__3__9_), .QN(n267500) );
  DFF_X1 matrix_mul_2D_reg_6__3__10_ ( .D(n7753), .CK(clk), .Q(
        matrix_mul_2D_6__3__10_), .QN(n267400) );
  DFF_X1 matrix_mul_2D_reg_6__3__11_ ( .D(n77490), .CK(clk), .Q(
        matrix_mul_2D_6__3__11_), .QN(n2673) );
  DFF_X1 matrix_mul_2D_reg_6__3__12_ ( .D(n77450), .CK(clk), .Q(
        matrix_mul_2D_6__3__12_), .QN(n2672) );
  DFF_X1 matrix_mul_2D_reg_6__3__13_ ( .D(n77410), .CK(clk), .Q(
        matrix_mul_2D_6__3__13_), .QN(n2671) );
  DFF_X1 matrix_mul_2D_reg_6__3__14_ ( .D(n77370), .CK(clk), .Q(
        matrix_mul_2D_6__3__14_), .QN(n2670) );
  DFF_X1 matrix_mul_2D_reg_6__3__15_ ( .D(n77360), .CK(clk), .Q(
        matrix_mul_2D_6__3__15_), .QN(n17424) );
  DFF_X1 matrix_mul_2D_reg_6__3__16_ ( .D(n77350), .CK(clk), .Q(
        matrix_mul_2D_6__3__16_), .QN(n17422) );
  DFF_X1 matrix_mul_2D_reg_6__3__17_ ( .D(n77340), .CK(clk), .Q(
        matrix_mul_2D_6__3__17_), .QN(n17420) );
  DFF_X1 matrix_mul_2D_reg_6__3__18_ ( .D(n77330), .CK(clk), .Q(
        matrix_mul_2D_6__3__18_), .QN(n17418) );
  DFF_X1 matrix_mul_2D_reg_6__3__19_ ( .D(n77320), .CK(clk), .Q(
        matrix_mul_2D_6__3__19_), .QN(n17416) );
  DFF_X1 matrix_mul_2D_reg_6__3__20_ ( .D(n77310), .CK(clk), .Q(
        matrix_mul_2D_6__3__20_), .QN(n17414) );
  DFF_X1 matrix_mul_2D_reg_6__4__0_ ( .D(n7726), .CK(clk), .Q(
        matrix_mul_2D_6__4__0_), .QN(n2705) );
  DFF_X1 matrix_mul_2D_reg_6__4__1_ ( .D(n7722), .CK(clk), .Q(
        matrix_mul_2D_6__4__1_), .QN(n2704) );
  DFF_X1 matrix_mul_2D_reg_6__4__2_ ( .D(n7718), .CK(clk), .Q(
        matrix_mul_2D_6__4__2_), .QN(n2703) );
  DFF_X1 matrix_mul_2D_reg_6__4__3_ ( .D(n7714), .CK(clk), .Q(
        matrix_mul_2D_6__4__3_), .QN(n2702) );
  DFF_X1 matrix_mul_2D_reg_6__4__4_ ( .D(n77100), .CK(clk), .Q(
        matrix_mul_2D_6__4__4_), .QN(n2701) );
  DFF_X1 matrix_mul_2D_reg_6__4__5_ ( .D(n77060), .CK(clk), .Q(
        matrix_mul_2D_6__4__5_), .QN(n2700) );
  DFF_X1 matrix_mul_2D_reg_6__4__6_ ( .D(n77020), .CK(clk), .Q(
        matrix_mul_2D_6__4__6_), .QN(n2699) );
  DFF_X1 matrix_mul_2D_reg_6__4__7_ ( .D(n76980), .CK(clk), .Q(
        matrix_mul_2D_6__4__7_), .QN(n2698) );
  DFF_X1 matrix_mul_2D_reg_6__4__8_ ( .D(n7694), .CK(clk), .Q(
        matrix_mul_2D_6__4__8_), .QN(n2697) );
  DFF_X1 matrix_mul_2D_reg_6__4__9_ ( .D(n7690), .CK(clk), .Q(
        matrix_mul_2D_6__4__9_), .QN(n2696) );
  DFF_X1 matrix_mul_2D_reg_6__4__10_ ( .D(n7686), .CK(clk), .Q(
        matrix_mul_2D_6__4__10_), .QN(n2695) );
  DFF_X1 matrix_mul_2D_reg_6__4__11_ ( .D(n7682), .CK(clk), .Q(
        matrix_mul_2D_6__4__11_), .QN(n269400) );
  DFF_X1 matrix_mul_2D_reg_6__4__12_ ( .D(n7678), .CK(clk), .Q(
        matrix_mul_2D_6__4__12_), .QN(n269300) );
  DFF_X1 matrix_mul_2D_reg_6__4__13_ ( .D(n7674), .CK(clk), .Q(
        matrix_mul_2D_6__4__13_), .QN(n269200) );
  DFF_X1 matrix_mul_2D_reg_6__4__14_ ( .D(n7670), .CK(clk), .Q(
        matrix_mul_2D_6__4__14_), .QN(n269100) );
  DFF_X1 matrix_mul_2D_reg_6__4__15_ ( .D(n7669), .CK(clk), .Q(
        matrix_mul_2D_6__4__15_), .QN(n17412) );
  DFF_X1 matrix_mul_2D_reg_6__4__16_ ( .D(n7668), .CK(clk), .Q(
        matrix_mul_2D_6__4__16_), .QN(n17410) );
  DFF_X1 matrix_mul_2D_reg_6__4__17_ ( .D(n7667), .CK(clk), .Q(
        matrix_mul_2D_6__4__17_), .QN(n17408) );
  DFF_X1 matrix_mul_2D_reg_6__4__18_ ( .D(n7666), .CK(clk), .Q(
        matrix_mul_2D_6__4__18_), .QN(n17406) );
  DFF_X1 matrix_mul_2D_reg_6__4__19_ ( .D(n7665), .CK(clk), .Q(
        matrix_mul_2D_6__4__19_), .QN(n17404) );
  DFF_X1 matrix_mul_2D_reg_6__4__20_ ( .D(n7664), .CK(clk), .Q(
        matrix_mul_2D_6__4__20_), .QN(n17402) );
  DFF_X1 matrix_mul_2D_reg_6__5__0_ ( .D(n76600), .CK(clk), .Q(
        matrix_mul_2D_6__5__0_), .QN(n2720) );
  DFF_X1 matrix_mul_2D_reg_6__5__1_ ( .D(n76550), .CK(clk), .Q(
        matrix_mul_2D_6__5__1_), .QN(n2719) );
  DFF_X1 matrix_mul_2D_reg_6__5__2_ ( .D(n76500), .CK(clk), .Q(
        matrix_mul_2D_6__5__2_), .QN(n2718) );
  DFF_X1 matrix_mul_2D_reg_6__5__3_ ( .D(n76450), .CK(clk), .Q(
        matrix_mul_2D_6__5__3_), .QN(n2717) );
  DFF_X1 matrix_mul_2D_reg_6__5__4_ ( .D(n76400), .CK(clk), .Q(
        matrix_mul_2D_6__5__4_), .QN(n2716) );
  DFF_X1 matrix_mul_2D_reg_6__5__5_ ( .D(n7635), .CK(clk), .Q(
        matrix_mul_2D_6__5__5_), .QN(n2715) );
  DFF_X1 matrix_mul_2D_reg_6__5__6_ ( .D(n7630), .CK(clk), .Q(
        matrix_mul_2D_6__5__6_), .QN(n2714) );
  DFF_X1 matrix_mul_2D_reg_6__5__7_ ( .D(n7625), .CK(clk), .Q(
        matrix_mul_2D_6__5__7_), .QN(n2713) );
  DFF_X1 matrix_mul_2D_reg_6__5__8_ ( .D(n76200), .CK(clk), .Q(
        matrix_mul_2D_6__5__8_), .QN(n2712) );
  DFF_X1 matrix_mul_2D_reg_6__5__9_ ( .D(n76150), .CK(clk), .Q(
        matrix_mul_2D_6__5__9_), .QN(n2711) );
  DFF_X1 matrix_mul_2D_reg_6__5__10_ ( .D(n76100), .CK(clk), .Q(
        matrix_mul_2D_6__5__10_), .QN(n2710) );
  DFF_X1 matrix_mul_2D_reg_6__5__11_ ( .D(n7605), .CK(clk), .Q(
        matrix_mul_2D_6__5__11_), .QN(n2709) );
  DFF_X1 matrix_mul_2D_reg_6__5__12_ ( .D(n7600), .CK(clk), .Q(
        matrix_mul_2D_6__5__12_), .QN(n2708) );
  DFF_X1 matrix_mul_2D_reg_6__5__13_ ( .D(n7595), .CK(clk), .Q(
        matrix_mul_2D_6__5__13_), .QN(n2707) );
  DFF_X1 matrix_mul_2D_reg_6__5__14_ ( .D(n7590), .CK(clk), .Q(
        matrix_mul_2D_6__5__14_), .QN(n2706) );
  DFF_X1 matrix_mul_2D_reg_6__5__15_ ( .D(n7589), .CK(clk), .Q(
        matrix_mul_2D_6__5__15_), .QN(n17400) );
  DFF_X1 matrix_mul_2D_reg_6__5__16_ ( .D(n7588), .CK(clk), .Q(
        matrix_mul_2D_6__5__16_), .QN(n17398) );
  DFF_X1 matrix_mul_2D_reg_6__5__17_ ( .D(n7587), .CK(clk), .Q(
        matrix_mul_2D_6__5__17_), .QN(n17396) );
  DFF_X1 matrix_mul_2D_reg_6__5__18_ ( .D(n7586), .CK(clk), .Q(
        matrix_mul_2D_6__5__18_), .QN(n17394) );
  DFF_X1 matrix_mul_2D_reg_6__5__19_ ( .D(n7585), .CK(clk), .Q(
        matrix_mul_2D_6__5__19_), .QN(n17392) );
  DFF_X1 matrix_mul_2D_reg_6__5__20_ ( .D(n7584), .CK(clk), .Q(
        matrix_mul_2D_6__5__20_), .QN(n17390) );
  DFF_X1 matrix_mul_2D_reg_6__6__0_ ( .D(n75790), .CK(clk), .Q(
        matrix_mul_2D_6__6__0_), .QN(n273500) );
  DFF_X1 matrix_mul_2D_reg_6__6__1_ ( .D(n75750), .CK(clk), .Q(
        matrix_mul_2D_6__6__1_), .QN(n273400) );
  DFF_X1 matrix_mul_2D_reg_6__6__2_ ( .D(n75710), .CK(clk), .Q(
        matrix_mul_2D_6__6__2_), .QN(n273300) );
  DFF_X1 matrix_mul_2D_reg_6__6__3_ ( .D(n75670), .CK(clk), .Q(
        matrix_mul_2D_6__6__3_), .QN(n2732) );
  DFF_X1 matrix_mul_2D_reg_6__6__4_ ( .D(n75630), .CK(clk), .Q(
        matrix_mul_2D_6__6__4_), .QN(n2731) );
  DFF_X1 matrix_mul_2D_reg_6__6__5_ ( .D(n7559), .CK(clk), .Q(
        matrix_mul_2D_6__6__5_), .QN(n2730) );
  DFF_X1 matrix_mul_2D_reg_6__6__6_ ( .D(n7555), .CK(clk), .Q(
        matrix_mul_2D_6__6__6_), .QN(n272900) );
  DFF_X1 matrix_mul_2D_reg_6__6__7_ ( .D(n7551), .CK(clk), .Q(
        matrix_mul_2D_6__6__7_), .QN(n2728) );
  DFF_X1 matrix_mul_2D_reg_6__6__8_ ( .D(n7547), .CK(clk), .Q(
        matrix_mul_2D_6__6__8_), .QN(n2727) );
  DFF_X1 matrix_mul_2D_reg_6__6__9_ ( .D(n75430), .CK(clk), .Q(
        matrix_mul_2D_6__6__9_), .QN(n2726) );
  DFF_X1 matrix_mul_2D_reg_6__6__10_ ( .D(n75390), .CK(clk), .Q(
        matrix_mul_2D_6__6__10_), .QN(n2725) );
  DFF_X1 matrix_mul_2D_reg_6__6__11_ ( .D(n75350), .CK(clk), .Q(
        matrix_mul_2D_6__6__11_), .QN(n2724) );
  DFF_X1 matrix_mul_2D_reg_6__6__12_ ( .D(n75310), .CK(clk), .Q(
        matrix_mul_2D_6__6__12_), .QN(n2723) );
  DFF_X1 matrix_mul_2D_reg_6__6__13_ ( .D(n7527), .CK(clk), .Q(
        matrix_mul_2D_6__6__13_), .QN(n2722) );
  DFF_X1 matrix_mul_2D_reg_6__6__14_ ( .D(n7523), .CK(clk), .Q(
        matrix_mul_2D_6__6__14_), .QN(n2721) );
  DFF_X1 matrix_mul_2D_reg_6__6__15_ ( .D(n7522), .CK(clk), .Q(
        matrix_mul_2D_6__6__15_), .QN(n17388) );
  DFF_X1 matrix_mul_2D_reg_6__6__16_ ( .D(n7521), .CK(clk), .Q(
        matrix_mul_2D_6__6__16_), .QN(n17386) );
  DFF_X1 matrix_mul_2D_reg_6__6__17_ ( .D(n7520), .CK(clk), .Q(
        matrix_mul_2D_6__6__17_), .QN(n17384) );
  DFF_X1 matrix_mul_2D_reg_6__6__18_ ( .D(n7519), .CK(clk), .Q(
        matrix_mul_2D_6__6__18_), .QN(n17382) );
  DFF_X1 matrix_mul_2D_reg_6__6__19_ ( .D(n7518), .CK(clk), .Q(
        matrix_mul_2D_6__6__19_), .QN(n17380) );
  DFF_X1 matrix_mul_2D_reg_6__6__20_ ( .D(n7517), .CK(clk), .Q(
        matrix_mul_2D_6__6__20_), .QN(n17378) );
  DFF_X1 matrix_mul_2D_reg_6__7__13_ ( .D(n7512), .CK(clk), .Q(
        matrix_mul_2D_6__7__13_), .QN(n273700) );
  DFF_X1 matrix_mul_2D_reg_6__7__15_ ( .D(n7511), .CK(clk), .Q(
        matrix_mul_2D_6__7__15_), .QN(n17376) );
  DFF_X1 matrix_mul_2D_reg_6__7__16_ ( .D(n7510), .CK(clk), .Q(
        matrix_mul_2D_6__7__16_), .QN(n17374) );
  DFF_X1 matrix_mul_2D_reg_6__7__17_ ( .D(n7509), .CK(clk), .Q(
        matrix_mul_2D_6__7__17_), .QN(n17372) );
  DFF_X1 matrix_mul_2D_reg_6__7__18_ ( .D(n7508), .CK(clk), .Q(
        matrix_mul_2D_6__7__18_), .QN(n17370) );
  DFF_X1 matrix_mul_2D_reg_6__7__19_ ( .D(n7507), .CK(clk), .Q(
        matrix_mul_2D_6__7__19_), .QN(n17368) );
  DFF_X1 matrix_mul_2D_reg_6__7__20_ ( .D(n7506), .CK(clk), .Q(
        matrix_mul_2D_6__7__20_), .QN(n17366) );
  DFF_X1 matrix_mul_2D_reg_7__0__0_ ( .D(n7502), .CK(clk), .Q(
        matrix_mul_2D_7__0__0_), .QN(n2765) );
  DFF_X1 matrix_mul_2D_reg_7__0__1_ ( .D(n7497), .CK(clk), .Q(
        matrix_mul_2D_7__0__1_), .QN(n2764) );
  DFF_X1 matrix_mul_2D_reg_7__0__2_ ( .D(n74920), .CK(clk), .Q(
        matrix_mul_2D_7__0__2_), .QN(n2763) );
  DFF_X1 matrix_mul_2D_reg_7__0__3_ ( .D(n74870), .CK(clk), .Q(
        matrix_mul_2D_7__0__3_), .QN(n2762) );
  DFF_X1 matrix_mul_2D_reg_7__0__4_ ( .D(n74820), .CK(clk), .Q(
        matrix_mul_2D_7__0__4_), .QN(n2761) );
  DFF_X1 matrix_mul_2D_reg_7__0__5_ ( .D(n74770), .CK(clk), .Q(
        matrix_mul_2D_7__0__5_), .QN(n2760) );
  DFF_X1 matrix_mul_2D_reg_7__0__6_ ( .D(n74720), .CK(clk), .Q(
        matrix_mul_2D_7__0__6_), .QN(n2759) );
  DFF_X1 matrix_mul_2D_reg_7__0__7_ ( .D(n7467), .CK(clk), .Q(
        matrix_mul_2D_7__0__7_), .QN(n2758) );
  DFF_X1 matrix_mul_2D_reg_7__0__8_ ( .D(n7462), .CK(clk), .Q(
        matrix_mul_2D_7__0__8_), .QN(n2757) );
  DFF_X1 matrix_mul_2D_reg_7__0__9_ ( .D(n7457), .CK(clk), .Q(
        matrix_mul_2D_7__0__9_), .QN(n2756) );
  DFF_X1 matrix_mul_2D_reg_7__0__10_ ( .D(n74520), .CK(clk), .Q(
        matrix_mul_2D_7__0__10_), .QN(n2755) );
  DFF_X1 matrix_mul_2D_reg_7__0__11_ ( .D(n74470), .CK(clk), .Q(
        matrix_mul_2D_7__0__11_), .QN(n2754) );
  DFF_X1 matrix_mul_2D_reg_7__0__12_ ( .D(n74420), .CK(clk), .Q(
        matrix_mul_2D_7__0__12_), .QN(n2753) );
  DFF_X1 matrix_mul_2D_reg_7__0__13_ ( .D(n7437), .CK(clk), .Q(
        matrix_mul_2D_7__0__13_), .QN(n2752) );
  DFF_X1 matrix_mul_2D_reg_7__0__14_ ( .D(n7432), .CK(clk), .Q(
        matrix_mul_2D_7__0__14_), .QN(n2751) );
  DFF_X1 matrix_mul_2D_reg_7__0__15_ ( .D(n7431), .CK(clk), .Q(
        matrix_mul_2D_7__0__15_), .QN(n17364) );
  DFF_X1 matrix_mul_2D_reg_7__0__16_ ( .D(n7430), .CK(clk), .Q(
        matrix_mul_2D_7__0__16_), .QN(n17362) );
  DFF_X1 matrix_mul_2D_reg_7__0__17_ ( .D(n7429), .CK(clk), .Q(
        matrix_mul_2D_7__0__17_), .QN(n17360) );
  DFF_X1 matrix_mul_2D_reg_7__0__18_ ( .D(n7428), .CK(clk), .Q(
        matrix_mul_2D_7__0__18_), .QN(n17358) );
  DFF_X1 matrix_mul_2D_reg_7__0__19_ ( .D(n7427), .CK(clk), .Q(
        matrix_mul_2D_7__0__19_), .QN(n17356) );
  DFF_X1 matrix_mul_2D_reg_7__0__20_ ( .D(n7426), .CK(clk), .Q(
        matrix_mul_2D_7__0__20_), .QN(n17354) );
  DFF_X1 matrix_mul_2D_reg_7__1__0_ ( .D(n7422), .CK(clk), .Q(
        matrix_mul_2D_7__1__0_), .QN(n278000) );
  DFF_X1 matrix_mul_2D_reg_7__1__1_ ( .D(n7417), .CK(clk), .Q(
        matrix_mul_2D_7__1__1_), .QN(n277900) );
  DFF_X1 matrix_mul_2D_reg_7__1__2_ ( .D(n74120), .CK(clk), .Q(
        matrix_mul_2D_7__1__2_), .QN(n277800) );
  DFF_X1 matrix_mul_2D_reg_7__1__3_ ( .D(n5296), .CK(clk), .Q(
        matrix_mul_2D_7__1__3_), .QN(n277700) );
  DFF_X1 matrix_mul_2D_reg_7__1__4_ ( .D(n4888), .CK(clk), .Q(
        matrix_mul_2D_7__1__4_), .QN(n277600) );
  DFF_X1 matrix_mul_2D_reg_7__1__5_ ( .D(n47080), .CK(clk), .Q(
        matrix_mul_2D_7__1__5_), .QN(n277500) );
  DFF_X1 matrix_mul_2D_reg_7__1__6_ ( .D(n43540), .CK(clk), .Q(
        matrix_mul_2D_7__1__6_), .QN(n277400) );
  DFF_X1 matrix_mul_2D_reg_7__1__7_ ( .D(n3617), .CK(clk), .Q(
        matrix_mul_2D_7__1__7_), .QN(n277300) );
  DFF_X1 matrix_mul_2D_reg_7__1__8_ ( .D(n32530), .CK(clk), .Q(
        matrix_mul_2D_7__1__8_), .QN(n277200) );
  DFF_X1 matrix_mul_2D_reg_7__1__9_ ( .D(n3153), .CK(clk), .Q(
        matrix_mul_2D_7__1__9_), .QN(n277100) );
  DFF_X1 matrix_mul_2D_reg_7__1__10_ ( .D(n3100), .CK(clk), .Q(
        matrix_mul_2D_7__1__10_), .QN(n277000) );
  DFF_X1 matrix_mul_2D_reg_7__1__11_ ( .D(n3067), .CK(clk), .Q(
        matrix_mul_2D_7__1__11_), .QN(n276900) );
  DFF_X1 matrix_mul_2D_reg_7__1__12_ ( .D(n3062), .CK(clk), .Q(
        matrix_mul_2D_7__1__12_), .QN(n276800) );
  DFF_X1 matrix_mul_2D_reg_7__1__13_ ( .D(n3057), .CK(clk), .Q(
        matrix_mul_2D_7__1__13_), .QN(n276700) );
  DFF_X1 matrix_mul_2D_reg_7__1__14_ ( .D(n3052), .CK(clk), .Q(
        matrix_mul_2D_7__1__14_), .QN(n276600) );
  DFF_X1 matrix_mul_2D_reg_7__1__15_ ( .D(n3051), .CK(clk), .Q(
        matrix_mul_2D_7__1__15_), .QN(n17352) );
  DFF_X1 matrix_mul_2D_reg_7__1__16_ ( .D(n3050), .CK(clk), .Q(
        matrix_mul_2D_7__1__16_), .QN(n17350) );
  DFF_X1 matrix_mul_2D_reg_7__1__17_ ( .D(n3049), .CK(clk), .Q(
        matrix_mul_2D_7__1__17_), .QN(n17348) );
  DFF_X1 matrix_mul_2D_reg_7__1__18_ ( .D(n3048), .CK(clk), .Q(
        matrix_mul_2D_7__1__18_), .QN(n17346) );
  DFF_X1 matrix_mul_2D_reg_7__1__19_ ( .D(n3047), .CK(clk), .Q(
        matrix_mul_2D_7__1__19_), .QN(n17344) );
  DFF_X1 matrix_mul_2D_reg_7__1__20_ ( .D(n3046), .CK(clk), .Q(
        matrix_mul_2D_7__1__20_), .QN(n17342) );
  DFF_X1 matrix_mul_2D_reg_7__2__0_ ( .D(n30410), .CK(clk), .Q(
        matrix_mul_2D_7__2__0_), .QN(n2801) );
  DFF_X1 matrix_mul_2D_reg_7__2__1_ ( .D(n30370), .CK(clk), .Q(
        matrix_mul_2D_7__2__1_), .QN(n2800) );
  DFF_X1 matrix_mul_2D_reg_7__2__2_ ( .D(n30330), .CK(clk), .Q(
        matrix_mul_2D_7__2__2_), .QN(n2799) );
  DFF_X1 matrix_mul_2D_reg_7__2__3_ ( .D(n30290), .CK(clk), .Q(
        matrix_mul_2D_7__2__3_), .QN(n2798) );
  DFF_X1 matrix_mul_2D_reg_7__2__4_ ( .D(n30250), .CK(clk), .Q(
        matrix_mul_2D_7__2__4_), .QN(n2797) );
  DFF_X1 matrix_mul_2D_reg_7__2__5_ ( .D(n3021), .CK(clk), .Q(
        matrix_mul_2D_7__2__5_), .QN(n2796) );
  DFF_X1 matrix_mul_2D_reg_7__2__6_ ( .D(n3017), .CK(clk), .Q(
        matrix_mul_2D_7__2__6_), .QN(n2795) );
  DFF_X1 matrix_mul_2D_reg_7__2__7_ ( .D(n3013), .CK(clk), .Q(
        matrix_mul_2D_7__2__7_), .QN(n2794) );
  DFF_X1 matrix_mul_2D_reg_7__2__8_ ( .D(n3009), .CK(clk), .Q(
        matrix_mul_2D_7__2__8_), .QN(n2793) );
  DFF_X1 matrix_mul_2D_reg_7__2__9_ ( .D(n3005), .CK(clk), .Q(
        matrix_mul_2D_7__2__9_), .QN(n2792) );
  DFF_X1 matrix_mul_2D_reg_7__2__10_ ( .D(n30010), .CK(clk), .Q(
        matrix_mul_2D_7__2__10_), .QN(n2791) );
  DFF_X1 matrix_mul_2D_reg_7__2__11_ ( .D(n29970), .CK(clk), .Q(
        matrix_mul_2D_7__2__11_), .QN(n2790) );
  DFF_X1 matrix_mul_2D_reg_7__2__12_ ( .D(n29930), .CK(clk), .Q(
        matrix_mul_2D_7__2__12_), .QN(n2789) );
  DFF_X1 matrix_mul_2D_reg_7__2__13_ ( .D(n29890), .CK(clk), .Q(
        matrix_mul_2D_7__2__13_), .QN(n2788) );
  DFF_X1 matrix_mul_2D_reg_7__2__14_ ( .D(n29850), .CK(clk), .Q(
        matrix_mul_2D_7__2__14_), .QN(n2787) );
  DFF_X1 matrix_mul_2D_reg_7__2__15_ ( .D(n2984), .CK(clk), .Q(
        matrix_mul_2D_7__2__15_), .QN(n17340) );
  DFF_X1 matrix_mul_2D_reg_7__2__16_ ( .D(n2983), .CK(clk), .Q(
        matrix_mul_2D_7__2__16_), .QN(n17338) );
  DFF_X1 matrix_mul_2D_reg_7__2__17_ ( .D(n2982), .CK(clk), .Q(
        matrix_mul_2D_7__2__17_), .QN(n17336) );
  DFF_X1 matrix_mul_2D_reg_7__2__18_ ( .D(n2981), .CK(clk), .Q(
        matrix_mul_2D_7__2__18_), .QN(n17334) );
  DFF_X1 matrix_mul_2D_reg_7__2__19_ ( .D(n2980), .CK(clk), .Q(
        matrix_mul_2D_7__2__19_), .QN(n17332) );
  DFF_X1 matrix_mul_2D_reg_7__2__20_ ( .D(n2979), .CK(clk), .Q(
        matrix_mul_2D_7__2__20_), .QN(n17330) );
  DFF_X1 matrix_mul_2D_reg_7__3__0_ ( .D(n2974), .CK(clk), .Q(
        matrix_mul_2D_7__3__0_), .QN(n28160) );
  DFF_X1 matrix_mul_2D_reg_7__3__1_ ( .D(n2970), .CK(clk), .Q(
        matrix_mul_2D_7__3__1_), .QN(n28150) );
  DFF_X1 matrix_mul_2D_reg_7__3__2_ ( .D(n2966), .CK(clk), .Q(
        matrix_mul_2D_7__3__2_), .QN(n2814) );
  DFF_X1 matrix_mul_2D_reg_7__3__3_ ( .D(n2962), .CK(clk), .Q(
        matrix_mul_2D_7__3__3_), .QN(n2813) );
  DFF_X1 matrix_mul_2D_reg_7__3__4_ ( .D(n29580), .CK(clk), .Q(
        matrix_mul_2D_7__3__4_), .QN(n2812) );
  DFF_X1 matrix_mul_2D_reg_7__3__5_ ( .D(n29540), .CK(clk), .Q(
        matrix_mul_2D_7__3__5_), .QN(n28110) );
  DFF_X1 matrix_mul_2D_reg_7__3__6_ ( .D(n29500), .CK(clk), .Q(
        matrix_mul_2D_7__3__6_), .QN(n2810) );
  DFF_X1 matrix_mul_2D_reg_7__3__7_ ( .D(n29460), .CK(clk), .Q(
        matrix_mul_2D_7__3__7_), .QN(n2809) );
  DFF_X1 matrix_mul_2D_reg_7__3__8_ ( .D(n29420), .CK(clk), .Q(
        matrix_mul_2D_7__3__8_), .QN(n2808) );
  DFF_X1 matrix_mul_2D_reg_7__3__9_ ( .D(n2938), .CK(clk), .Q(
        matrix_mul_2D_7__3__9_), .QN(n2807) );
  DFF_X1 matrix_mul_2D_reg_7__3__10_ ( .D(n2934), .CK(clk), .Q(
        matrix_mul_2D_7__3__10_), .QN(n2806) );
  DFF_X1 matrix_mul_2D_reg_7__3__11_ ( .D(n2930), .CK(clk), .Q(
        matrix_mul_2D_7__3__11_), .QN(n2805) );
  DFF_X1 matrix_mul_2D_reg_7__3__12_ ( .D(n2926), .CK(clk), .Q(
        matrix_mul_2D_7__3__12_), .QN(n2804) );
  DFF_X1 matrix_mul_2D_reg_7__3__13_ ( .D(n29220), .CK(clk), .Q(
        matrix_mul_2D_7__3__13_), .QN(n2803) );
  DFF_X1 matrix_mul_2D_reg_7__3__14_ ( .D(n29180), .CK(clk), .Q(
        matrix_mul_2D_7__3__14_), .QN(n2802) );
  DFF_X1 matrix_mul_2D_reg_7__3__15_ ( .D(n29170), .CK(clk), .Q(
        matrix_mul_2D_7__3__15_), .QN(n17328) );
  DFF_X1 matrix_mul_2D_reg_7__3__16_ ( .D(n29160), .CK(clk), .Q(
        matrix_mul_2D_7__3__16_), .QN(n17326) );
  DFF_X1 matrix_mul_2D_reg_7__3__17_ ( .D(n29150), .CK(clk), .Q(
        matrix_mul_2D_7__3__17_), .QN(n17324) );
  DFF_X1 matrix_mul_2D_reg_7__3__18_ ( .D(n29140), .CK(clk), .Q(
        matrix_mul_2D_7__3__18_), .QN(n17322) );
  DFF_X1 matrix_mul_2D_reg_7__3__19_ ( .D(n29130), .CK(clk), .Q(
        matrix_mul_2D_7__3__19_), .QN(n17320) );
  DFF_X1 matrix_mul_2D_reg_7__3__20_ ( .D(n29120), .CK(clk), .Q(
        matrix_mul_2D_7__3__20_), .QN(n17318) );
  DFF_X1 matrix_mul_2D_reg_7__4__0_ ( .D(n29070), .CK(clk), .Q(
        matrix_mul_2D_7__4__0_), .QN(n2837) );
  DFF_X1 matrix_mul_2D_reg_7__4__1_ ( .D(n29030), .CK(clk), .Q(
        matrix_mul_2D_7__4__1_), .QN(n2836) );
  DFF_X1 matrix_mul_2D_reg_7__4__2_ ( .D(n2899), .CK(clk), .Q(
        matrix_mul_2D_7__4__2_), .QN(n2835) );
  DFF_X1 matrix_mul_2D_reg_7__4__3_ ( .D(n2895), .CK(clk), .Q(
        matrix_mul_2D_7__4__3_), .QN(n2834) );
  DFF_X1 matrix_mul_2D_reg_7__4__4_ ( .D(n2891), .CK(clk), .Q(
        matrix_mul_2D_7__4__4_), .QN(n2833) );
  DFF_X1 matrix_mul_2D_reg_7__4__5_ ( .D(n2887), .CK(clk), .Q(
        matrix_mul_2D_7__4__5_), .QN(n2832) );
  DFF_X1 matrix_mul_2D_reg_7__4__6_ ( .D(n2883), .CK(clk), .Q(
        matrix_mul_2D_7__4__6_), .QN(n2831) );
  DFF_X1 matrix_mul_2D_reg_7__4__7_ ( .D(n28190), .CK(clk), .Q(
        matrix_mul_2D_7__4__7_), .QN(n28300) );
  DFF_X1 matrix_mul_2D_reg_7__4__8_ ( .D(n278500), .CK(clk), .Q(
        matrix_mul_2D_7__4__8_), .QN(n28290) );
  DFF_X1 matrix_mul_2D_reg_7__4__9_ ( .D(n278100), .CK(clk), .Q(
        matrix_mul_2D_7__4__9_), .QN(n28280) );
  DFF_X1 matrix_mul_2D_reg_7__4__10_ ( .D(n268700), .CK(clk), .Q(
        matrix_mul_2D_7__4__10_), .QN(n28270) );
  DFF_X1 matrix_mul_2D_reg_7__4__11_ ( .D(n265300), .CK(clk), .Q(
        matrix_mul_2D_7__4__11_), .QN(n28260) );
  DFF_X1 matrix_mul_2D_reg_7__4__12_ ( .D(n264900), .CK(clk), .Q(
        matrix_mul_2D_7__4__12_), .QN(n28250) );
  DFF_X1 matrix_mul_2D_reg_7__4__13_ ( .D(n2555), .CK(clk), .Q(
        matrix_mul_2D_7__4__13_), .QN(n28240) );
  DFF_X1 matrix_mul_2D_reg_7__4__14_ ( .D(n2431), .CK(clk), .Q(
        matrix_mul_2D_7__4__14_), .QN(n28230) );
  DFF_X1 matrix_mul_2D_reg_7__4__15_ ( .D(n2430), .CK(clk), .Q(
        matrix_mul_2D_7__4__15_), .QN(n17316) );
  DFF_X1 matrix_mul_2D_reg_7__4__16_ ( .D(n2429), .CK(clk), .Q(
        matrix_mul_2D_7__4__16_), .QN(n17314) );
  DFF_X1 matrix_mul_2D_reg_7__4__17_ ( .D(n2428), .CK(clk), .Q(
        matrix_mul_2D_7__4__17_), .QN(n17312) );
  DFF_X1 matrix_mul_2D_reg_7__4__18_ ( .D(n2427), .CK(clk), .Q(
        matrix_mul_2D_7__4__18_), .QN(n17310) );
  DFF_X1 matrix_mul_2D_reg_7__4__19_ ( .D(n2291), .CK(clk), .Q(
        matrix_mul_2D_7__4__19_), .QN(n17308) );
  DFF_X1 matrix_mul_2D_reg_7__4__20_ ( .D(n2290), .CK(clk), .Q(
        matrix_mul_2D_7__4__20_), .QN(n17306) );
  DFF_X1 matrix_mul_2D_reg_7__5__0_ ( .D(n2210), .CK(clk), .Q(
        matrix_mul_2D_7__5__0_), .QN(n28520) );
  DFF_X1 matrix_mul_2D_reg_7__5__1_ ( .D(n2206), .CK(clk), .Q(
        matrix_mul_2D_7__5__1_), .QN(n28510) );
  DFF_X1 matrix_mul_2D_reg_7__5__2_ ( .D(n1923), .CK(clk), .Q(
        matrix_mul_2D_7__5__2_), .QN(n28500) );
  DFF_X1 matrix_mul_2D_reg_7__5__3_ ( .D(n948), .CK(clk), .Q(
        matrix_mul_2D_7__5__3_), .QN(n28490) );
  DFF_X1 matrix_mul_2D_reg_7__5__4_ ( .D(n944), .CK(clk), .Q(
        matrix_mul_2D_7__5__4_), .QN(n28480) );
  DFF_X1 matrix_mul_2D_reg_7__5__5_ ( .D(n940), .CK(clk), .Q(
        matrix_mul_2D_7__5__5_), .QN(n2847) );
  DFF_X1 matrix_mul_2D_reg_7__5__6_ ( .D(n936), .CK(clk), .Q(
        matrix_mul_2D_7__5__6_), .QN(n2846) );
  DFF_X1 matrix_mul_2D_reg_7__5__7_ ( .D(n932), .CK(clk), .Q(
        matrix_mul_2D_7__5__7_), .QN(n2845) );
  DFF_X1 matrix_mul_2D_reg_7__5__8_ ( .D(n928), .CK(clk), .Q(
        matrix_mul_2D_7__5__8_), .QN(n2844) );
  DFF_X1 matrix_mul_2D_reg_7__5__9_ ( .D(n924), .CK(clk), .Q(
        matrix_mul_2D_7__5__9_), .QN(n2843) );
  DFF_X1 matrix_mul_2D_reg_7__5__10_ ( .D(n920), .CK(clk), .Q(
        matrix_mul_2D_7__5__10_), .QN(n2842) );
  DFF_X1 matrix_mul_2D_reg_7__5__11_ ( .D(n916), .CK(clk), .Q(
        matrix_mul_2D_7__5__11_), .QN(n2841) );
  DFF_X1 matrix_mul_2D_reg_7__5__12_ ( .D(n912), .CK(clk), .Q(
        matrix_mul_2D_7__5__12_), .QN(n2840) );
  DFF_X1 matrix_mul_2D_reg_7__5__13_ ( .D(n908), .CK(clk), .Q(
        matrix_mul_2D_7__5__13_), .QN(n2839) );
  DFF_X1 matrix_mul_2D_reg_7__5__14_ ( .D(n904), .CK(clk), .Q(
        matrix_mul_2D_7__5__14_), .QN(n2838) );
  DFF_X1 matrix_mul_2D_reg_7__5__15_ ( .D(n903), .CK(clk), .Q(
        matrix_mul_2D_7__5__15_), .QN(n17304) );
  DFF_X1 matrix_mul_2D_reg_7__5__16_ ( .D(n902), .CK(clk), .Q(
        matrix_mul_2D_7__5__16_), .QN(n17302) );
  DFF_X1 matrix_mul_2D_reg_7__5__17_ ( .D(n901), .CK(clk), .Q(
        matrix_mul_2D_7__5__17_), .QN(n17300) );
  DFF_X1 matrix_mul_2D_reg_7__5__18_ ( .D(n900), .CK(clk), .Q(
        matrix_mul_2D_7__5__18_), .QN(n17298) );
  DFF_X1 matrix_mul_2D_reg_7__5__19_ ( .D(n899), .CK(clk), .Q(
        matrix_mul_2D_7__5__19_), .QN(n17296) );
  DFF_X1 matrix_mul_2D_reg_7__5__20_ ( .D(n898), .CK(clk), .Q(
        matrix_mul_2D_7__5__20_), .QN(n17294) );
  DFF_X1 matrix_mul_2D_reg_7__6__15_ ( .D(n897), .CK(clk), .Q(
        matrix_mul_2D_7__6__15_), .QN(n17292) );
  DFF_X1 matrix_mul_2D_reg_7__6__16_ ( .D(n896), .CK(clk), .Q(
        matrix_mul_2D_7__6__16_), .QN(n17290) );
  DFF_X1 matrix_mul_2D_reg_7__6__17_ ( .D(n895), .CK(clk), .Q(
        matrix_mul_2D_7__6__17_), .QN(n17288) );
  DFF_X1 matrix_mul_2D_reg_7__6__18_ ( .D(n894), .CK(clk), .Q(
        matrix_mul_2D_7__6__18_), .QN(n17286) );
  DFF_X1 matrix_mul_2D_reg_7__6__19_ ( .D(n893), .CK(clk), .Q(
        matrix_mul_2D_7__6__19_), .QN(n17284) );
  DFF_X1 matrix_mul_2D_reg_7__6__20_ ( .D(n892), .CK(clk), .Q(
        matrix_mul_2D_7__6__20_), .QN(n17282) );
  DFF_X1 matrix_mul_2D_reg_7__7__15_ ( .D(n891), .CK(clk), .Q(
        matrix_mul_2D_7__7__15_), .QN(n17280) );
  DFF_X1 matrix_mul_2D_reg_7__7__16_ ( .D(n890), .CK(clk), .Q(
        matrix_mul_2D_7__7__16_), .QN(n17278) );
  DFF_X1 matrix_mul_2D_reg_7__7__17_ ( .D(n889), .CK(clk), .Q(
        matrix_mul_2D_7__7__17_), .QN(n17276) );
  DFF_X1 matrix_mul_2D_reg_7__7__18_ ( .D(n888), .CK(clk), .Q(
        matrix_mul_2D_7__7__18_), .QN(n17274) );
  DFF_X1 matrix_mul_2D_reg_7__7__19_ ( .D(n887), .CK(clk), .Q(
        matrix_mul_2D_7__7__19_), .QN(n17272) );
  DFF_X1 matrix_mul_2D_reg_7__7__20_ ( .D(n886), .CK(clk), .Q(
        matrix_mul_2D_7__7__20_), .QN(n17270) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_1 add_103_I8_I8 ( 
        .A({matrix_mul_2D_7__7__20_, matrix_mul_2D_7__7__19_, 
        matrix_mul_2D_7__7__18_, matrix_mul_2D_7__7__17_, 
        matrix_mul_2D_7__7__16_, matrix_mul_2D_7__7__15_, 
        matrix_mul_2D_7__7__14_, matrix_mul_2D_7__7__13_, 
        matrix_mul_2D_7__7__12_, matrix_mul_2D_7__7__11_, 
        matrix_mul_2D_7__7__10_, matrix_mul_2D_7__7__9_, 
        matrix_mul_2D_7__7__8_, matrix_mul_2D_7__7__7_, matrix_mul_2D_7__7__6_, 
        matrix_mul_2D_7__7__5_, matrix_mul_2D_7__7__4_, matrix_mul_2D_7__7__3_, 
        matrix_mul_2D_7__7__2_, matrix_mul_2D_7__7__1_, n19328}), .B({n872, 
        n870, n873, n872, n871, n870, N7960, N7959, N7958, N7957, N7956, N7955, 
        N7954, N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946}), .SUM(
        {N7999, N7998, N7997, N7996, N7995, N7994, N7993, N7992, N7991, N7990, 
        N7989, N7988, N7987, N7986, N7985, N7984, N7983, N7982, N7981, N7980, 
        N7979}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_2 add_103_I7_I8 ( 
        .A({matrix_mul_2D_7__6__20_, matrix_mul_2D_7__6__19_, 
        matrix_mul_2D_7__6__18_, matrix_mul_2D_7__6__17_, 
        matrix_mul_2D_7__6__16_, matrix_mul_2D_7__6__15_, 
        matrix_mul_2D_7__6__14_, matrix_mul_2D_7__6__13_, 
        matrix_mul_2D_7__6__12_, matrix_mul_2D_7__6__11_, 
        matrix_mul_2D_7__6__10_, matrix_mul_2D_7__6__9_, 
        matrix_mul_2D_7__6__8_, matrix_mul_2D_7__6__7_, matrix_mul_2D_7__6__6_, 
        matrix_mul_2D_7__6__5_, matrix_mul_2D_7__6__4_, matrix_mul_2D_7__6__3_, 
        matrix_mul_2D_7__6__2_, matrix_mul_2D_7__6__1_, n19325}), .B({n867, 
        n865, n868, n867, n866, n865, N7878, N7877, N7876, N7875, N7874, N7873, 
        N7872, N7871, N7870, N7869, N7868, N7867, N7866, N7865, N7864}), .SUM(
        {N7917, N7916, N7915, N7914, N7913, N7912, N7911, N7910, N7909, N7908, 
        N7907, N7906, N7905, N7904, N7903, N7902, N7901, N7900, N7899, N7898, 
        N7897}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_3 add_103_I6_I8 ( 
        .A({matrix_mul_2D_7__5__20_, matrix_mul_2D_7__5__19_, 
        matrix_mul_2D_7__5__18_, matrix_mul_2D_7__5__17_, 
        matrix_mul_2D_7__5__16_, matrix_mul_2D_7__5__15_, 
        matrix_mul_2D_7__5__14_, matrix_mul_2D_7__5__13_, 
        matrix_mul_2D_7__5__12_, matrix_mul_2D_7__5__11_, 
        matrix_mul_2D_7__5__10_, matrix_mul_2D_7__5__9_, 
        matrix_mul_2D_7__5__8_, matrix_mul_2D_7__5__7_, matrix_mul_2D_7__5__6_, 
        matrix_mul_2D_7__5__5_, matrix_mul_2D_7__5__4_, matrix_mul_2D_7__5__3_, 
        matrix_mul_2D_7__5__2_, matrix_mul_2D_7__5__1_, matrix_mul_2D_7__5__0_}), .B({n862, n860, n863, n862, n861, n860, N7789, N7788, N7787, N7786, N7785, 
        N7784, N7783, N7782, N7781, N7780, N7779, N7778, N7777, N7776, N7775}), 
        .SUM({N7828, N7827, N7826, N7825, N7824, N7823, N7822, N7821, N7820, 
        N7819, N7818, N7817, N7816, N7815, N7814, N7813, N7812, N7811, N7810, 
        N7809, N7808}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_4 add_103_I5_I8 ( 
        .A({matrix_mul_2D_7__4__20_, matrix_mul_2D_7__4__19_, 
        matrix_mul_2D_7__4__18_, matrix_mul_2D_7__4__17_, 
        matrix_mul_2D_7__4__16_, matrix_mul_2D_7__4__15_, 
        matrix_mul_2D_7__4__14_, matrix_mul_2D_7__4__13_, 
        matrix_mul_2D_7__4__12_, matrix_mul_2D_7__4__11_, 
        matrix_mul_2D_7__4__10_, matrix_mul_2D_7__4__9_, 
        matrix_mul_2D_7__4__8_, matrix_mul_2D_7__4__7_, matrix_mul_2D_7__4__6_, 
        matrix_mul_2D_7__4__5_, matrix_mul_2D_7__4__4_, matrix_mul_2D_7__4__3_, 
        matrix_mul_2D_7__4__2_, matrix_mul_2D_7__4__1_, matrix_mul_2D_7__4__0_}), .B({n857, n855, n858, n857, n856, n855, N7710, N7709, N7708, N7707, N7706, 
        N7705, N7704, N7703, N7702, N7701, N7700, N7699, N7698, N7697, N7696}), 
        .SUM({N7749, N7748, N7747, N7746, N7745, N7744, N7743, N7742, N7741, 
        N7740, N7739, N7738, N7737, N7736, N7735, N7734, N7733, N7732, N7731, 
        N7730, N7729}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_5 add_103_I4_I8 ( 
        .A({matrix_mul_2D_7__3__20_, matrix_mul_2D_7__3__19_, 
        matrix_mul_2D_7__3__18_, matrix_mul_2D_7__3__17_, 
        matrix_mul_2D_7__3__16_, matrix_mul_2D_7__3__15_, 
        matrix_mul_2D_7__3__14_, matrix_mul_2D_7__3__13_, 
        matrix_mul_2D_7__3__12_, matrix_mul_2D_7__3__11_, 
        matrix_mul_2D_7__3__10_, matrix_mul_2D_7__3__9_, 
        matrix_mul_2D_7__3__8_, matrix_mul_2D_7__3__7_, matrix_mul_2D_7__3__6_, 
        matrix_mul_2D_7__3__5_, matrix_mul_2D_7__3__4_, matrix_mul_2D_7__3__3_, 
        matrix_mul_2D_7__3__2_, matrix_mul_2D_7__3__1_, matrix_mul_2D_7__3__0_}), .B({n852, n850, n853, n852, n851, n850, N7621, N7620, N7619, N7618, N7617, 
        N7616, N7615, N7614, N7613, N7612, N7611, N7610, N7609, N7608, N7607}), 
        .SUM({N7660, N7659, N7658, N7657, N7656, N7655, N7654, N7653, N7652, 
        N7651, N7650, N7649, N7648, N7647, N7646, N7645, N7644, N7643, N7642, 
        N7641, N7640}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_6 add_103_I3_I8 ( 
        .A({matrix_mul_2D_7__2__20_, matrix_mul_2D_7__2__19_, 
        matrix_mul_2D_7__2__18_, matrix_mul_2D_7__2__17_, 
        matrix_mul_2D_7__2__16_, matrix_mul_2D_7__2__15_, 
        matrix_mul_2D_7__2__14_, matrix_mul_2D_7__2__13_, 
        matrix_mul_2D_7__2__12_, matrix_mul_2D_7__2__11_, 
        matrix_mul_2D_7__2__10_, matrix_mul_2D_7__2__9_, 
        matrix_mul_2D_7__2__8_, matrix_mul_2D_7__2__7_, matrix_mul_2D_7__2__6_, 
        matrix_mul_2D_7__2__5_, matrix_mul_2D_7__2__4_, matrix_mul_2D_7__2__3_, 
        matrix_mul_2D_7__2__2_, matrix_mul_2D_7__2__1_, matrix_mul_2D_7__2__0_}), .B({n847, n845, n848, n847, n846, n845, N7542, N7541, N7540, N7539, N7538, 
        N7537, N7536, N7535, N7534, N7533, N7532, N7531, N7530, N7529, N7528}), 
        .SUM({N7581, N7580, N7579, N7578, N7577, N7576, N7575, N7574, N7573, 
        N7572, N7571, N7570, N7569, N7568, N7567, N7566, N7565, N7564, N7563, 
        N7562, N7561}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_7 add_103_I2_I8 ( 
        .A({matrix_mul_2D_7__1__20_, matrix_mul_2D_7__1__19_, 
        matrix_mul_2D_7__1__18_, matrix_mul_2D_7__1__17_, 
        matrix_mul_2D_7__1__16_, matrix_mul_2D_7__1__15_, 
        matrix_mul_2D_7__1__14_, matrix_mul_2D_7__1__13_, 
        matrix_mul_2D_7__1__12_, matrix_mul_2D_7__1__11_, 
        matrix_mul_2D_7__1__10_, matrix_mul_2D_7__1__9_, 
        matrix_mul_2D_7__1__8_, matrix_mul_2D_7__1__7_, matrix_mul_2D_7__1__6_, 
        matrix_mul_2D_7__1__5_, matrix_mul_2D_7__1__4_, matrix_mul_2D_7__1__3_, 
        matrix_mul_2D_7__1__2_, matrix_mul_2D_7__1__1_, n19329}), .B({n842, 
        n840, n843, n842, n841, n840, N7453, N7452, N7451, N7450, N7449, N7448, 
        N7447, N7446, N7445, N7444, N7443, N7442, N7441, N7440, N7439}), .SUM(
        {N7492, N7491, N7490, N7489, N7488, N7487, N7486, N7485, N7484, N7483, 
        N7482, N7481, N7480, N7479, N7478, N7477, N7476, N7475, N7474, N7473, 
        N7472}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_8 add_103_I8 ( 
        .A({matrix_mul_2D_7__0__20_, matrix_mul_2D_7__0__19_, 
        matrix_mul_2D_7__0__18_, matrix_mul_2D_7__0__17_, 
        matrix_mul_2D_7__0__16_, matrix_mul_2D_7__0__15_, 
        matrix_mul_2D_7__0__14_, matrix_mul_2D_7__0__13_, 
        matrix_mul_2D_7__0__12_, matrix_mul_2D_7__0__11_, 
        matrix_mul_2D_7__0__10_, matrix_mul_2D_7__0__9_, 
        matrix_mul_2D_7__0__8_, matrix_mul_2D_7__0__7_, matrix_mul_2D_7__0__6_, 
        matrix_mul_2D_7__0__5_, matrix_mul_2D_7__0__4_, matrix_mul_2D_7__0__3_, 
        matrix_mul_2D_7__0__2_, matrix_mul_2D_7__0__1_, n19330}), .B({n837, 
        n835, n838, n837, n836, n835, N7374, N7373, N7372, N7371, N7370, N7369, 
        N7368, N7367, N7366, N7365, N7364, N7363, N7362, N7361, N7360}), .SUM(
        {N7413, N7412, N7411, N7410, N7409, N7408, N7407, N7406, N7405, N7404, 
        N7403, N7402, N7401, N7400, N7399, N7398, N7397, N7396, N7395, N7394, 
        N7393}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_9 add_103_I8_I7 ( 
        .A({matrix_mul_2D_6__7__20_, matrix_mul_2D_6__7__19_, 
        matrix_mul_2D_6__7__18_, matrix_mul_2D_6__7__17_, 
        matrix_mul_2D_6__7__16_, matrix_mul_2D_6__7__15_, 
        matrix_mul_2D_6__7__14_, matrix_mul_2D_6__7__13_, 
        matrix_mul_2D_6__7__12_, matrix_mul_2D_6__7__11_, 
        matrix_mul_2D_6__7__10_, matrix_mul_2D_6__7__9_, 
        matrix_mul_2D_6__7__8_, matrix_mul_2D_6__7__7_, matrix_mul_2D_6__7__6_, 
        matrix_mul_2D_6__7__5_, matrix_mul_2D_6__7__4_, matrix_mul_2D_6__7__3_, 
        matrix_mul_2D_6__7__2_, matrix_mul_2D_6__7__1_, n19326}), .B({n832, 
        n830, n833, n832, n831, n830, N7285, N7284, N7283, N7282, N7281, N7280, 
        N7279, N7278, N7277, N7276, N7275, N7274, N7273, N7272, N7271}), .SUM(
        {N7324, N7323, N7322, N7321, N7320, N7319, N7318, N7317, N7316, N7315, 
        N7314, N7313, N7312, N7311, N7310, N7309, N7308, N7307, N7306, N7305, 
        N7304}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_10 add_103_I7_I7 ( 
        .A({matrix_mul_2D_6__6__20_, matrix_mul_2D_6__6__19_, 
        matrix_mul_2D_6__6__18_, matrix_mul_2D_6__6__17_, 
        matrix_mul_2D_6__6__16_, matrix_mul_2D_6__6__15_, 
        matrix_mul_2D_6__6__14_, matrix_mul_2D_6__6__13_, 
        matrix_mul_2D_6__6__12_, matrix_mul_2D_6__6__11_, 
        matrix_mul_2D_6__6__10_, matrix_mul_2D_6__6__9_, 
        matrix_mul_2D_6__6__8_, matrix_mul_2D_6__6__7_, matrix_mul_2D_6__6__6_, 
        matrix_mul_2D_6__6__5_, matrix_mul_2D_6__6__4_, matrix_mul_2D_6__6__3_, 
        matrix_mul_2D_6__6__2_, matrix_mul_2D_6__6__1_, matrix_mul_2D_6__6__0_}), .B({n827, n825, n828, n827, n826, n825, N7203, N7202, N7201, N7200, N7199, 
        N7198, N7197, N7196, N7195, N7194, N7193, N7192, N7191, N7190, N7189}), 
        .SUM({N7242, N7241, N7240, N7239, N7238, N7237, N7236, N7235, N7234, 
        N7233, N7232, N7231, N7230, N7229, N7228, N7227, N7226, N7225, N7224, 
        N7223, N7222}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_11 add_103_I6_I7 ( 
        .A({matrix_mul_2D_6__5__20_, matrix_mul_2D_6__5__19_, 
        matrix_mul_2D_6__5__18_, matrix_mul_2D_6__5__17_, 
        matrix_mul_2D_6__5__16_, matrix_mul_2D_6__5__15_, 
        matrix_mul_2D_6__5__14_, matrix_mul_2D_6__5__13_, 
        matrix_mul_2D_6__5__12_, matrix_mul_2D_6__5__11_, 
        matrix_mul_2D_6__5__10_, matrix_mul_2D_6__5__9_, 
        matrix_mul_2D_6__5__8_, matrix_mul_2D_6__5__7_, matrix_mul_2D_6__5__6_, 
        matrix_mul_2D_6__5__5_, matrix_mul_2D_6__5__4_, matrix_mul_2D_6__5__3_, 
        matrix_mul_2D_6__5__2_, matrix_mul_2D_6__5__1_, n19331}), .B({n822, 
        n820, n823, n822, n821, n820, N7111, N7110, N7109, N7108, N7107, N7106, 
        N7105, N7104, N7103, N7102, N7101, N7100, N7099, N7098, N7097}), .SUM(
        {N7150, N7149, N7148, N7147, N7146, N7145, N7144, N7143, N7142, N7141, 
        N7140, N7139, N7138, N7137, N7136, N7135, N7134, N7133, N7132, N7131, 
        N7130}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_12 add_103_I5_I7 ( 
        .A({matrix_mul_2D_6__4__20_, matrix_mul_2D_6__4__19_, 
        matrix_mul_2D_6__4__18_, matrix_mul_2D_6__4__17_, 
        matrix_mul_2D_6__4__16_, matrix_mul_2D_6__4__15_, 
        matrix_mul_2D_6__4__14_, matrix_mul_2D_6__4__13_, 
        matrix_mul_2D_6__4__12_, matrix_mul_2D_6__4__11_, 
        matrix_mul_2D_6__4__10_, matrix_mul_2D_6__4__9_, 
        matrix_mul_2D_6__4__8_, matrix_mul_2D_6__4__7_, matrix_mul_2D_6__4__6_, 
        matrix_mul_2D_6__4__5_, matrix_mul_2D_6__4__4_, matrix_mul_2D_6__4__3_, 
        matrix_mul_2D_6__4__2_, matrix_mul_2D_6__4__1_, matrix_mul_2D_6__4__0_}), .B({n817, n815, n818, n817, n816, n815, N7029, N7028, N7027, N7026, N7025, 
        N7024, N7023, N7022, N7021, N7020, N7019, N7018, N7017, N7016, N7015}), 
        .SUM({N7068, N7067, N7066, N7065, N7064, N7063, N7062, N7061, N7060, 
        N7059, N7058, N7057, N7056, N7055, N7054, N7053, N7052, N7051, N7050, 
        N7049, N7048}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_13 add_103_I4_I7 ( 
        .A({matrix_mul_2D_6__3__20_, matrix_mul_2D_6__3__19_, 
        matrix_mul_2D_6__3__18_, matrix_mul_2D_6__3__17_, 
        matrix_mul_2D_6__3__16_, matrix_mul_2D_6__3__15_, 
        matrix_mul_2D_6__3__14_, matrix_mul_2D_6__3__13_, 
        matrix_mul_2D_6__3__12_, matrix_mul_2D_6__3__11_, 
        matrix_mul_2D_6__3__10_, matrix_mul_2D_6__3__9_, 
        matrix_mul_2D_6__3__8_, matrix_mul_2D_6__3__7_, matrix_mul_2D_6__3__6_, 
        matrix_mul_2D_6__3__5_, matrix_mul_2D_6__3__4_, matrix_mul_2D_6__3__3_, 
        matrix_mul_2D_6__3__2_, matrix_mul_2D_6__3__1_, matrix_mul_2D_6__3__0_}), .B({n812, n810, n813, n812, n811, n810, N6937, N6936, N6935, N6934, N6933, 
        N6932, N6931, N6930, N6929, N6928, N6927, N6926, N6925, N6924, N6923}), 
        .SUM({N6976, N6975, N6974, N6973, N6972, N6971, N6970, N6969, N6968, 
        N6967, N6966, N6965, N6964, N6963, N6962, N6961, N6960, N6959, N6958, 
        N6957, N6956}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_14 add_103_I3_I7 ( 
        .A({matrix_mul_2D_6__2__20_, matrix_mul_2D_6__2__19_, 
        matrix_mul_2D_6__2__18_, matrix_mul_2D_6__2__17_, 
        matrix_mul_2D_6__2__16_, matrix_mul_2D_6__2__15_, 
        matrix_mul_2D_6__2__14_, matrix_mul_2D_6__2__13_, 
        matrix_mul_2D_6__2__12_, matrix_mul_2D_6__2__11_, 
        matrix_mul_2D_6__2__10_, matrix_mul_2D_6__2__9_, 
        matrix_mul_2D_6__2__8_, matrix_mul_2D_6__2__7_, matrix_mul_2D_6__2__6_, 
        matrix_mul_2D_6__2__5_, matrix_mul_2D_6__2__4_, matrix_mul_2D_6__2__3_, 
        matrix_mul_2D_6__2__2_, matrix_mul_2D_6__2__1_, matrix_mul_2D_6__2__0_}), .B({n807, n805, n808, n807, n806, n805, N6855, N6854, N6853, N6852, N6851, 
        N6850, N6849, N6848, N6847, N6846, N6845, N6844, N6843, N6842, N6841}), 
        .SUM({N6894, N6893, N6892, N6891, N6890, N6889, N6888, N6887, N6886, 
        N6885, N6884, N6883, N6882, N6881, N6880, N6879, N6878, N6877, N6876, 
        N6875, N6874}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_15 add_103_I2_I7 ( 
        .A({matrix_mul_2D_6__1__20_, matrix_mul_2D_6__1__19_, 
        matrix_mul_2D_6__1__18_, matrix_mul_2D_6__1__17_, 
        matrix_mul_2D_6__1__16_, matrix_mul_2D_6__1__15_, 
        matrix_mul_2D_6__1__14_, matrix_mul_2D_6__1__13_, 
        matrix_mul_2D_6__1__12_, matrix_mul_2D_6__1__11_, 
        matrix_mul_2D_6__1__10_, matrix_mul_2D_6__1__9_, 
        matrix_mul_2D_6__1__8_, matrix_mul_2D_6__1__7_, matrix_mul_2D_6__1__6_, 
        matrix_mul_2D_6__1__5_, matrix_mul_2D_6__1__4_, matrix_mul_2D_6__1__3_, 
        matrix_mul_2D_6__1__2_, matrix_mul_2D_6__1__1_, n19332}), .B({n802, 
        n800, n803, n802, n801, n800, N6763, N6762, N6761, N6760, N6759, N6758, 
        N6757, N6756, N6755, N6754, N6753, N6752, N6751, N6750, N6749}), .SUM(
        {N6802, N6801, N6800, N6799, N6798, N6797, N6796, N6795, N6794, N6793, 
        N6792, N6791, N6790, N6789, N6788, N6787, N6786, N6785, N6784, N6783, 
        N6782}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_16 add_103_I7 ( 
        .A({matrix_mul_2D_6__0__20_, matrix_mul_2D_6__0__19_, 
        matrix_mul_2D_6__0__18_, matrix_mul_2D_6__0__17_, 
        matrix_mul_2D_6__0__16_, matrix_mul_2D_6__0__15_, 
        matrix_mul_2D_6__0__14_, matrix_mul_2D_6__0__13_, 
        matrix_mul_2D_6__0__12_, matrix_mul_2D_6__0__11_, 
        matrix_mul_2D_6__0__10_, matrix_mul_2D_6__0__9_, 
        matrix_mul_2D_6__0__8_, matrix_mul_2D_6__0__7_, matrix_mul_2D_6__0__6_, 
        matrix_mul_2D_6__0__5_, matrix_mul_2D_6__0__4_, matrix_mul_2D_6__0__3_, 
        matrix_mul_2D_6__0__2_, matrix_mul_2D_6__0__1_, n19333}), .B({n797, 
        n795, n798, n797, n796, n795, N6681, N6680, N6679, N6678, N6677, N6676, 
        N6675, N6674, N6673, N6672, N6671, N6670, N6669, N6668, N6667}), .SUM(
        {N6720, N6719, N6718, N6717, N6716, N6715, N6714, N6713, N6712, N6711, 
        N6710, N6709, N6708, N6707, N6706, N6705, N6704, N6703, N6702, N6701, 
        N6700}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_17 add_103_I8_I6 ( 
        .A({matrix_mul_2D_5__7__20_, matrix_mul_2D_5__7__19_, 
        matrix_mul_2D_5__7__18_, matrix_mul_2D_5__7__17_, 
        matrix_mul_2D_5__7__16_, matrix_mul_2D_5__7__15_, 
        matrix_mul_2D_5__7__14_, matrix_mul_2D_5__7__13_, 
        matrix_mul_2D_5__7__12_, matrix_mul_2D_5__7__11_, 
        matrix_mul_2D_5__7__10_, matrix_mul_2D_5__7__9_, 
        matrix_mul_2D_5__7__8_, matrix_mul_2D_5__7__7_, matrix_mul_2D_5__7__6_, 
        matrix_mul_2D_5__7__5_, matrix_mul_2D_5__7__4_, matrix_mul_2D_5__7__3_, 
        matrix_mul_2D_5__7__2_, matrix_mul_2D_5__7__1_, n19334}), .B({n792, 
        n790, n793, n792, n791, n790, N6581, N6580, N6579, N6578, N6577, N6576, 
        N6575, N6574, N6573, N6572, N6571, N6570, N6569, N6568, N6567}), .SUM(
        {N6620, N6619, N6618, N6617, N6616, N6615, N6614, N6613, N6612, N6611, 
        N6610, N6609, N6608, N6607, N6606, N6605, N6604, N6603, N6602, N6601, 
        N6600}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_18 add_103_I7_I6 ( 
        .A({matrix_mul_2D_5__6__20_, matrix_mul_2D_5__6__19_, 
        matrix_mul_2D_5__6__18_, matrix_mul_2D_5__6__17_, 
        matrix_mul_2D_5__6__16_, matrix_mul_2D_5__6__15_, 
        matrix_mul_2D_5__6__14_, matrix_mul_2D_5__6__13_, 
        matrix_mul_2D_5__6__12_, matrix_mul_2D_5__6__11_, 
        matrix_mul_2D_5__6__10_, matrix_mul_2D_5__6__9_, 
        matrix_mul_2D_5__6__8_, matrix_mul_2D_5__6__7_, matrix_mul_2D_5__6__6_, 
        matrix_mul_2D_5__6__5_, matrix_mul_2D_5__6__4_, matrix_mul_2D_5__6__3_, 
        matrix_mul_2D_5__6__2_, matrix_mul_2D_5__6__1_, n19335}), .B({n787, 
        n785, n788, n787, n786, n785, N6499, N6498, N6497, N6496, N6495, N6494, 
        N6493, N6492, N6491, N6490, N6489, N6488, N6487, N6486, N6485}), .SUM(
        {N6538, N6537, N6536, N6535, N6534, N6533, N6532, N6531, N6530, N6529, 
        N6528, N6527, N6526, N6525, N6524, N6523, N6522, N6521, N6520, N6519, 
        N6518}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_19 add_103_I6_I6 ( 
        .A({matrix_mul_2D_5__5__20_, matrix_mul_2D_5__5__19_, 
        matrix_mul_2D_5__5__18_, matrix_mul_2D_5__5__17_, 
        matrix_mul_2D_5__5__16_, matrix_mul_2D_5__5__15_, 
        matrix_mul_2D_5__5__14_, matrix_mul_2D_5__5__13_, 
        matrix_mul_2D_5__5__12_, matrix_mul_2D_5__5__11_, 
        matrix_mul_2D_5__5__10_, matrix_mul_2D_5__5__9_, 
        matrix_mul_2D_5__5__8_, matrix_mul_2D_5__5__7_, matrix_mul_2D_5__5__6_, 
        matrix_mul_2D_5__5__5_, matrix_mul_2D_5__5__4_, matrix_mul_2D_5__5__3_, 
        matrix_mul_2D_5__5__2_, matrix_mul_2D_5__5__1_, matrix_mul_2D_5__5__0_}), .B({n782, n780, n783, n782, n781, n780, N6410, N6409, N6408, N6407, N6406, 
        N6405, N6404, N6403, N6402, N6401, N6400, N6399, N6398, N6397, N6396}), 
        .SUM({N6449, N6448, N6447, N6446, N6445, N6444, N6443, N6442, N6441, 
        N6440, N6439, N6438, N6437, N6436, N6435, N6434, N6433, N6432, N6431, 
        N6430, N6429}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_20 add_103_I5_I6 ( 
        .A({matrix_mul_2D_5__4__20_, matrix_mul_2D_5__4__19_, 
        matrix_mul_2D_5__4__18_, matrix_mul_2D_5__4__17_, 
        matrix_mul_2D_5__4__16_, matrix_mul_2D_5__4__15_, 
        matrix_mul_2D_5__4__14_, matrix_mul_2D_5__4__13_, 
        matrix_mul_2D_5__4__12_, matrix_mul_2D_5__4__11_, 
        matrix_mul_2D_5__4__10_, matrix_mul_2D_5__4__9_, 
        matrix_mul_2D_5__4__8_, matrix_mul_2D_5__4__7_, matrix_mul_2D_5__4__6_, 
        matrix_mul_2D_5__4__5_, matrix_mul_2D_5__4__4_, matrix_mul_2D_5__4__3_, 
        matrix_mul_2D_5__4__2_, matrix_mul_2D_5__4__1_, matrix_mul_2D_5__4__0_}), .B({n777, n775, n778, n777, n776, n775, N6331, N6330, N6329, N6328, N6327, 
        N6326, N6325, N6324, N6323, N6322, N6321, N6320, N6319, N6318, N6317}), 
        .SUM({N6370, N6369, N6368, N6367, N6366, N6365, N6364, N6363, N6362, 
        N6361, N6360, N6359, N6358, N6357, N6356, N6355, N6354, N6353, N6352, 
        N6351, N6350}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_21 add_103_I4_I6 ( 
        .A({matrix_mul_2D_5__3__20_, matrix_mul_2D_5__3__19_, 
        matrix_mul_2D_5__3__18_, matrix_mul_2D_5__3__17_, 
        matrix_mul_2D_5__3__16_, matrix_mul_2D_5__3__15_, 
        matrix_mul_2D_5__3__14_, matrix_mul_2D_5__3__13_, 
        matrix_mul_2D_5__3__12_, matrix_mul_2D_5__3__11_, 
        matrix_mul_2D_5__3__10_, matrix_mul_2D_5__3__9_, 
        matrix_mul_2D_5__3__8_, matrix_mul_2D_5__3__7_, matrix_mul_2D_5__3__6_, 
        matrix_mul_2D_5__3__5_, matrix_mul_2D_5__3__4_, matrix_mul_2D_5__3__3_, 
        matrix_mul_2D_5__3__2_, matrix_mul_2D_5__3__1_, n19336}), .B({n772, 
        n770, n773, n772, n771, n770, N6242, N6241, N6240, N6239, N6238, N6237, 
        N6236, N6235, N6234, N6233, N6232, N6231, N6230, N6229, N6228}), .SUM(
        {N6281, N6280, N6279, N6278, N6277, N6276, N6275, N6274, N6273, N6272, 
        N6271, N6270, N6269, N6268, N6267, N6266, N6265, N6264, N6263, N6262, 
        N6261}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_22 add_103_I3_I6 ( 
        .A({matrix_mul_2D_5__2__20_, matrix_mul_2D_5__2__19_, 
        matrix_mul_2D_5__2__18_, matrix_mul_2D_5__2__17_, 
        matrix_mul_2D_5__2__16_, matrix_mul_2D_5__2__15_, 
        matrix_mul_2D_5__2__14_, matrix_mul_2D_5__2__13_, 
        matrix_mul_2D_5__2__12_, matrix_mul_2D_5__2__11_, 
        matrix_mul_2D_5__2__10_, matrix_mul_2D_5__2__9_, 
        matrix_mul_2D_5__2__8_, matrix_mul_2D_5__2__7_, matrix_mul_2D_5__2__6_, 
        matrix_mul_2D_5__2__5_, matrix_mul_2D_5__2__4_, matrix_mul_2D_5__2__3_, 
        matrix_mul_2D_5__2__2_, matrix_mul_2D_5__2__1_, n19337}), .B({n767, 
        n765, n768, n767, n766, n765, N6163, N6162, N6161, N6160, N6159, N6158, 
        N6157, N6156, N6155, N6154, N6153, N6152, N6151, N6150, N6149}), .SUM(
        {N6202, N6201, N6200, N6199, N6198, N6197, N6196, N6195, N6194, N6193, 
        N6192, N6191, N6190, N6189, N6188, N6187, N6186, N6185, N6184, N6183, 
        N6182}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_23 add_103_I2_I6 ( 
        .A({matrix_mul_2D_5__1__20_, matrix_mul_2D_5__1__19_, 
        matrix_mul_2D_5__1__18_, matrix_mul_2D_5__1__17_, 
        matrix_mul_2D_5__1__16_, matrix_mul_2D_5__1__15_, 
        matrix_mul_2D_5__1__14_, matrix_mul_2D_5__1__13_, 
        matrix_mul_2D_5__1__12_, matrix_mul_2D_5__1__11_, 
        matrix_mul_2D_5__1__10_, matrix_mul_2D_5__1__9_, 
        matrix_mul_2D_5__1__8_, matrix_mul_2D_5__1__7_, matrix_mul_2D_5__1__6_, 
        matrix_mul_2D_5__1__5_, matrix_mul_2D_5__1__4_, matrix_mul_2D_5__1__3_, 
        matrix_mul_2D_5__1__2_, matrix_mul_2D_5__1__1_, n19338}), .B({n762, 
        n760, n763, n762, n761, n760, N6074, N6073, N6072, N6071, N6070, N6069, 
        N6068, N6067, N6066, N6065, N6064, N6063, N6062, N6061, N6060}), .SUM(
        {N6113, N6112, N6111, N6110, N6109, N6108, N6107, N6106, N6105, N6104, 
        N6103, N6102, N6101, N6100, N6099, N6098, N6097, N6096, N6095, N6094, 
        N6093}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_24 add_103_I6 ( 
        .A({matrix_mul_2D_5__0__20_, matrix_mul_2D_5__0__19_, 
        matrix_mul_2D_5__0__18_, matrix_mul_2D_5__0__17_, 
        matrix_mul_2D_5__0__16_, matrix_mul_2D_5__0__15_, 
        matrix_mul_2D_5__0__14_, matrix_mul_2D_5__0__13_, 
        matrix_mul_2D_5__0__12_, matrix_mul_2D_5__0__11_, 
        matrix_mul_2D_5__0__10_, matrix_mul_2D_5__0__9_, 
        matrix_mul_2D_5__0__8_, matrix_mul_2D_5__0__7_, matrix_mul_2D_5__0__6_, 
        matrix_mul_2D_5__0__5_, matrix_mul_2D_5__0__4_, matrix_mul_2D_5__0__3_, 
        matrix_mul_2D_5__0__2_, matrix_mul_2D_5__0__1_, n19339}), .B({n757, 
        n755, n758, n757, n756, n755, N5995, N5994, N5993, N5992, N5991, N5990, 
        N5989, N5988, N5987, N5986, N5985, N5984, N5983, N5982, N5981}), .SUM(
        {N6034, N6033, N6032, N6031, N6030, N6029, N6028, N6027, N6026, N6025, 
        N6024, N6023, N6022, N6021, N6020, N6019, N6018, N6017, N6016, N6015, 
        N6014}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_25 add_103_I8_I5 ( 
        .A({matrix_mul_2D_4__7__20_, matrix_mul_2D_4__7__19_, 
        matrix_mul_2D_4__7__18_, matrix_mul_2D_4__7__17_, 
        matrix_mul_2D_4__7__16_, matrix_mul_2D_4__7__15_, 
        matrix_mul_2D_4__7__14_, matrix_mul_2D_4__7__13_, 
        matrix_mul_2D_4__7__12_, matrix_mul_2D_4__7__11_, 
        matrix_mul_2D_4__7__10_, matrix_mul_2D_4__7__9_, 
        matrix_mul_2D_4__7__8_, matrix_mul_2D_4__7__7_, matrix_mul_2D_4__7__6_, 
        matrix_mul_2D_4__7__5_, matrix_mul_2D_4__7__4_, matrix_mul_2D_4__7__3_, 
        matrix_mul_2D_4__7__2_, matrix_mul_2D_4__7__1_, n19340}), .B({n752, 
        n750, n753, n752, n751, n750, N5906, N5905, N5904, N5903, N5902, N5901, 
        N5900, N5899, N5898, N5897, N5896, N5895, N5894, N5893, N5892}), .SUM(
        {N5945, N5944, N5943, N5942, N5941, N5940, N5939, N5938, N5937, N5936, 
        N5935, N5934, N5933, N5932, N5931, N5930, N5929, N5928, N5927, N5926, 
        N5925}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_26 add_103_I7_I5 ( 
        .A({matrix_mul_2D_4__6__20_, matrix_mul_2D_4__6__19_, 
        matrix_mul_2D_4__6__18_, matrix_mul_2D_4__6__17_, 
        matrix_mul_2D_4__6__16_, matrix_mul_2D_4__6__15_, 
        matrix_mul_2D_4__6__14_, matrix_mul_2D_4__6__13_, 
        matrix_mul_2D_4__6__12_, matrix_mul_2D_4__6__11_, 
        matrix_mul_2D_4__6__10_, matrix_mul_2D_4__6__9_, 
        matrix_mul_2D_4__6__8_, matrix_mul_2D_4__6__7_, matrix_mul_2D_4__6__6_, 
        matrix_mul_2D_4__6__5_, matrix_mul_2D_4__6__4_, matrix_mul_2D_4__6__3_, 
        matrix_mul_2D_4__6__2_, matrix_mul_2D_4__6__1_, n19341}), .B({n747, 
        n745, n748, n747, n746, n745, N5824, N5823, N5822, N5821, N5820, N5819, 
        N5818, N5817, N5816, N5815, N5814, N5813, N5812, N5811, N5810}), .SUM(
        {N5863, N5862, N5861, N5860, N5859, N5858, N5857, N5856, N5855, N5854, 
        N5853, N5852, N5851, N5850, N5849, N5848, N5847, N5846, N5845, N5844, 
        N5843}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_27 add_103_I6_I5 ( 
        .A({matrix_mul_2D_4__5__20_, matrix_mul_2D_4__5__19_, 
        matrix_mul_2D_4__5__18_, matrix_mul_2D_4__5__17_, 
        matrix_mul_2D_4__5__16_, matrix_mul_2D_4__5__15_, 
        matrix_mul_2D_4__5__14_, matrix_mul_2D_4__5__13_, 
        matrix_mul_2D_4__5__12_, matrix_mul_2D_4__5__11_, 
        matrix_mul_2D_4__5__10_, matrix_mul_2D_4__5__9_, 
        matrix_mul_2D_4__5__8_, matrix_mul_2D_4__5__7_, matrix_mul_2D_4__5__6_, 
        matrix_mul_2D_4__5__5_, matrix_mul_2D_4__5__4_, matrix_mul_2D_4__5__3_, 
        matrix_mul_2D_4__5__2_, matrix_mul_2D_4__5__1_, matrix_mul_2D_4__5__0_}), .B({n742, n740, n743, n742, n741, n740, N5735, N5734, N5733, N5732, N5731, 
        N5730, N5729, N5728, N5727, N5726, N5725, N5724, N5723, N5722, N5721}), 
        .SUM({N5774, N5773, N5772, N5771, N5770, N5769, N5768, N5767, N5766, 
        N5765, N5764, N5763, N5762, N5761, N5760, N5759, N5758, N5757, N5756, 
        N5755, N5754}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_28 add_103_I5_I5 ( 
        .A({matrix_mul_2D_4__4__20_, matrix_mul_2D_4__4__19_, 
        matrix_mul_2D_4__4__18_, matrix_mul_2D_4__4__17_, 
        matrix_mul_2D_4__4__16_, matrix_mul_2D_4__4__15_, 
        matrix_mul_2D_4__4__14_, matrix_mul_2D_4__4__13_, 
        matrix_mul_2D_4__4__12_, matrix_mul_2D_4__4__11_, 
        matrix_mul_2D_4__4__10_, matrix_mul_2D_4__4__9_, 
        matrix_mul_2D_4__4__8_, matrix_mul_2D_4__4__7_, matrix_mul_2D_4__4__6_, 
        matrix_mul_2D_4__4__5_, matrix_mul_2D_4__4__4_, matrix_mul_2D_4__4__3_, 
        matrix_mul_2D_4__4__2_, matrix_mul_2D_4__4__1_, matrix_mul_2D_4__4__0_}), .B({n737, n735, n738, n737, n736, n735, N5656, N5655, N5654, N5653, N5652, 
        N5651, N5650, N5649, N5648, N5647, N5646, N5645, N5644, N5643, N5642}), 
        .SUM({N5695, N5694, N5693, N5692, N5691, N5690, N5689, N5688, N5687, 
        N5686, N5685, N5684, N5683, N5682, N5681, N5680, N5679, N5678, N5677, 
        N5676, N5675}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_29 add_103_I4_I5 ( 
        .A({matrix_mul_2D_4__3__20_, matrix_mul_2D_4__3__19_, 
        matrix_mul_2D_4__3__18_, matrix_mul_2D_4__3__17_, 
        matrix_mul_2D_4__3__16_, matrix_mul_2D_4__3__15_, 
        matrix_mul_2D_4__3__14_, matrix_mul_2D_4__3__13_, 
        matrix_mul_2D_4__3__12_, matrix_mul_2D_4__3__11_, 
        matrix_mul_2D_4__3__10_, matrix_mul_2D_4__3__9_, 
        matrix_mul_2D_4__3__8_, matrix_mul_2D_4__3__7_, matrix_mul_2D_4__3__6_, 
        matrix_mul_2D_4__3__5_, matrix_mul_2D_4__3__4_, matrix_mul_2D_4__3__3_, 
        matrix_mul_2D_4__3__2_, matrix_mul_2D_4__3__1_, n19342}), .B({n732, 
        n730, n733, n732, n731, n730, N5567, N5566, N5565, N5564, N5563, N5562, 
        N5561, N5560, N5559, N5558, N5557, N5556, N5555, N5554, N5553}), .SUM(
        {N5606, N5605, N5604, N5603, N5602, N5601, N5600, N5599, N5598, N5597, 
        N5596, N5595, N5594, N5593, N5592, N5591, N5590, N5589, N5588, N5587, 
        N5586}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_30 add_103_I3_I5 ( 
        .A({matrix_mul_2D_4__2__20_, matrix_mul_2D_4__2__19_, 
        matrix_mul_2D_4__2__18_, matrix_mul_2D_4__2__17_, 
        matrix_mul_2D_4__2__16_, matrix_mul_2D_4__2__15_, 
        matrix_mul_2D_4__2__14_, matrix_mul_2D_4__2__13_, 
        matrix_mul_2D_4__2__12_, matrix_mul_2D_4__2__11_, 
        matrix_mul_2D_4__2__10_, matrix_mul_2D_4__2__9_, 
        matrix_mul_2D_4__2__8_, matrix_mul_2D_4__2__7_, matrix_mul_2D_4__2__6_, 
        matrix_mul_2D_4__2__5_, matrix_mul_2D_4__2__4_, matrix_mul_2D_4__2__3_, 
        matrix_mul_2D_4__2__2_, matrix_mul_2D_4__2__1_, n19343}), .B({n727, 
        n725, n728, n727, n726, n725, N5488, N5487, N5486, N5485, N5484, N5483, 
        N5482, N5481, N5480, N5479, N5478, N5477, N5476, N5475, N5474}), .SUM(
        {N5527, N5526, N5525, N5524, N5523, N5522, N5521, N5520, N5519, N5518, 
        N5517, N5516, N5515, N5514, N5513, N5512, N5511, N5510, N5509, N5508, 
        N5507}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_31 add_103_I2_I5 ( 
        .A({matrix_mul_2D_4__1__20_, matrix_mul_2D_4__1__19_, 
        matrix_mul_2D_4__1__18_, matrix_mul_2D_4__1__17_, 
        matrix_mul_2D_4__1__16_, matrix_mul_2D_4__1__15_, 
        matrix_mul_2D_4__1__14_, matrix_mul_2D_4__1__13_, 
        matrix_mul_2D_4__1__12_, matrix_mul_2D_4__1__11_, 
        matrix_mul_2D_4__1__10_, matrix_mul_2D_4__1__9_, 
        matrix_mul_2D_4__1__8_, matrix_mul_2D_4__1__7_, matrix_mul_2D_4__1__6_, 
        matrix_mul_2D_4__1__5_, matrix_mul_2D_4__1__4_, matrix_mul_2D_4__1__3_, 
        matrix_mul_2D_4__1__2_, matrix_mul_2D_4__1__1_, n19344}), .B({n722, 
        n720, n723, n722, n721, n720, N5399, N5398, N5397, N5396, N5395, N5394, 
        N5393, N5392, N5391, N5390, N5389, N5388, N5387, N5386, N5385}), .SUM(
        {N5438, N5437, N5436, N5435, N5434, N5433, N5432, N5431, N5430, N5429, 
        N5428, N5427, N5426, N5425, N5424, N5423, N5422, N5421, N5420, N5419, 
        N5418}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_32 add_103_I5 ( 
        .A({matrix_mul_2D_4__0__20_, matrix_mul_2D_4__0__19_, 
        matrix_mul_2D_4__0__18_, matrix_mul_2D_4__0__17_, 
        matrix_mul_2D_4__0__16_, matrix_mul_2D_4__0__15_, 
        matrix_mul_2D_4__0__14_, matrix_mul_2D_4__0__13_, 
        matrix_mul_2D_4__0__12_, matrix_mul_2D_4__0__11_, 
        matrix_mul_2D_4__0__10_, matrix_mul_2D_4__0__9_, 
        matrix_mul_2D_4__0__8_, matrix_mul_2D_4__0__7_, matrix_mul_2D_4__0__6_, 
        matrix_mul_2D_4__0__5_, matrix_mul_2D_4__0__4_, matrix_mul_2D_4__0__3_, 
        matrix_mul_2D_4__0__2_, matrix_mul_2D_4__0__1_, n19345}), .B({n717, 
        n715, n718, n717, n716, n715, N5320, N5319, N5318, N5317, N5316, N5315, 
        N5314, N5313, N5312, N5311, N5310, N5309, N5308, N5307, N5306}), .SUM(
        {N5359, N5358, N5357, N5356, N5355, N5354, N5353, N5352, N5351, N5350, 
        N5349, N5348, N5347, N5346, N5345, N5344, N5343, N5342, N5341, N5340, 
        N5339}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_33 add_103_I8_I4 ( 
        .A({matrix_mul_2D_3__7__20_, matrix_mul_2D_3__7__19_, 
        matrix_mul_2D_3__7__18_, matrix_mul_2D_3__7__17_, 
        matrix_mul_2D_3__7__16_, matrix_mul_2D_3__7__15_, 
        matrix_mul_2D_3__7__14_, matrix_mul_2D_3__7__13_, 
        matrix_mul_2D_3__7__12_, matrix_mul_2D_3__7__11_, 
        matrix_mul_2D_3__7__10_, matrix_mul_2D_3__7__9_, 
        matrix_mul_2D_3__7__8_, matrix_mul_2D_3__7__7_, matrix_mul_2D_3__7__6_, 
        matrix_mul_2D_3__7__5_, matrix_mul_2D_3__7__4_, matrix_mul_2D_3__7__3_, 
        matrix_mul_2D_3__7__2_, matrix_mul_2D_3__7__1_, n19346}), .B({n712, 
        n710, n713, n712, n711, n710, N5231, N5230, N5229, N5228, N5227, N5226, 
        N5225, N5224, N5223, N5222, N5221, N5220, N5219, N5218, N5217}), .SUM(
        {N5270, N5269, N5268, N5267, N5266, N5265, N5264, N5263, N5262, N5261, 
        N5260, N5259, N5258, N5257, N5256, N5255, N5254, N5253, N5252, N5251, 
        N5250}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_34 add_103_I7_I4 ( 
        .A({matrix_mul_2D_3__6__20_, matrix_mul_2D_3__6__19_, 
        matrix_mul_2D_3__6__18_, matrix_mul_2D_3__6__17_, 
        matrix_mul_2D_3__6__16_, matrix_mul_2D_3__6__15_, 
        matrix_mul_2D_3__6__14_, matrix_mul_2D_3__6__13_, 
        matrix_mul_2D_3__6__12_, matrix_mul_2D_3__6__11_, 
        matrix_mul_2D_3__6__10_, matrix_mul_2D_3__6__9_, 
        matrix_mul_2D_3__6__8_, matrix_mul_2D_3__6__7_, matrix_mul_2D_3__6__6_, 
        matrix_mul_2D_3__6__5_, matrix_mul_2D_3__6__4_, matrix_mul_2D_3__6__3_, 
        matrix_mul_2D_3__6__2_, matrix_mul_2D_3__6__1_, n19347}), .B({n707, 
        n705, n708, n707, n706, n705, N5149, N5148, N5147, N5146, N5145, N5144, 
        N5143, N5142, N5141, N5140, N5139, N5138, N5137, N5136, N5135}), .SUM(
        {N5188, N5187, N5186, N5185, N5184, N5183, N5182, N5181, N5180, N5179, 
        N5178, N5177, N5176, N5175, N5174, N5173, N5172, N5171, N5170, N5169, 
        N5168}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_35 add_103_I6_I4 ( 
        .A({matrix_mul_2D_3__5__20_, matrix_mul_2D_3__5__19_, 
        matrix_mul_2D_3__5__18_, matrix_mul_2D_3__5__17_, 
        matrix_mul_2D_3__5__16_, matrix_mul_2D_3__5__15_, 
        matrix_mul_2D_3__5__14_, matrix_mul_2D_3__5__13_, 
        matrix_mul_2D_3__5__12_, matrix_mul_2D_3__5__11_, 
        matrix_mul_2D_3__5__10_, matrix_mul_2D_3__5__9_, 
        matrix_mul_2D_3__5__8_, matrix_mul_2D_3__5__7_, matrix_mul_2D_3__5__6_, 
        matrix_mul_2D_3__5__5_, matrix_mul_2D_3__5__4_, matrix_mul_2D_3__5__3_, 
        matrix_mul_2D_3__5__2_, matrix_mul_2D_3__5__1_, n19348}), .B({n702, 
        n700, n703, n702, n701, n700, N5057, N5056, N5055, N5054, N5053, N5052, 
        N5051, N5050, N5049, N5048, N5047, N5046, N5045, N5044, N5043}), .SUM(
        {N5096, N5095, N5094, N5093, N5092, N5091, N5090, N5089, N5088, N5087, 
        N5086, N5085, N5084, N5083, N5082, N5081, N5080, N5079, N5078, N5077, 
        N5076}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_36 add_103_I5_I4 ( 
        .A({matrix_mul_2D_3__4__20_, matrix_mul_2D_3__4__19_, 
        matrix_mul_2D_3__4__18_, matrix_mul_2D_3__4__17_, 
        matrix_mul_2D_3__4__16_, matrix_mul_2D_3__4__15_, 
        matrix_mul_2D_3__4__14_, matrix_mul_2D_3__4__13_, 
        matrix_mul_2D_3__4__12_, matrix_mul_2D_3__4__11_, 
        matrix_mul_2D_3__4__10_, matrix_mul_2D_3__4__9_, 
        matrix_mul_2D_3__4__8_, matrix_mul_2D_3__4__7_, matrix_mul_2D_3__4__6_, 
        matrix_mul_2D_3__4__5_, matrix_mul_2D_3__4__4_, matrix_mul_2D_3__4__3_, 
        matrix_mul_2D_3__4__2_, matrix_mul_2D_3__4__1_, matrix_mul_2D_3__4__0_}), .B({n697, n695, n698, n697, n696, n695, N4975, N4974, N4973, N4972, N4971, 
        N4970, N4969, N4968, N4967, N4966, N4965, N4964, N4963, N4962, N4961}), 
        .SUM({N5014, N5013, N5012, N5011, N5010, N5009, N5008, N5007, N5006, 
        N5005, N5004, N5003, N5002, N5001, N5000, N4999, N4998, N4997, N4996, 
        N4995, N4994}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_37 add_103_I4_I4 ( 
        .A({matrix_mul_2D_3__3__20_, matrix_mul_2D_3__3__19_, 
        matrix_mul_2D_3__3__18_, matrix_mul_2D_3__3__17_, 
        matrix_mul_2D_3__3__16_, matrix_mul_2D_3__3__15_, 
        matrix_mul_2D_3__3__14_, matrix_mul_2D_3__3__13_, 
        matrix_mul_2D_3__3__12_, matrix_mul_2D_3__3__11_, 
        matrix_mul_2D_3__3__10_, matrix_mul_2D_3__3__9_, 
        matrix_mul_2D_3__3__8_, matrix_mul_2D_3__3__7_, matrix_mul_2D_3__3__6_, 
        matrix_mul_2D_3__3__5_, matrix_mul_2D_3__3__4_, matrix_mul_2D_3__3__3_, 
        matrix_mul_2D_3__3__2_, matrix_mul_2D_3__3__1_, matrix_mul_2D_3__3__0_}), .B({n692, n690, n693, n692, n691, n690, N4883, N4882, N4881, N4880, N4879, 
        N4878, N4877, N4876, N4875, N4874, N4873, N4872, N4871, N4870, N4869}), 
        .SUM({N4922, N4921, N4920, N4919, N4918, N4917, N4916, N4915, N4914, 
        N4913, N4912, N4911, N4910, N4909, N4908, N4907, N4906, N4905, N4904, 
        N4903, N4902}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_38 add_103_I3_I4 ( 
        .A({matrix_mul_2D_3__2__20_, matrix_mul_2D_3__2__19_, 
        matrix_mul_2D_3__2__18_, matrix_mul_2D_3__2__17_, 
        matrix_mul_2D_3__2__16_, matrix_mul_2D_3__2__15_, 
        matrix_mul_2D_3__2__14_, matrix_mul_2D_3__2__13_, 
        matrix_mul_2D_3__2__12_, matrix_mul_2D_3__2__11_, 
        matrix_mul_2D_3__2__10_, matrix_mul_2D_3__2__9_, 
        matrix_mul_2D_3__2__8_, matrix_mul_2D_3__2__7_, matrix_mul_2D_3__2__6_, 
        matrix_mul_2D_3__2__5_, matrix_mul_2D_3__2__4_, matrix_mul_2D_3__2__3_, 
        matrix_mul_2D_3__2__2_, matrix_mul_2D_3__2__1_, n19349}), .B({n687, 
        n685, n688, n687, n686, n685, N4801, N4800, N4799, N4798, N4797, N4796, 
        N4795, N4794, N4793, N4792, N4791, N4790, N4789, N4788, N4787}), .SUM(
        {N4840, N4839, N4838, N4837, N4836, N4835, N4834, N4833, N4832, N4831, 
        N4830, N4829, N4828, N4827, N4826, N4825, N4824, N4823, N4822, N4821, 
        N4820}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_39 add_103_I2_I4 ( 
        .A({matrix_mul_2D_3__1__20_, matrix_mul_2D_3__1__19_, 
        matrix_mul_2D_3__1__18_, matrix_mul_2D_3__1__17_, 
        matrix_mul_2D_3__1__16_, matrix_mul_2D_3__1__15_, 
        matrix_mul_2D_3__1__14_, matrix_mul_2D_3__1__13_, 
        matrix_mul_2D_3__1__12_, matrix_mul_2D_3__1__11_, 
        matrix_mul_2D_3__1__10_, matrix_mul_2D_3__1__9_, 
        matrix_mul_2D_3__1__8_, matrix_mul_2D_3__1__7_, matrix_mul_2D_3__1__6_, 
        matrix_mul_2D_3__1__5_, matrix_mul_2D_3__1__4_, matrix_mul_2D_3__1__3_, 
        matrix_mul_2D_3__1__2_, matrix_mul_2D_3__1__1_, n19350}), .B({n682, 
        n680, n683, n682, n681, n680, N4709, N4708, N4707, N4706, N4705, N4704, 
        N4703, N4702, N4701, N4700, N4699, N4698, N4697, N4696, N4695}), .SUM(
        {N4748, N4747, N4746, N4745, N4744, N4743, N4742, N4741, N4740, N4739, 
        N4738, N4737, N4736, N4735, N4734, N4733, N4732, N4731, N4730, N4729, 
        N4728}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_40 add_103_I4 ( 
        .A({matrix_mul_2D_3__0__20_, matrix_mul_2D_3__0__19_, 
        matrix_mul_2D_3__0__18_, matrix_mul_2D_3__0__17_, 
        matrix_mul_2D_3__0__16_, matrix_mul_2D_3__0__15_, 
        matrix_mul_2D_3__0__14_, matrix_mul_2D_3__0__13_, 
        matrix_mul_2D_3__0__12_, matrix_mul_2D_3__0__11_, 
        matrix_mul_2D_3__0__10_, matrix_mul_2D_3__0__9_, 
        matrix_mul_2D_3__0__8_, matrix_mul_2D_3__0__7_, matrix_mul_2D_3__0__6_, 
        matrix_mul_2D_3__0__5_, matrix_mul_2D_3__0__4_, matrix_mul_2D_3__0__3_, 
        matrix_mul_2D_3__0__2_, matrix_mul_2D_3__0__1_, n19351}), .B({n677, 
        n675, n678, n677, n676, n675, N4627, N4626, N4625, N4624, N4623, N4622, 
        N4621, N4620, N4619, N4618, N4617, N4616, N4615, N4614, N4613}), .SUM(
        {N4666, N4665, N4664, N4663, N4662, N4661, N4660, N4659, N4658, N4657, 
        N4656, N4655, N4654, N4653, N4652, N4651, N4650, N4649, N4648, N4647, 
        N4646}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_41 add_103_I8_I3 ( 
        .A({matrix_mul_2D_2__7__20_, matrix_mul_2D_2__7__19_, 
        matrix_mul_2D_2__7__18_, matrix_mul_2D_2__7__17_, 
        matrix_mul_2D_2__7__16_, matrix_mul_2D_2__7__15_, 
        matrix_mul_2D_2__7__14_, matrix_mul_2D_2__7__13_, 
        matrix_mul_2D_2__7__12_, matrix_mul_2D_2__7__11_, 
        matrix_mul_2D_2__7__10_, matrix_mul_2D_2__7__9_, 
        matrix_mul_2D_2__7__8_, matrix_mul_2D_2__7__7_, matrix_mul_2D_2__7__6_, 
        matrix_mul_2D_2__7__5_, matrix_mul_2D_2__7__4_, matrix_mul_2D_2__7__3_, 
        matrix_mul_2D_2__7__2_, matrix_mul_2D_2__7__1_, matrix_mul_2D_2__7__0_}), .B({n672, n670, n673, n672, n671, n670, N4527, N4526, N4525, N4524, N4523, 
        N4522, N4521, N4520, N4519, N4518, N4517, N4516, N4515, N4514, N4513}), 
        .SUM({N4566, N4565, N4564, N4563, N4562, N4561, N4560, N4559, N4558, 
        N4557, N4556, N4555, N4554, N4553, N4552, N4551, N4550, N4549, N4548, 
        N4547, N4546}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_42 add_103_I7_I3 ( 
        .A({matrix_mul_2D_2__6__20_, matrix_mul_2D_2__6__19_, 
        matrix_mul_2D_2__6__18_, matrix_mul_2D_2__6__17_, 
        matrix_mul_2D_2__6__16_, matrix_mul_2D_2__6__15_, 
        matrix_mul_2D_2__6__14_, matrix_mul_2D_2__6__13_, 
        matrix_mul_2D_2__6__12_, matrix_mul_2D_2__6__11_, 
        matrix_mul_2D_2__6__10_, matrix_mul_2D_2__6__9_, 
        matrix_mul_2D_2__6__8_, matrix_mul_2D_2__6__7_, matrix_mul_2D_2__6__6_, 
        matrix_mul_2D_2__6__5_, matrix_mul_2D_2__6__4_, matrix_mul_2D_2__6__3_, 
        matrix_mul_2D_2__6__2_, matrix_mul_2D_2__6__1_, matrix_mul_2D_2__6__0_}), .B({n667, n665, n668, n667, n666, n665, N4445, N4444, N4443, N4442, N4441, 
        N4440, N4439, N4438, N4437, N4436, N4435, N4434, N4433, N4432, N4431}), 
        .SUM({N4484, N4483, N4482, N4481, N4480, N4479, N4478, N4477, N4476, 
        N4475, N4474, N4473, N4472, N4471, N4470, N4469, N4468, N4467, N4466, 
        N4465, N4464}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_43 add_103_I6_I3 ( 
        .A({matrix_mul_2D_2__5__20_, matrix_mul_2D_2__5__19_, 
        matrix_mul_2D_2__5__18_, matrix_mul_2D_2__5__17_, 
        matrix_mul_2D_2__5__16_, matrix_mul_2D_2__5__15_, 
        matrix_mul_2D_2__5__14_, matrix_mul_2D_2__5__13_, 
        matrix_mul_2D_2__5__12_, matrix_mul_2D_2__5__11_, 
        matrix_mul_2D_2__5__10_, matrix_mul_2D_2__5__9_, 
        matrix_mul_2D_2__5__8_, matrix_mul_2D_2__5__7_, matrix_mul_2D_2__5__6_, 
        matrix_mul_2D_2__5__5_, matrix_mul_2D_2__5__4_, matrix_mul_2D_2__5__3_, 
        matrix_mul_2D_2__5__2_, matrix_mul_2D_2__5__1_, n19352}), .B({n662, 
        n660, n663, n662, n661, n660, N4356, N4355, N4354, N4353, N4352, N4351, 
        N4350, N4349, N4348, N4347, N4346, N4345, N4344, N4343, N4342}), .SUM(
        {N4395, N4394, N4393, N4392, N4391, N4390, N4389, N4388, N4387, N4386, 
        N4385, N4384, N4383, N4382, N4381, N4380, N4379, N4378, N4377, N4376, 
        N4375}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_44 add_103_I5_I3 ( 
        .A({matrix_mul_2D_2__4__20_, matrix_mul_2D_2__4__19_, 
        matrix_mul_2D_2__4__18_, matrix_mul_2D_2__4__17_, 
        matrix_mul_2D_2__4__16_, matrix_mul_2D_2__4__15_, 
        matrix_mul_2D_2__4__14_, matrix_mul_2D_2__4__13_, 
        matrix_mul_2D_2__4__12_, matrix_mul_2D_2__4__11_, 
        matrix_mul_2D_2__4__10_, matrix_mul_2D_2__4__9_, 
        matrix_mul_2D_2__4__8_, matrix_mul_2D_2__4__7_, matrix_mul_2D_2__4__6_, 
        matrix_mul_2D_2__4__5_, matrix_mul_2D_2__4__4_, matrix_mul_2D_2__4__3_, 
        matrix_mul_2D_2__4__2_, matrix_mul_2D_2__4__1_, n19353}), .B({n657, 
        n655, n658, n657, n656, n655, N4277, N4276, N4275, N4274, N4273, N4272, 
        N4271, N4270, N4269, N4268, N4267, N4266, N4265, N4264, N4263}), .SUM(
        {N4316, N4315, N4314, N4313, N4312, N4311, N4310, N4309, N4308, N4307, 
        N4306, N4305, N4304, N4303, N4302, N4301, N4300, N4299, N4298, N4297, 
        N4296}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_45 add_103_I4_I3 ( 
        .A({matrix_mul_2D_2__3__20_, matrix_mul_2D_2__3__19_, 
        matrix_mul_2D_2__3__18_, matrix_mul_2D_2__3__17_, 
        matrix_mul_2D_2__3__16_, matrix_mul_2D_2__3__15_, 
        matrix_mul_2D_2__3__14_, matrix_mul_2D_2__3__13_, 
        matrix_mul_2D_2__3__12_, matrix_mul_2D_2__3__11_, 
        matrix_mul_2D_2__3__10_, matrix_mul_2D_2__3__9_, 
        matrix_mul_2D_2__3__8_, matrix_mul_2D_2__3__7_, matrix_mul_2D_2__3__6_, 
        matrix_mul_2D_2__3__5_, matrix_mul_2D_2__3__4_, matrix_mul_2D_2__3__3_, 
        matrix_mul_2D_2__3__2_, matrix_mul_2D_2__3__1_, n19354}), .B({n652, 
        n650, n653, n652, n651, n650, N4188, N4187, N4186, N4185, N4184, N4183, 
        N4182, N4181, N4180, N4179, N4178, N4177, N4176, N4175, N4174}), .SUM(
        {N4227, N4226, N4225, N4224, N4223, N4222, N4221, N4220, N4219, N4218, 
        N4217, N4216, N4215, N4214, N4213, N4212, N4211, N4210, N4209, N4208, 
        N4207}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_46 add_103_I3_I3 ( 
        .A({matrix_mul_2D_2__2__20_, matrix_mul_2D_2__2__19_, 
        matrix_mul_2D_2__2__18_, matrix_mul_2D_2__2__17_, 
        matrix_mul_2D_2__2__16_, matrix_mul_2D_2__2__15_, 
        matrix_mul_2D_2__2__14_, matrix_mul_2D_2__2__13_, 
        matrix_mul_2D_2__2__12_, matrix_mul_2D_2__2__11_, 
        matrix_mul_2D_2__2__10_, matrix_mul_2D_2__2__9_, 
        matrix_mul_2D_2__2__8_, matrix_mul_2D_2__2__7_, matrix_mul_2D_2__2__6_, 
        matrix_mul_2D_2__2__5_, matrix_mul_2D_2__2__4_, matrix_mul_2D_2__2__3_, 
        matrix_mul_2D_2__2__2_, matrix_mul_2D_2__2__1_, n19355}), .B({n647, 
        n645, n648, n647, n646, n645, N4109, N4108, N4107, N4106, N4105, N4104, 
        N4103, N4102, N4101, N4100, N4099, N4098, N4097, N4096, N4095}), .SUM(
        {N4148, N4147, N4146, N4145, N4144, N4143, N4142, N4141, N4140, N4139, 
        N4138, N4137, N4136, N4135, N4134, N4133, N4132, N4131, N4130, N4129, 
        N4128}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_47 add_103_I2_I3 ( 
        .A({matrix_mul_2D_2__1__20_, matrix_mul_2D_2__1__19_, 
        matrix_mul_2D_2__1__18_, matrix_mul_2D_2__1__17_, 
        matrix_mul_2D_2__1__16_, matrix_mul_2D_2__1__15_, 
        matrix_mul_2D_2__1__14_, matrix_mul_2D_2__1__13_, 
        matrix_mul_2D_2__1__12_, matrix_mul_2D_2__1__11_, 
        matrix_mul_2D_2__1__10_, matrix_mul_2D_2__1__9_, 
        matrix_mul_2D_2__1__8_, matrix_mul_2D_2__1__7_, matrix_mul_2D_2__1__6_, 
        matrix_mul_2D_2__1__5_, matrix_mul_2D_2__1__4_, matrix_mul_2D_2__1__3_, 
        matrix_mul_2D_2__1__2_, matrix_mul_2D_2__1__1_, n19356}), .B({n642, 
        n640, n643, n642, n641, n640, N4020, N4019, N4018, N4017, N4016, N4015, 
        N4014, N4013, N4012, N4011, N4010, N4009, N4008, N4007, N4006}), .SUM(
        {N4059, N4058, N4057, N4056, N4055, N4054, N4053, N4052, N4051, N4050, 
        N4049, N4048, N4047, N4046, N4045, N4044, N4043, N4042, N4041, N4040, 
        N4039}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_48 add_103_I3 ( 
        .A({matrix_mul_2D_2__0__20_, matrix_mul_2D_2__0__19_, 
        matrix_mul_2D_2__0__18_, matrix_mul_2D_2__0__17_, 
        matrix_mul_2D_2__0__16_, matrix_mul_2D_2__0__15_, 
        matrix_mul_2D_2__0__14_, matrix_mul_2D_2__0__13_, 
        matrix_mul_2D_2__0__12_, matrix_mul_2D_2__0__11_, 
        matrix_mul_2D_2__0__10_, matrix_mul_2D_2__0__9_, 
        matrix_mul_2D_2__0__8_, matrix_mul_2D_2__0__7_, matrix_mul_2D_2__0__6_, 
        matrix_mul_2D_2__0__5_, matrix_mul_2D_2__0__4_, matrix_mul_2D_2__0__3_, 
        matrix_mul_2D_2__0__2_, matrix_mul_2D_2__0__1_, n19357}), .B({n637, 
        n635, n638, n637, n636, n635, N3941, N3940, N3939, N3938, N3937, N3936, 
        N3935, N3934, N3933, N3932, N3931, N3930, N3929, N3928, N3927}), .SUM(
        {N3980, N3979, N3978, N3977, N3976, N3975, N3974, N3973, N3972, N3971, 
        N3970, N3969, N3968, N3967, N3966, N3965, N3964, N3963, N3962, N3961, 
        N3960}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_49 add_103_I8_I2 ( 
        .A({matrix_mul_2D_1__7__20_, matrix_mul_2D_1__7__19_, 
        matrix_mul_2D_1__7__18_, matrix_mul_2D_1__7__17_, 
        matrix_mul_2D_1__7__16_, matrix_mul_2D_1__7__15_, 
        matrix_mul_2D_1__7__14_, matrix_mul_2D_1__7__13_, 
        matrix_mul_2D_1__7__12_, matrix_mul_2D_1__7__11_, 
        matrix_mul_2D_1__7__10_, matrix_mul_2D_1__7__9_, 
        matrix_mul_2D_1__7__8_, matrix_mul_2D_1__7__7_, matrix_mul_2D_1__7__6_, 
        matrix_mul_2D_1__7__5_, matrix_mul_2D_1__7__4_, matrix_mul_2D_1__7__3_, 
        matrix_mul_2D_1__7__2_, matrix_mul_2D_1__7__1_, n19358}), .B({n632, 
        n630, n633, n632, n631, n630, N3852, N3851, N3850, N3849, N3848, N3847, 
        N3846, N3845, N3844, N3843, N3842, N3841, N3840, N3839, N3838}), .SUM(
        {N3891, N3890, N3889, N3888, N3887, N3886, N3885, N3884, N3883, N3882, 
        N3881, N3880, N3879, N3878, N3877, N3876, N3875, N3874, N3873, N3872, 
        N3871}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_50 add_103_I7_I2 ( 
        .A({matrix_mul_2D_1__6__20_, matrix_mul_2D_1__6__19_, 
        matrix_mul_2D_1__6__18_, matrix_mul_2D_1__6__17_, 
        matrix_mul_2D_1__6__16_, matrix_mul_2D_1__6__15_, 
        matrix_mul_2D_1__6__14_, matrix_mul_2D_1__6__13_, 
        matrix_mul_2D_1__6__12_, matrix_mul_2D_1__6__11_, 
        matrix_mul_2D_1__6__10_, matrix_mul_2D_1__6__9_, 
        matrix_mul_2D_1__6__8_, matrix_mul_2D_1__6__7_, matrix_mul_2D_1__6__6_, 
        matrix_mul_2D_1__6__5_, matrix_mul_2D_1__6__4_, matrix_mul_2D_1__6__3_, 
        matrix_mul_2D_1__6__2_, matrix_mul_2D_1__6__1_, n19359}), .B({n627, 
        n625, n628, n627, n626, n625, N3770, N3769, N3768, N3767, N3766, N3765, 
        N3764, N3763, N3762, N3761, N3760, N3759, N3758, N3757, N3756}), .SUM(
        {N3809, N3808, N3807, N3806, N3805, N3804, N3803, N3802, N3801, N3800, 
        N3799, N3798, N3797, N3796, N3795, N3794, N3793, N3792, N3791, N3790, 
        N3789}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_51 add_103_I6_I2 ( 
        .A({matrix_mul_2D_1__5__20_, matrix_mul_2D_1__5__19_, 
        matrix_mul_2D_1__5__18_, matrix_mul_2D_1__5__17_, 
        matrix_mul_2D_1__5__16_, matrix_mul_2D_1__5__15_, 
        matrix_mul_2D_1__5__14_, matrix_mul_2D_1__5__13_, 
        matrix_mul_2D_1__5__12_, matrix_mul_2D_1__5__11_, 
        matrix_mul_2D_1__5__10_, matrix_mul_2D_1__5__9_, 
        matrix_mul_2D_1__5__8_, matrix_mul_2D_1__5__7_, matrix_mul_2D_1__5__6_, 
        matrix_mul_2D_1__5__5_, matrix_mul_2D_1__5__4_, matrix_mul_2D_1__5__3_, 
        matrix_mul_2D_1__5__2_, matrix_mul_2D_1__5__1_, matrix_mul_2D_1__5__0_}), .B({n622, n620, n623, n622, n621, n620, N3681, N3680, N3679, N3678, N3677, 
        N3676, N3675, N3674, N3673, N3672, N3671, N3670, N3669, N3668, N3667}), 
        .SUM({N3720, N3719, N3718, N3717, N3716, N3715, N3714, N3713, N3712, 
        N3711, N3710, N3709, N3708, N3707, N3706, N3705, N3704, N3703, N3702, 
        N3701, N3700}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_52 add_103_I5_I2 ( 
        .A({matrix_mul_2D_1__4__20_, matrix_mul_2D_1__4__19_, 
        matrix_mul_2D_1__4__18_, matrix_mul_2D_1__4__17_, 
        matrix_mul_2D_1__4__16_, matrix_mul_2D_1__4__15_, 
        matrix_mul_2D_1__4__14_, matrix_mul_2D_1__4__13_, 
        matrix_mul_2D_1__4__12_, matrix_mul_2D_1__4__11_, 
        matrix_mul_2D_1__4__10_, matrix_mul_2D_1__4__9_, 
        matrix_mul_2D_1__4__8_, matrix_mul_2D_1__4__7_, matrix_mul_2D_1__4__6_, 
        matrix_mul_2D_1__4__5_, matrix_mul_2D_1__4__4_, matrix_mul_2D_1__4__3_, 
        matrix_mul_2D_1__4__2_, matrix_mul_2D_1__4__1_, matrix_mul_2D_1__4__0_}), .B({n617, n615, n618, n617, n616, n615, N3602, N3601, N3600, N3599, N3598, 
        N3597, N3596, N3595, N3594, N3593, N3592, N3591, N3590, N3589, N3588}), 
        .SUM({N3641, N3640, N3639, N3638, N3637, N3636, N3635, N3634, N3633, 
        N3632, N3631, N3630, N3629, N3628, N3627, N3626, N3625, N3624, N3623, 
        N3622, N3621}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_53 add_103_I4_I2 ( 
        .A({matrix_mul_2D_1__3__20_, matrix_mul_2D_1__3__19_, 
        matrix_mul_2D_1__3__18_, matrix_mul_2D_1__3__17_, 
        matrix_mul_2D_1__3__16_, matrix_mul_2D_1__3__15_, 
        matrix_mul_2D_1__3__14_, matrix_mul_2D_1__3__13_, 
        matrix_mul_2D_1__3__12_, matrix_mul_2D_1__3__11_, 
        matrix_mul_2D_1__3__10_, matrix_mul_2D_1__3__9_, 
        matrix_mul_2D_1__3__8_, matrix_mul_2D_1__3__7_, matrix_mul_2D_1__3__6_, 
        matrix_mul_2D_1__3__5_, matrix_mul_2D_1__3__4_, matrix_mul_2D_1__3__3_, 
        matrix_mul_2D_1__3__2_, matrix_mul_2D_1__3__1_, matrix_mul_2D_1__3__0_}), .B({n612, n610, n613, n612, n611, n610, N3513, N3512, N3511, N3510, N3509, 
        N3508, N3507, N3506, N3505, N3504, N3503, N3502, N3501, N3500, N3499}), 
        .SUM({N3552, N3551, N3550, N3549, N3548, N3547, N3546, N3545, N3544, 
        N3543, N3542, N3541, N3540, N3539, N3538, N3537, N3536, N3535, N3534, 
        N3533, N3532}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_54 add_103_I3_I2 ( 
        .A({matrix_mul_2D_1__2__20_, matrix_mul_2D_1__2__19_, 
        matrix_mul_2D_1__2__18_, matrix_mul_2D_1__2__17_, 
        matrix_mul_2D_1__2__16_, matrix_mul_2D_1__2__15_, 
        matrix_mul_2D_1__2__14_, matrix_mul_2D_1__2__13_, 
        matrix_mul_2D_1__2__12_, matrix_mul_2D_1__2__11_, 
        matrix_mul_2D_1__2__10_, matrix_mul_2D_1__2__9_, 
        matrix_mul_2D_1__2__8_, matrix_mul_2D_1__2__7_, matrix_mul_2D_1__2__6_, 
        matrix_mul_2D_1__2__5_, matrix_mul_2D_1__2__4_, matrix_mul_2D_1__2__3_, 
        matrix_mul_2D_1__2__2_, matrix_mul_2D_1__2__1_, matrix_mul_2D_1__2__0_}), .B({n607, n605, n608, n607, n606, n605, N3434, N3433, N3432, N3431, N3430, 
        N3429, N3428, N3427, N3426, N3425, N3424, N3423, N3422, N3421, N3420}), 
        .SUM({N3473, N3472, N3471, N3470, N3469, N3468, N3467, N3466, N3465, 
        N3464, N3463, N3462, N3461, N3460, N3459, N3458, N3457, N3456, N3455, 
        N3454, N3453}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_55 add_103_I2_I2 ( 
        .A({matrix_mul_2D_1__1__20_, matrix_mul_2D_1__1__19_, 
        matrix_mul_2D_1__1__18_, matrix_mul_2D_1__1__17_, 
        matrix_mul_2D_1__1__16_, matrix_mul_2D_1__1__15_, 
        matrix_mul_2D_1__1__14_, matrix_mul_2D_1__1__13_, 
        matrix_mul_2D_1__1__12_, matrix_mul_2D_1__1__11_, 
        matrix_mul_2D_1__1__10_, matrix_mul_2D_1__1__9_, 
        matrix_mul_2D_1__1__8_, matrix_mul_2D_1__1__7_, matrix_mul_2D_1__1__6_, 
        matrix_mul_2D_1__1__5_, matrix_mul_2D_1__1__4_, matrix_mul_2D_1__1__3_, 
        matrix_mul_2D_1__1__2_, matrix_mul_2D_1__1__1_, n19360}), .B({n602, 
        n600, n603, n602, n601, n600, N3345, N3344, N3343, N3342, N3341, N3340, 
        N3339, N3338, N3337, N3336, N3335, N3334, N3333, N3332, N3331}), .SUM(
        {N3384, N3383, N3382, N3381, N3380, N3379, N3378, N3377, N3376, N3375, 
        N3374, N3373, N3372, N3371, N3370, N3369, N3368, N3367, N3366, N3365, 
        N3364}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_56 add_103_I2 ( 
        .A({matrix_mul_2D_1__0__20_, matrix_mul_2D_1__0__19_, 
        matrix_mul_2D_1__0__18_, matrix_mul_2D_1__0__17_, 
        matrix_mul_2D_1__0__16_, matrix_mul_2D_1__0__15_, 
        matrix_mul_2D_1__0__14_, matrix_mul_2D_1__0__13_, 
        matrix_mul_2D_1__0__12_, matrix_mul_2D_1__0__11_, 
        matrix_mul_2D_1__0__10_, matrix_mul_2D_1__0__9_, 
        matrix_mul_2D_1__0__8_, matrix_mul_2D_1__0__7_, matrix_mul_2D_1__0__6_, 
        matrix_mul_2D_1__0__5_, matrix_mul_2D_1__0__4_, matrix_mul_2D_1__0__3_, 
        matrix_mul_2D_1__0__2_, matrix_mul_2D_1__0__1_, n19361}), .B({n597, 
        n595, n598, n597, n596, n595, N3266, N3265, N3264, N3263, N3262, N3261, 
        N3260, N3259, N3258, N3257, N3256, N3255, N3254, N3253, N3252}), .SUM(
        {N3305, N3304, N3303, N3302, N3301, N3300, N3299, N3298, N3297, N3296, 
        N3295, N3294, N3293, N3292, N3291, N3290, N3289, N3288, N3287, N3286, 
        N3285}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_57 add_103_I8_I1 ( 
        .A({matrix_mul_2D_0__7__20_, matrix_mul_2D_0__7__19_, 
        matrix_mul_2D_0__7__18_, matrix_mul_2D_0__7__17_, 
        matrix_mul_2D_0__7__16_, matrix_mul_2D_0__7__15_, 
        matrix_mul_2D_0__7__14_, matrix_mul_2D_0__7__13_, 
        matrix_mul_2D_0__7__12_, matrix_mul_2D_0__7__11_, 
        matrix_mul_2D_0__7__10_, matrix_mul_2D_0__7__9_, 
        matrix_mul_2D_0__7__8_, matrix_mul_2D_0__7__7_, matrix_mul_2D_0__7__6_, 
        matrix_mul_2D_0__7__5_, matrix_mul_2D_0__7__4_, matrix_mul_2D_0__7__3_, 
        matrix_mul_2D_0__7__2_, matrix_mul_2D_0__7__1_, matrix_mul_2D_0__7__0_}), .B({n592, n590, n593, n592, n591, n590, N3177, N3176, N3175, N3174, N3173, 
        N3172, N3171, N3170, N3169, N3168, N3167, N3166, N3165, N3164, N3163}), 
        .SUM({N3216, N3215, N3214, N3213, N3212, N3211, N3210, N3209, N3208, 
        N3207, N3206, N3205, N3204, N3203, N3202, N3201, N3200, N3199, N3198, 
        N3197, N3196}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_58 add_103_I7_I1 ( 
        .A({matrix_mul_2D_0__6__20_, matrix_mul_2D_0__6__19_, 
        matrix_mul_2D_0__6__18_, matrix_mul_2D_0__6__17_, 
        matrix_mul_2D_0__6__16_, matrix_mul_2D_0__6__15_, 
        matrix_mul_2D_0__6__14_, matrix_mul_2D_0__6__13_, 
        matrix_mul_2D_0__6__12_, matrix_mul_2D_0__6__11_, 
        matrix_mul_2D_0__6__10_, matrix_mul_2D_0__6__9_, 
        matrix_mul_2D_0__6__8_, matrix_mul_2D_0__6__7_, matrix_mul_2D_0__6__6_, 
        matrix_mul_2D_0__6__5_, matrix_mul_2D_0__6__4_, matrix_mul_2D_0__6__3_, 
        matrix_mul_2D_0__6__2_, matrix_mul_2D_0__6__1_, n19362}), .B({n587, 
        n585, n588, n587, n586, n585, N3095, N3094, N3093, N3092, N3091, N3090, 
        N3089, N3088, N3087, N3086, N3085, N3084, N3083, N3082, N3081}), .SUM(
        {N3134, N3133, N3132, N3131, N3130, N3129, N3128, N3127, N3126, N3125, 
        N3124, N3123, N3122, N3121, N3120, N3119, N3118, N3117, N3116, N3115, 
        N3114}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_59 add_103_I6_I1 ( 
        .A({matrix_mul_2D_0__5__20_, matrix_mul_2D_0__5__19_, 
        matrix_mul_2D_0__5__18_, matrix_mul_2D_0__5__17_, 
        matrix_mul_2D_0__5__16_, matrix_mul_2D_0__5__15_, 
        matrix_mul_2D_0__5__14_, matrix_mul_2D_0__5__13_, 
        matrix_mul_2D_0__5__12_, matrix_mul_2D_0__5__11_, 
        matrix_mul_2D_0__5__10_, matrix_mul_2D_0__5__9_, 
        matrix_mul_2D_0__5__8_, matrix_mul_2D_0__5__7_, matrix_mul_2D_0__5__6_, 
        matrix_mul_2D_0__5__5_, matrix_mul_2D_0__5__4_, matrix_mul_2D_0__5__3_, 
        matrix_mul_2D_0__5__2_, matrix_mul_2D_0__5__1_, matrix_mul_2D_0__5__0_}), .B({n582, n580, n583, n582, n581, n580, N3003, N3002, N3001, N3000, N2999, 
        N2998, N2997, N2996, N2995, N2994, N2993, N2992, N2991, N2990, N2989}), 
        .SUM({N3042, N3041, N3040, N3039, N3038, N3037, N3036, N3035, N3034, 
        N3033, N3032, N3031, N3030, N3029, N3028, N3027, N3026, N3025, N3024, 
        N3023, N3022}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_60 add_103_I5_I1 ( 
        .A({matrix_mul_2D_0__4__20_, matrix_mul_2D_0__4__19_, 
        matrix_mul_2D_0__4__18_, matrix_mul_2D_0__4__17_, 
        matrix_mul_2D_0__4__16_, matrix_mul_2D_0__4__15_, 
        matrix_mul_2D_0__4__14_, matrix_mul_2D_0__4__13_, 
        matrix_mul_2D_0__4__12_, matrix_mul_2D_0__4__11_, 
        matrix_mul_2D_0__4__10_, matrix_mul_2D_0__4__9_, 
        matrix_mul_2D_0__4__8_, matrix_mul_2D_0__4__7_, matrix_mul_2D_0__4__6_, 
        matrix_mul_2D_0__4__5_, matrix_mul_2D_0__4__4_, matrix_mul_2D_0__4__3_, 
        matrix_mul_2D_0__4__2_, matrix_mul_2D_0__4__1_, n19363}), .B({n577, 
        n575, n578, n577, n576, n575, N2921, N2920, N2919, N2918, N2917, N2916, 
        N2915, N2914, N2913, N2912, N2911, N2910, N2909, N2908, N2907}), .SUM(
        {N2960, N2959, N2958, N2957, N2956, N2955, N2954, N2953, N2952, N2951, 
        N2950, N2949, N2948, N2947, N2946, N2945, N2944, N2943, N2942, N2941, 
        N2940}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_61 add_103_I4_I1 ( 
        .A({matrix_mul_2D_0__3__20_, matrix_mul_2D_0__3__19_, 
        matrix_mul_2D_0__3__18_, matrix_mul_2D_0__3__17_, 
        matrix_mul_2D_0__3__16_, matrix_mul_2D_0__3__15_, 
        matrix_mul_2D_0__3__14_, matrix_mul_2D_0__3__13_, 
        matrix_mul_2D_0__3__12_, matrix_mul_2D_0__3__11_, 
        matrix_mul_2D_0__3__10_, matrix_mul_2D_0__3__9_, 
        matrix_mul_2D_0__3__8_, matrix_mul_2D_0__3__7_, matrix_mul_2D_0__3__6_, 
        matrix_mul_2D_0__3__5_, matrix_mul_2D_0__3__4_, matrix_mul_2D_0__3__3_, 
        matrix_mul_2D_0__3__2_, matrix_mul_2D_0__3__1_, n19364}), .B({n572, 
        n570, n573, n572, n571, n570, N2829, N2828, N2827, N2826, N2825, N2824, 
        N2823, N2822, N2821, N2820, N2819, N2818, N2817, N2816, N2815}), .SUM(
        {N2868, N2867, N2866, N2865, N2864, N2863, N2862, N2861, N2860, N2859, 
        N2858, N2857, N2856, N2855, N2854, N2853, N2852, N2851, N2850, N2849, 
        N2848}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_62 add_103_I3_I1 ( 
        .A({matrix_mul_2D_0__2__20_, matrix_mul_2D_0__2__19_, 
        matrix_mul_2D_0__2__18_, matrix_mul_2D_0__2__17_, 
        matrix_mul_2D_0__2__16_, matrix_mul_2D_0__2__15_, 
        matrix_mul_2D_0__2__14_, matrix_mul_2D_0__2__13_, 
        matrix_mul_2D_0__2__12_, matrix_mul_2D_0__2__11_, 
        matrix_mul_2D_0__2__10_, matrix_mul_2D_0__2__9_, 
        matrix_mul_2D_0__2__8_, matrix_mul_2D_0__2__7_, matrix_mul_2D_0__2__6_, 
        matrix_mul_2D_0__2__5_, matrix_mul_2D_0__2__4_, matrix_mul_2D_0__2__3_, 
        matrix_mul_2D_0__2__2_, matrix_mul_2D_0__2__1_, n19365}), .B({n567, 
        n565, n568, n567, n566, n565, N2747, N2746, N2745, N2744, N2743, N2742, 
        N2741, N2740, N2739, N2738, N2737, N2736, N2735, N2734, N2733}), .SUM(
        {N2786, N2785, N2784, N2783, N2782, N2781, N2780, N2779, N2778, N2777, 
        N2776, N2775, N2774, N2773, N2772, N2771, N2770, N2769, N2768, N2767, 
        N2766}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_63 add_103_I2_I1 ( 
        .A({matrix_mul_2D_0__1__20_, matrix_mul_2D_0__1__19_, 
        matrix_mul_2D_0__1__18_, matrix_mul_2D_0__1__17_, 
        matrix_mul_2D_0__1__16_, matrix_mul_2D_0__1__15_, 
        matrix_mul_2D_0__1__14_, matrix_mul_2D_0__1__13_, 
        matrix_mul_2D_0__1__12_, matrix_mul_2D_0__1__11_, 
        matrix_mul_2D_0__1__10_, matrix_mul_2D_0__1__9_, 
        matrix_mul_2D_0__1__8_, matrix_mul_2D_0__1__7_, matrix_mul_2D_0__1__6_, 
        matrix_mul_2D_0__1__5_, matrix_mul_2D_0__1__4_, matrix_mul_2D_0__1__3_, 
        matrix_mul_2D_0__1__2_, matrix_mul_2D_0__1__1_, n19366}), .B({n562, 
        n560, n563, n562, n561, n560, N2655, N2654, N2653, N2652, N2651, N2650, 
        N2649, N2648, N2647, N2646, N2645, N2644, N2643, N2642, N2641}), .SUM(
        {N2694, N2693, N2692, N2691, N2690, N2689, N2688, N2687, N2686, N2685, 
        N2684, N2683, N2682, N2681, N2680, N2679, N2678, N2677, N2676, N2675, 
        N2674}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW01_add_64 add_103 ( .A(
        {matrix_mul_2D_0__0__20_, matrix_mul_2D_0__0__19_, 
        matrix_mul_2D_0__0__18_, matrix_mul_2D_0__0__17_, 
        matrix_mul_2D_0__0__16_, matrix_mul_2D_0__0__15_, 
        matrix_mul_2D_0__0__14_, matrix_mul_2D_0__0__13_, 
        matrix_mul_2D_0__0__12_, matrix_mul_2D_0__0__11_, 
        matrix_mul_2D_0__0__10_, matrix_mul_2D_0__0__9_, 
        matrix_mul_2D_0__0__8_, matrix_mul_2D_0__0__7_, matrix_mul_2D_0__0__6_, 
        matrix_mul_2D_0__0__5_, matrix_mul_2D_0__0__4_, matrix_mul_2D_0__0__3_, 
        matrix_mul_2D_0__0__2_, matrix_mul_2D_0__0__1_, n19327}), .B({n557, 
        n555, n558, n557, n556, n555, N2573, N2572, N2571, N2570, N2569, N2568, 
        N2567, N2566, N2565, N2564, N2563, N2562, N2561, N2560, N2559}), .SUM(
        {N2612, N2611, N2610, N2609, N2608, N2607, N2606, N2605, N2604, N2603, 
        N2602, N2601, N2600, N2599, N2598, N2597, N2596, N2595, N2594, N2593, 
        N2592}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_63 r895 ( .A({
        weight_queue_0__0__7_, weight_queue_0__0__6_, weight_queue_0__0__5_, 
        weight_queue_0__0__4_, weight_queue_0__0__3_, weight_queue_0__0__2_, 
        weight_queue_0__0__1_, weight_queue_0__0__0_}), .B({
        data_queue_0__0__7_, data_queue_0__0__6_, data_queue_0__0__5_, 
        data_queue_0__0__4_, data_queue_0__0__3_, data_queue_0__0__2_, 
        data_queue_0__0__1_, data_queue_0__0__0_}), .PRODUCT({N2574, N2573, 
        N2572, N2571, N2570, N2569, N2568, N2567, N2566, N2565, N2564, N2563, 
        N2562, N2561, N2560, N2559}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_62 r900 ( .A({
        weight_queue_0__1__7_, weight_queue_0__1__6_, weight_queue_0__1__5_, 
        weight_queue_0__1__4_, weight_queue_0__1__3_, weight_queue_0__1__2_, 
        weight_queue_0__1__1_, weight_queue_0__1__0_}), .B({
        data_queue_0__1__7_, data_queue_0__1__6_, data_queue_0__1__5_, 
        data_queue_0__1__4_, data_queue_0__1__3_, data_queue_0__1__2_, 
        data_queue_0__1__1_, data_queue_0__1__0_}), .PRODUCT({N2656, N2655, 
        N2654, N2653, N2652, N2651, N2650, N2649, N2648, N2647, N2646, N2645, 
        N2644, N2643, N2642, N2641}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_61 r905 ( .A({
        weight_queue_0__2__7_, weight_queue_0__2__6_, weight_queue_0__2__5_, 
        weight_queue_0__2__4_, weight_queue_0__2__3_, weight_queue_0__2__2_, 
        weight_queue_0__2__1_, weight_queue_0__2__0_}), .B({
        data_queue_0__2__7_, data_queue_0__2__6_, data_queue_0__2__5_, 
        data_queue_0__2__4_, data_queue_0__2__3_, data_queue_0__2__2_, 
        data_queue_0__2__1_, data_queue_0__2__0_}), .PRODUCT({N2748, N2747, 
        N2746, N2745, N2744, N2743, N2742, N2741, N2740, N2739, N2738, N2737, 
        N2736, N2735, N2734, N2733}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_60 r910 ( .A({
        weight_queue_0__3__7_, weight_queue_0__3__6_, weight_queue_0__3__5_, 
        weight_queue_0__3__4_, weight_queue_0__3__3_, weight_queue_0__3__2_, 
        weight_queue_0__3__1_, weight_queue_0__3__0_}), .B({
        data_queue_0__3__7_, data_queue_0__3__6_, data_queue_0__3__5_, 
        data_queue_0__3__4_, data_queue_0__3__3_, data_queue_0__3__2_, 
        data_queue_0__3__1_, data_queue_0__3__0_}), .PRODUCT({N2830, N2829, 
        N2828, N2827, N2826, N2825, N2824, N2823, N2822, N2821, N2820, N2819, 
        N2818, N2817, N2816, N2815}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_59 r915 ( .A({
        weight_queue_0__4__7_, weight_queue_0__4__6_, weight_queue_0__4__5_, 
        weight_queue_0__4__4_, weight_queue_0__4__3_, weight_queue_0__4__2_, 
        weight_queue_0__4__1_, weight_queue_0__4__0_}), .B({
        data_queue_0__4__7_, data_queue_0__4__6_, data_queue_0__4__5_, 
        data_queue_0__4__4_, data_queue_0__4__3_, data_queue_0__4__2_, 
        data_queue_0__4__1_, data_queue_0__4__0_}), .PRODUCT({N2922, N2921, 
        N2920, N2919, N2918, N2917, N2916, N2915, N2914, N2913, N2912, N2911, 
        N2910, N2909, N2908, N2907}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_58 r920 ( .A({
        weight_queue_0__5__7_, weight_queue_0__5__6_, weight_queue_0__5__5_, 
        weight_queue_0__5__4_, weight_queue_0__5__3_, weight_queue_0__5__2_, 
        weight_queue_0__5__1_, weight_queue_0__5__0_}), .B({
        data_queue_0__5__7_, data_queue_0__5__6_, data_queue_0__5__5_, 
        data_queue_0__5__4_, data_queue_0__5__3_, data_queue_0__5__2_, 
        data_queue_0__5__1_, data_queue_0__5__0_}), .PRODUCT({N3004, N3003, 
        N3002, N3001, N3000, N2999, N2998, N2997, N2996, N2995, N2994, N2993, 
        N2992, N2991, N2990, N2989}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_57 r925 ( .A({
        weight_queue_0__6__7_, weight_queue_0__6__6_, weight_queue_0__6__5_, 
        weight_queue_0__6__4_, weight_queue_0__6__3_, weight_queue_0__6__2_, 
        weight_queue_0__6__1_, weight_queue_0__6__0_}), .B({
        data_queue_0__6__7_, data_queue_0__6__6_, data_queue_0__6__5_, 
        data_queue_0__6__4_, data_queue_0__6__3_, data_queue_0__6__2_, 
        data_queue_0__6__1_, data_queue_0__6__0_}), .PRODUCT({N3096, N3095, 
        N3094, N3093, N3092, N3091, N3090, N3089, N3088, N3087, N3086, N3085, 
        N3084, N3083, N3082, N3081}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_56 r930 ( .A({
        weight_queue_0__7__7_, weight_queue_0__7__6_, weight_queue_0__7__5_, 
        weight_queue_0__7__4_, weight_queue_0__7__3_, weight_queue_0__7__2_, 
        weight_queue_0__7__1_, weight_queue_0__7__0_}), .B({n19750, n19747, 
        n19744, n19741, n19738, n19735, n19732, n19729}), .PRODUCT({N3178, 
        N3177, N3176, N3175, N3174, N3173, N3172, N3171, N3170, N3169, N3168, 
        N3167, N3166, N3165, N3164, N3163}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_55 r932 ( .A({
        weight_queue_1__0__7_, weight_queue_1__0__6_, weight_queue_1__0__5_, 
        weight_queue_1__0__4_, weight_queue_1__0__3_, weight_queue_1__0__2_, 
        weight_queue_1__0__1_, weight_queue_1__0__0_}), .B({
        data_queue_1__0__7_, data_queue_1__0__6_, data_queue_1__0__5_, 
        data_queue_1__0__4_, data_queue_1__0__3_, data_queue_1__0__2_, 
        data_queue_1__0__1_, data_queue_1__0__0_}), .PRODUCT({N3267, N3266, 
        N3265, N3264, N3263, N3262, N3261, N3260, N3259, N3258, N3257, N3256, 
        N3255, N3254, N3253, N3252}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_54 r934 ( .A({
        weight_queue_1__1__7_, weight_queue_1__1__6_, weight_queue_1__1__5_, 
        weight_queue_1__1__4_, weight_queue_1__1__3_, weight_queue_1__1__2_, 
        weight_queue_1__1__1_, weight_queue_1__1__0_}), .B({
        data_queue_1__1__7_, data_queue_1__1__6_, data_queue_1__1__5_, 
        data_queue_1__1__4_, data_queue_1__1__3_, data_queue_1__1__2_, 
        data_queue_1__1__1_, data_queue_1__1__0_}), .PRODUCT({N3346, N3345, 
        N3344, N3343, N3342, N3341, N3340, N3339, N3338, N3337, N3336, N3335, 
        N3334, N3333, N3332, N3331}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_53 r936 ( .A({
        weight_queue_1__2__7_, weight_queue_1__2__6_, weight_queue_1__2__5_, 
        weight_queue_1__2__4_, weight_queue_1__2__3_, weight_queue_1__2__2_, 
        weight_queue_1__2__1_, weight_queue_1__2__0_}), .B({
        data_queue_1__2__7_, data_queue_1__2__6_, data_queue_1__2__5_, 
        data_queue_1__2__4_, data_queue_1__2__3_, data_queue_1__2__2_, 
        data_queue_1__2__1_, data_queue_1__2__0_}), .PRODUCT({N3435, N3434, 
        N3433, N3432, N3431, N3430, N3429, N3428, N3427, N3426, N3425, N3424, 
        N3423, N3422, N3421, N3420}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_52 r938 ( .A({
        weight_queue_1__3__7_, weight_queue_1__3__6_, weight_queue_1__3__5_, 
        weight_queue_1__3__4_, weight_queue_1__3__3_, weight_queue_1__3__2_, 
        weight_queue_1__3__1_, weight_queue_1__3__0_}), .B({
        data_queue_1__3__7_, data_queue_1__3__6_, data_queue_1__3__5_, 
        data_queue_1__3__4_, data_queue_1__3__3_, data_queue_1__3__2_, 
        data_queue_1__3__1_, data_queue_1__3__0_}), .PRODUCT({N3514, N3513, 
        N3512, N3511, N3510, N3509, N3508, N3507, N3506, N3505, N3504, N3503, 
        N3502, N3501, N3500, N3499}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_51 r940 ( .A({
        weight_queue_1__4__7_, weight_queue_1__4__6_, weight_queue_1__4__5_, 
        weight_queue_1__4__4_, weight_queue_1__4__3_, weight_queue_1__4__2_, 
        weight_queue_1__4__1_, weight_queue_1__4__0_}), .B({
        data_queue_1__4__7_, data_queue_1__4__6_, data_queue_1__4__5_, 
        data_queue_1__4__4_, data_queue_1__4__3_, data_queue_1__4__2_, 
        data_queue_1__4__1_, data_queue_1__4__0_}), .PRODUCT({N3603, N3602, 
        N3601, N3600, N3599, N3598, N3597, N3596, N3595, N3594, N3593, N3592, 
        N3591, N3590, N3589, N3588}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_50 r942 ( .A({
        weight_queue_1__5__7_, weight_queue_1__5__6_, weight_queue_1__5__5_, 
        weight_queue_1__5__4_, weight_queue_1__5__3_, weight_queue_1__5__2_, 
        weight_queue_1__5__1_, weight_queue_1__5__0_}), .B({
        data_queue_1__5__7_, data_queue_1__5__6_, data_queue_1__5__5_, 
        data_queue_1__5__4_, data_queue_1__5__3_, data_queue_1__5__2_, 
        data_queue_1__5__1_, data_queue_1__5__0_}), .PRODUCT({N3682, N3681, 
        N3680, N3679, N3678, N3677, N3676, N3675, N3674, N3673, N3672, N3671, 
        N3670, N3669, N3668, N3667}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_49 r944 ( .A({
        weight_queue_1__6__7_, weight_queue_1__6__6_, weight_queue_1__6__5_, 
        weight_queue_1__6__4_, weight_queue_1__6__3_, weight_queue_1__6__2_, 
        weight_queue_1__6__1_, weight_queue_1__6__0_}), .B({
        data_queue_1__6__7_, data_queue_1__6__6_, data_queue_1__6__5_, 
        data_queue_1__6__4_, data_queue_1__6__3_, data_queue_1__6__2_, 
        data_queue_1__6__1_, data_queue_1__6__0_}), .PRODUCT({N3771, N3770, 
        N3769, N3768, N3767, N3766, N3765, N3764, N3763, N3762, N3761, N3760, 
        N3759, N3758, N3757, N3756}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_48 r949 ( .A({
        weight_queue_1__7__7_, weight_queue_1__7__6_, weight_queue_1__7__5_, 
        weight_queue_1__7__4_, weight_queue_1__7__3_, weight_queue_1__7__2_, 
        weight_queue_1__7__1_, weight_queue_1__7__0_}), .B({n19726, n19723, 
        n19720, n19717, n19714, n19711, n19708, n19705}), .PRODUCT({N3853, 
        N3852, N3851, N3850, N3849, N3848, N3847, N3846, N3845, N3844, N3843, 
        N3842, N3841, N3840, N3839, N3838}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_47 r951 ( .A({
        weight_queue_2__0__7_, weight_queue_2__0__6_, weight_queue_2__0__5_, 
        weight_queue_2__0__4_, weight_queue_2__0__3_, weight_queue_2__0__2_, 
        weight_queue_2__0__1_, weight_queue_2__0__0_}), .B({
        data_queue_2__0__7_, data_queue_2__0__6_, data_queue_2__0__5_, 
        data_queue_2__0__4_, data_queue_2__0__3_, data_queue_2__0__2_, 
        data_queue_2__0__1_, data_queue_2__0__0_}), .PRODUCT({N3942, N3941, 
        N3940, N3939, N3938, N3937, N3936, N3935, N3934, N3933, N3932, N3931, 
        N3930, N3929, N3928, N3927}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_46 r953 ( .A({
        weight_queue_2__1__7_, weight_queue_2__1__6_, weight_queue_2__1__5_, 
        weight_queue_2__1__4_, weight_queue_2__1__3_, weight_queue_2__1__2_, 
        weight_queue_2__1__1_, weight_queue_2__1__0_}), .B({
        data_queue_2__1__7_, data_queue_2__1__6_, data_queue_2__1__5_, 
        data_queue_2__1__4_, data_queue_2__1__3_, data_queue_2__1__2_, 
        data_queue_2__1__1_, data_queue_2__1__0_}), .PRODUCT({N4021, N4020, 
        N4019, N4018, N4017, N4016, N4015, N4014, N4013, N4012, N4011, N4010, 
        N4009, N4008, N4007, N4006}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_45 r955 ( .A({
        weight_queue_2__2__7_, weight_queue_2__2__6_, weight_queue_2__2__5_, 
        weight_queue_2__2__4_, weight_queue_2__2__3_, weight_queue_2__2__2_, 
        weight_queue_2__2__1_, weight_queue_2__2__0_}), .B({
        data_queue_2__2__7_, data_queue_2__2__6_, data_queue_2__2__5_, 
        data_queue_2__2__4_, data_queue_2__2__3_, data_queue_2__2__2_, 
        data_queue_2__2__1_, data_queue_2__2__0_}), .PRODUCT({N4110, N4109, 
        N4108, N4107, N4106, N4105, N4104, N4103, N4102, N4101, N4100, N4099, 
        N4098, N4097, N4096, N4095}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_44 r957 ( .A({
        weight_queue_2__3__7_, weight_queue_2__3__6_, weight_queue_2__3__5_, 
        weight_queue_2__3__4_, weight_queue_2__3__3_, weight_queue_2__3__2_, 
        weight_queue_2__3__1_, weight_queue_2__3__0_}), .B({
        data_queue_2__3__7_, data_queue_2__3__6_, data_queue_2__3__5_, 
        data_queue_2__3__4_, data_queue_2__3__3_, data_queue_2__3__2_, 
        data_queue_2__3__1_, data_queue_2__3__0_}), .PRODUCT({N4189, N4188, 
        N4187, N4186, N4185, N4184, N4183, N4182, N4181, N4180, N4179, N4178, 
        N4177, N4176, N4175, N4174}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_43 r959 ( .A({
        weight_queue_2__4__7_, weight_queue_2__4__6_, weight_queue_2__4__5_, 
        weight_queue_2__4__4_, weight_queue_2__4__3_, weight_queue_2__4__2_, 
        weight_queue_2__4__1_, weight_queue_2__4__0_}), .B({
        data_queue_2__4__7_, data_queue_2__4__6_, data_queue_2__4__5_, 
        data_queue_2__4__4_, data_queue_2__4__3_, data_queue_2__4__2_, 
        data_queue_2__4__1_, data_queue_2__4__0_}), .PRODUCT({N4278, N4277, 
        N4276, N4275, N4274, N4273, N4272, N4271, N4270, N4269, N4268, N4267, 
        N4266, N4265, N4264, N4263}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_42 r961 ( .A({
        weight_queue_2__5__7_, weight_queue_2__5__6_, weight_queue_2__5__5_, 
        weight_queue_2__5__4_, weight_queue_2__5__3_, weight_queue_2__5__2_, 
        weight_queue_2__5__1_, weight_queue_2__5__0_}), .B({
        data_queue_2__5__7_, data_queue_2__5__6_, data_queue_2__5__5_, 
        data_queue_2__5__4_, data_queue_2__5__3_, data_queue_2__5__2_, 
        data_queue_2__5__1_, data_queue_2__5__0_}), .PRODUCT({N4357, N4356, 
        N4355, N4354, N4353, N4352, N4351, N4350, N4349, N4348, N4347, N4346, 
        N4345, N4344, N4343, N4342}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_41 r963 ( .A({
        weight_queue_2__6__7_, weight_queue_2__6__6_, weight_queue_2__6__5_, 
        weight_queue_2__6__4_, weight_queue_2__6__3_, weight_queue_2__6__2_, 
        weight_queue_2__6__1_, weight_queue_2__6__0_}), .B({
        data_queue_2__6__7_, data_queue_2__6__6_, data_queue_2__6__5_, 
        data_queue_2__6__4_, data_queue_2__6__3_, data_queue_2__6__2_, 
        data_queue_2__6__1_, data_queue_2__6__0_}), .PRODUCT({N4446, N4445, 
        N4444, N4443, N4442, N4441, N4440, N4439, N4438, N4437, N4436, N4435, 
        N4434, N4433, N4432, N4431}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_40 r968 ( .A({
        weight_queue_2__7__7_, weight_queue_2__7__6_, weight_queue_2__7__5_, 
        weight_queue_2__7__4_, weight_queue_2__7__3_, weight_queue_2__7__2_, 
        weight_queue_2__7__1_, weight_queue_2__7__0_}), .B({n19702, n19699, 
        n19696, n19693, n19690, n19687, n19684, n19681}), .PRODUCT({N4528, 
        N4527, N4526, N4525, N4524, N4523, N4522, N4521, N4520, N4519, N4518, 
        N4517, N4516, N4515, N4514, N4513}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_39 r970 ( .A({
        weight_queue_3__0__7_, weight_queue_3__0__6_, weight_queue_3__0__5_, 
        weight_queue_3__0__4_, weight_queue_3__0__3_, weight_queue_3__0__2_, 
        weight_queue_3__0__1_, weight_queue_3__0__0_}), .B({
        data_queue_3__0__7_, data_queue_3__0__6_, data_queue_3__0__5_, 
        data_queue_3__0__4_, data_queue_3__0__3_, data_queue_3__0__2_, 
        data_queue_3__0__1_, data_queue_3__0__0_}), .PRODUCT({N4628, N4627, 
        N4626, N4625, N4624, N4623, N4622, N4621, N4620, N4619, N4618, N4617, 
        N4616, N4615, N4614, N4613}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_38 r972 ( .A({
        weight_queue_3__1__7_, weight_queue_3__1__6_, weight_queue_3__1__5_, 
        weight_queue_3__1__4_, weight_queue_3__1__3_, weight_queue_3__1__2_, 
        weight_queue_3__1__1_, weight_queue_3__1__0_}), .B({
        data_queue_3__1__7_, data_queue_3__1__6_, data_queue_3__1__5_, 
        data_queue_3__1__4_, data_queue_3__1__3_, data_queue_3__1__2_, 
        data_queue_3__1__1_, data_queue_3__1__0_}), .PRODUCT({N4710, N4709, 
        N4708, N4707, N4706, N4705, N4704, N4703, N4702, N4701, N4700, N4699, 
        N4698, N4697, N4696, N4695}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_37 r974 ( .A({
        weight_queue_3__2__7_, weight_queue_3__2__6_, weight_queue_3__2__5_, 
        weight_queue_3__2__4_, weight_queue_3__2__3_, weight_queue_3__2__2_, 
        weight_queue_3__2__1_, weight_queue_3__2__0_}), .B({
        data_queue_3__2__7_, data_queue_3__2__6_, data_queue_3__2__5_, 
        data_queue_3__2__4_, data_queue_3__2__3_, data_queue_3__2__2_, 
        data_queue_3__2__1_, data_queue_3__2__0_}), .PRODUCT({N4802, N4801, 
        N4800, N4799, N4798, N4797, N4796, N4795, N4794, N4793, N4792, N4791, 
        N4790, N4789, N4788, N4787}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_36 r976 ( .A({
        weight_queue_3__3__7_, weight_queue_3__3__6_, weight_queue_3__3__5_, 
        weight_queue_3__3__4_, weight_queue_3__3__3_, weight_queue_3__3__2_, 
        weight_queue_3__3__1_, weight_queue_3__3__0_}), .B({
        data_queue_3__3__7_, data_queue_3__3__6_, data_queue_3__3__5_, 
        data_queue_3__3__4_, data_queue_3__3__3_, data_queue_3__3__2_, 
        data_queue_3__3__1_, data_queue_3__3__0_}), .PRODUCT({N4884, N4883, 
        N4882, N4881, N4880, N4879, N4878, N4877, N4876, N4875, N4874, N4873, 
        N4872, N4871, N4870, N4869}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_35 r978 ( .A({
        weight_queue_3__4__7_, weight_queue_3__4__6_, weight_queue_3__4__5_, 
        weight_queue_3__4__4_, weight_queue_3__4__3_, weight_queue_3__4__2_, 
        weight_queue_3__4__1_, weight_queue_3__4__0_}), .B({
        data_queue_3__4__7_, data_queue_3__4__6_, data_queue_3__4__5_, 
        data_queue_3__4__4_, data_queue_3__4__3_, data_queue_3__4__2_, 
        data_queue_3__4__1_, data_queue_3__4__0_}), .PRODUCT({N4976, N4975, 
        N4974, N4973, N4972, N4971, N4970, N4969, N4968, N4967, N4966, N4965, 
        N4964, N4963, N4962, N4961}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_34 r980 ( .A({
        weight_queue_3__5__7_, weight_queue_3__5__6_, weight_queue_3__5__5_, 
        weight_queue_3__5__4_, weight_queue_3__5__3_, weight_queue_3__5__2_, 
        weight_queue_3__5__1_, weight_queue_3__5__0_}), .B({
        data_queue_3__5__7_, data_queue_3__5__6_, data_queue_3__5__5_, 
        data_queue_3__5__4_, data_queue_3__5__3_, data_queue_3__5__2_, 
        data_queue_3__5__1_, data_queue_3__5__0_}), .PRODUCT({N5058, N5057, 
        N5056, N5055, N5054, N5053, N5052, N5051, N5050, N5049, N5048, N5047, 
        N5046, N5045, N5044, N5043}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_33 r982 ( .A({
        weight_queue_3__6__7_, weight_queue_3__6__6_, weight_queue_3__6__5_, 
        weight_queue_3__6__4_, weight_queue_3__6__3_, weight_queue_3__6__2_, 
        weight_queue_3__6__1_, weight_queue_3__6__0_}), .B({
        data_queue_3__6__7_, data_queue_3__6__6_, data_queue_3__6__5_, 
        data_queue_3__6__4_, data_queue_3__6__3_, data_queue_3__6__2_, 
        data_queue_3__6__1_, data_queue_3__6__0_}), .PRODUCT({N5150, N5149, 
        N5148, N5147, N5146, N5145, N5144, N5143, N5142, N5141, N5140, N5139, 
        N5138, N5137, N5136, N5135}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_32 r987 ( .A({
        weight_queue_3__7__7_, weight_queue_3__7__6_, weight_queue_3__7__5_, 
        weight_queue_3__7__4_, weight_queue_3__7__3_, weight_queue_3__7__2_, 
        weight_queue_3__7__1_, weight_queue_3__7__0_}), .B({n19678, n19675, 
        n19672, n19669, n19666, n19663, n19660, n19657}), .PRODUCT({N5232, 
        N5231, N5230, N5229, N5228, N5227, N5226, N5225, N5224, N5223, N5222, 
        N5221, N5220, N5219, N5218, N5217}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_31 r989 ( .A({
        weight_queue_4__0__7_, weight_queue_4__0__6_, weight_queue_4__0__5_, 
        weight_queue_4__0__4_, weight_queue_4__0__3_, weight_queue_4__0__2_, 
        weight_queue_4__0__1_, weight_queue_4__0__0_}), .B({
        data_queue_4__0__7_, data_queue_4__0__6_, data_queue_4__0__5_, 
        data_queue_4__0__4_, data_queue_4__0__3_, data_queue_4__0__2_, 
        data_queue_4__0__1_, data_queue_4__0__0_}), .PRODUCT({N5321, N5320, 
        N5319, N5318, N5317, N5316, N5315, N5314, N5313, N5312, N5311, N5310, 
        N5309, N5308, N5307, N5306}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_30 r991 ( .A({
        weight_queue_4__1__7_, weight_queue_4__1__6_, weight_queue_4__1__5_, 
        weight_queue_4__1__4_, weight_queue_4__1__3_, weight_queue_4__1__2_, 
        weight_queue_4__1__1_, weight_queue_4__1__0_}), .B({
        data_queue_4__1__7_, data_queue_4__1__6_, data_queue_4__1__5_, 
        data_queue_4__1__4_, data_queue_4__1__3_, data_queue_4__1__2_, 
        data_queue_4__1__1_, data_queue_4__1__0_}), .PRODUCT({N5400, N5399, 
        N5398, N5397, N5396, N5395, N5394, N5393, N5392, N5391, N5390, N5389, 
        N5388, N5387, N5386, N5385}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_29 r993 ( .A({
        weight_queue_4__2__7_, weight_queue_4__2__6_, weight_queue_4__2__5_, 
        weight_queue_4__2__4_, weight_queue_4__2__3_, weight_queue_4__2__2_, 
        weight_queue_4__2__1_, weight_queue_4__2__0_}), .B({
        data_queue_4__2__7_, data_queue_4__2__6_, data_queue_4__2__5_, 
        data_queue_4__2__4_, data_queue_4__2__3_, data_queue_4__2__2_, 
        data_queue_4__2__1_, data_queue_4__2__0_}), .PRODUCT({N5489, N5488, 
        N5487, N5486, N5485, N5484, N5483, N5482, N5481, N5480, N5479, N5478, 
        N5477, N5476, N5475, N5474}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_28 r995 ( .A({
        weight_queue_4__3__7_, weight_queue_4__3__6_, weight_queue_4__3__5_, 
        weight_queue_4__3__4_, weight_queue_4__3__3_, weight_queue_4__3__2_, 
        weight_queue_4__3__1_, weight_queue_4__3__0_}), .B({
        data_queue_4__3__7_, data_queue_4__3__6_, data_queue_4__3__5_, 
        data_queue_4__3__4_, data_queue_4__3__3_, data_queue_4__3__2_, 
        data_queue_4__3__1_, data_queue_4__3__0_}), .PRODUCT({N5568, N5567, 
        N5566, N5565, N5564, N5563, N5562, N5561, N5560, N5559, N5558, N5557, 
        N5556, N5555, N5554, N5553}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_27 r997 ( .A({
        weight_queue_4__4__7_, weight_queue_4__4__6_, weight_queue_4__4__5_, 
        weight_queue_4__4__4_, weight_queue_4__4__3_, weight_queue_4__4__2_, 
        weight_queue_4__4__1_, weight_queue_4__4__0_}), .B({
        data_queue_4__4__7_, data_queue_4__4__6_, data_queue_4__4__5_, 
        data_queue_4__4__4_, data_queue_4__4__3_, data_queue_4__4__2_, 
        data_queue_4__4__1_, data_queue_4__4__0_}), .PRODUCT({N5657, N5656, 
        N5655, N5654, N5653, N5652, N5651, N5650, N5649, N5648, N5647, N5646, 
        N5645, N5644, N5643, N5642}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_26 r999 ( .A({
        weight_queue_4__5__7_, weight_queue_4__5__6_, weight_queue_4__5__5_, 
        weight_queue_4__5__4_, weight_queue_4__5__3_, weight_queue_4__5__2_, 
        weight_queue_4__5__1_, weight_queue_4__5__0_}), .B({
        data_queue_4__5__7_, data_queue_4__5__6_, data_queue_4__5__5_, 
        data_queue_4__5__4_, data_queue_4__5__3_, data_queue_4__5__2_, 
        data_queue_4__5__1_, data_queue_4__5__0_}), .PRODUCT({N5736, N5735, 
        N5734, N5733, N5732, N5731, N5730, N5729, N5728, N5727, N5726, N5725, 
        N5724, N5723, N5722, N5721}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_25 r1001 ( .A({
        weight_queue_4__6__7_, weight_queue_4__6__6_, weight_queue_4__6__5_, 
        weight_queue_4__6__4_, weight_queue_4__6__3_, weight_queue_4__6__2_, 
        weight_queue_4__6__1_, weight_queue_4__6__0_}), .B({
        data_queue_4__6__7_, data_queue_4__6__6_, data_queue_4__6__5_, 
        data_queue_4__6__4_, data_queue_4__6__3_, data_queue_4__6__2_, 
        data_queue_4__6__1_, data_queue_4__6__0_}), .PRODUCT({N5825, N5824, 
        N5823, N5822, N5821, N5820, N5819, N5818, N5817, N5816, N5815, N5814, 
        N5813, N5812, N5811, N5810}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_24 r1006 ( .A({
        weight_queue_4__7__7_, weight_queue_4__7__6_, weight_queue_4__7__5_, 
        weight_queue_4__7__4_, weight_queue_4__7__3_, weight_queue_4__7__2_, 
        weight_queue_4__7__1_, weight_queue_4__7__0_}), .B({n19654, n19651, 
        n19648, n19645, n19642, n19639, n19636, n19633}), .PRODUCT({N5907, 
        N5906, N5905, N5904, N5903, N5902, N5901, N5900, N5899, N5898, N5897, 
        N5896, N5895, N5894, N5893, N5892}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_23 r1008 ( .A({
        weight_queue_5__0__7_, weight_queue_5__0__6_, weight_queue_5__0__5_, 
        weight_queue_5__0__4_, weight_queue_5__0__3_, weight_queue_5__0__2_, 
        weight_queue_5__0__1_, weight_queue_5__0__0_}), .B({
        data_queue_5__0__7_, data_queue_5__0__6_, data_queue_5__0__5_, 
        data_queue_5__0__4_, data_queue_5__0__3_, data_queue_5__0__2_, 
        data_queue_5__0__1_, data_queue_5__0__0_}), .PRODUCT({N5996, N5995, 
        N5994, N5993, N5992, N5991, N5990, N5989, N5988, N5987, N5986, N5985, 
        N5984, N5983, N5982, N5981}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_22 r1010 ( .A({
        weight_queue_5__1__7_, weight_queue_5__1__6_, weight_queue_5__1__5_, 
        weight_queue_5__1__4_, weight_queue_5__1__3_, weight_queue_5__1__2_, 
        weight_queue_5__1__1_, weight_queue_5__1__0_}), .B({
        data_queue_5__1__7_, data_queue_5__1__6_, data_queue_5__1__5_, 
        data_queue_5__1__4_, data_queue_5__1__3_, data_queue_5__1__2_, 
        data_queue_5__1__1_, data_queue_5__1__0_}), .PRODUCT({N6075, N6074, 
        N6073, N6072, N6071, N6070, N6069, N6068, N6067, N6066, N6065, N6064, 
        N6063, N6062, N6061, N6060}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_21 r1012 ( .A({
        weight_queue_5__2__7_, weight_queue_5__2__6_, weight_queue_5__2__5_, 
        weight_queue_5__2__4_, weight_queue_5__2__3_, weight_queue_5__2__2_, 
        weight_queue_5__2__1_, weight_queue_5__2__0_}), .B({
        data_queue_5__2__7_, data_queue_5__2__6_, data_queue_5__2__5_, 
        data_queue_5__2__4_, data_queue_5__2__3_, data_queue_5__2__2_, 
        data_queue_5__2__1_, data_queue_5__2__0_}), .PRODUCT({N6164, N6163, 
        N6162, N6161, N6160, N6159, N6158, N6157, N6156, N6155, N6154, N6153, 
        N6152, N6151, N6150, N6149}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_20 r1014 ( .A({
        weight_queue_5__3__7_, weight_queue_5__3__6_, weight_queue_5__3__5_, 
        weight_queue_5__3__4_, weight_queue_5__3__3_, weight_queue_5__3__2_, 
        weight_queue_5__3__1_, weight_queue_5__3__0_}), .B({
        data_queue_5__3__7_, data_queue_5__3__6_, data_queue_5__3__5_, 
        data_queue_5__3__4_, data_queue_5__3__3_, data_queue_5__3__2_, 
        data_queue_5__3__1_, data_queue_5__3__0_}), .PRODUCT({N6243, N6242, 
        N6241, N6240, N6239, N6238, N6237, N6236, N6235, N6234, N6233, N6232, 
        N6231, N6230, N6229, N6228}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_19 r1016 ( .A({
        weight_queue_5__4__7_, weight_queue_5__4__6_, weight_queue_5__4__5_, 
        weight_queue_5__4__4_, weight_queue_5__4__3_, weight_queue_5__4__2_, 
        weight_queue_5__4__1_, weight_queue_5__4__0_}), .B({
        data_queue_5__4__7_, data_queue_5__4__6_, data_queue_5__4__5_, 
        data_queue_5__4__4_, data_queue_5__4__3_, data_queue_5__4__2_, 
        data_queue_5__4__1_, data_queue_5__4__0_}), .PRODUCT({N6332, N6331, 
        N6330, N6329, N6328, N6327, N6326, N6325, N6324, N6323, N6322, N6321, 
        N6320, N6319, N6318, N6317}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_18 r1018 ( .A({
        weight_queue_5__5__7_, weight_queue_5__5__6_, weight_queue_5__5__5_, 
        weight_queue_5__5__4_, weight_queue_5__5__3_, weight_queue_5__5__2_, 
        weight_queue_5__5__1_, weight_queue_5__5__0_}), .B({
        data_queue_5__5__7_, data_queue_5__5__6_, data_queue_5__5__5_, 
        data_queue_5__5__4_, data_queue_5__5__3_, data_queue_5__5__2_, 
        data_queue_5__5__1_, data_queue_5__5__0_}), .PRODUCT({N6411, N6410, 
        N6409, N6408, N6407, N6406, N6405, N6404, N6403, N6402, N6401, N6400, 
        N6399, N6398, N6397, N6396}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_17 r1020 ( .A({
        weight_queue_5__6__7_, weight_queue_5__6__6_, weight_queue_5__6__5_, 
        weight_queue_5__6__4_, weight_queue_5__6__3_, weight_queue_5__6__2_, 
        weight_queue_5__6__1_, weight_queue_5__6__0_}), .B({
        data_queue_5__6__7_, data_queue_5__6__6_, data_queue_5__6__5_, 
        data_queue_5__6__4_, data_queue_5__6__3_, data_queue_5__6__2_, 
        data_queue_5__6__1_, data_queue_5__6__0_}), .PRODUCT({N6500, N6499, 
        N6498, N6497, N6496, N6495, N6494, N6493, N6492, N6491, N6490, N6489, 
        N6488, N6487, N6486, N6485}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_16 r1025 ( .A({
        weight_queue_5__7__7_, weight_queue_5__7__6_, weight_queue_5__7__5_, 
        weight_queue_5__7__4_, weight_queue_5__7__3_, weight_queue_5__7__2_, 
        weight_queue_5__7__1_, weight_queue_5__7__0_}), .B({n19630, n19627, 
        n19624, n19621, n19618, n19615, n19612, n19609}), .PRODUCT({N6582, 
        N6581, N6580, N6579, N6578, N6577, N6576, N6575, N6574, N6573, N6572, 
        N6571, N6570, N6569, N6568, N6567}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_15 r1027 ( .A({
        weight_queue_6__0__7_, weight_queue_6__0__6_, weight_queue_6__0__5_, 
        weight_queue_6__0__4_, weight_queue_6__0__3_, weight_queue_6__0__2_, 
        weight_queue_6__0__1_, weight_queue_6__0__0_}), .B({
        data_queue_6__0__7_, data_queue_6__0__6_, data_queue_6__0__5_, 
        data_queue_6__0__4_, data_queue_6__0__3_, data_queue_6__0__2_, 
        data_queue_6__0__1_, data_queue_6__0__0_}), .PRODUCT({N6682, N6681, 
        N6680, N6679, N6678, N6677, N6676, N6675, N6674, N6673, N6672, N6671, 
        N6670, N6669, N6668, N6667}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_14 r1029 ( .A({
        weight_queue_6__1__7_, weight_queue_6__1__6_, weight_queue_6__1__5_, 
        weight_queue_6__1__4_, weight_queue_6__1__3_, weight_queue_6__1__2_, 
        weight_queue_6__1__1_, weight_queue_6__1__0_}), .B({
        data_queue_6__1__7_, data_queue_6__1__6_, data_queue_6__1__5_, 
        data_queue_6__1__4_, data_queue_6__1__3_, data_queue_6__1__2_, 
        data_queue_6__1__1_, data_queue_6__1__0_}), .PRODUCT({N6764, N6763, 
        N6762, N6761, N6760, N6759, N6758, N6757, N6756, N6755, N6754, N6753, 
        N6752, N6751, N6750, N6749}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_13 r1031 ( .A({
        weight_queue_6__2__7_, weight_queue_6__2__6_, weight_queue_6__2__5_, 
        weight_queue_6__2__4_, weight_queue_6__2__3_, weight_queue_6__2__2_, 
        weight_queue_6__2__1_, weight_queue_6__2__0_}), .B({
        data_queue_6__2__7_, data_queue_6__2__6_, data_queue_6__2__5_, 
        data_queue_6__2__4_, data_queue_6__2__3_, data_queue_6__2__2_, 
        data_queue_6__2__1_, data_queue_6__2__0_}), .PRODUCT({N6856, N6855, 
        N6854, N6853, N6852, N6851, N6850, N6849, N6848, N6847, N6846, N6845, 
        N6844, N6843, N6842, N6841}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_12 r1033 ( .A({
        weight_queue_6__3__7_, weight_queue_6__3__6_, weight_queue_6__3__5_, 
        weight_queue_6__3__4_, weight_queue_6__3__3_, weight_queue_6__3__2_, 
        weight_queue_6__3__1_, weight_queue_6__3__0_}), .B({
        data_queue_6__3__7_, data_queue_6__3__6_, data_queue_6__3__5_, 
        data_queue_6__3__4_, data_queue_6__3__3_, data_queue_6__3__2_, 
        data_queue_6__3__1_, data_queue_6__3__0_}), .PRODUCT({N6938, N6937, 
        N6936, N6935, N6934, N6933, N6932, N6931, N6930, N6929, N6928, N6927, 
        N6926, N6925, N6924, N6923}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_11 r1035 ( .A({
        weight_queue_6__4__7_, weight_queue_6__4__6_, weight_queue_6__4__5_, 
        weight_queue_6__4__4_, weight_queue_6__4__3_, weight_queue_6__4__2_, 
        weight_queue_6__4__1_, weight_queue_6__4__0_}), .B({
        data_queue_6__4__7_, data_queue_6__4__6_, data_queue_6__4__5_, 
        data_queue_6__4__4_, data_queue_6__4__3_, data_queue_6__4__2_, 
        data_queue_6__4__1_, data_queue_6__4__0_}), .PRODUCT({N7030, N7029, 
        N7028, N7027, N7026, N7025, N7024, N7023, N7022, N7021, N7020, N7019, 
        N7018, N7017, N7016, N7015}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_10 r1037 ( .A({
        weight_queue_6__5__7_, weight_queue_6__5__6_, weight_queue_6__5__5_, 
        weight_queue_6__5__4_, weight_queue_6__5__3_, weight_queue_6__5__2_, 
        weight_queue_6__5__1_, weight_queue_6__5__0_}), .B({
        data_queue_6__5__7_, data_queue_6__5__6_, data_queue_6__5__5_, 
        data_queue_6__5__4_, data_queue_6__5__3_, data_queue_6__5__2_, 
        data_queue_6__5__1_, data_queue_6__5__0_}), .PRODUCT({N7112, N7111, 
        N7110, N7109, N7108, N7107, N7106, N7105, N7104, N7103, N7102, N7101, 
        N7100, N7099, N7098, N7097}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_9 r1039 ( .A({
        weight_queue_6__6__7_, weight_queue_6__6__6_, weight_queue_6__6__5_, 
        weight_queue_6__6__4_, weight_queue_6__6__3_, weight_queue_6__6__2_, 
        weight_queue_6__6__1_, weight_queue_6__6__0_}), .B({
        data_queue_6__6__7_, data_queue_6__6__6_, data_queue_6__6__5_, 
        data_queue_6__6__4_, data_queue_6__6__3_, data_queue_6__6__2_, 
        data_queue_6__6__1_, data_queue_6__6__0_}), .PRODUCT({N7204, N7203, 
        N7202, N7201, N7200, N7199, N7198, N7197, N7196, N7195, N7194, N7193, 
        N7192, N7191, N7190, N7189}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_8 r1044 ( .A({
        weight_queue_6__7__7_, weight_queue_6__7__6_, weight_queue_6__7__5_, 
        weight_queue_6__7__4_, weight_queue_6__7__3_, weight_queue_6__7__2_, 
        weight_queue_6__7__1_, weight_queue_6__7__0_}), .B({n19606, n19603, 
        n19600, n19597, n19594, n19591, n19588, n19585}), .PRODUCT({N7286, 
        N7285, N7284, N7283, N7282, N7281, N7280, N7279, N7278, N7277, N7276, 
        N7275, N7274, N7273, N7272, N7271}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_7 r1046 ( .A({
        n19557, n19555, n19552, n19549, n19546, n19543, n19540, n19537}), .B({
        data_queue_7__0__7_, data_queue_7__0__6_, data_queue_7__0__5_, 
        data_queue_7__0__4_, data_queue_7__0__3_, data_queue_7__0__2_, 
        data_queue_7__0__1_, data_queue_7__0__0_}), .PRODUCT({N7375, N7374, 
        N7373, N7372, N7371, N7370, N7369, N7368, N7367, N7366, N7365, N7364, 
        N7363, N7362, N7361, N7360}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_6 r1048 ( .A({
        n19533, n19531, n19528, n19525, n19522, n19519, n19516, n19513}), .B({
        data_queue_7__1__7_, data_queue_7__1__6_, data_queue_7__1__5_, 
        data_queue_7__1__4_, data_queue_7__1__3_, data_queue_7__1__2_, 
        data_queue_7__1__1_, data_queue_7__1__0_}), .PRODUCT({N7454, N7453, 
        N7452, N7451, N7450, N7449, N7448, N7447, N7446, N7445, N7444, N7443, 
        N7442, N7441, N7440, N7439}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_5 r1050 ( .A({
        n19509, n19507, n19504, n19501, n19498, n19495, n19492, n19489}), .B({
        data_queue_7__2__7_, data_queue_7__2__6_, data_queue_7__2__5_, 
        data_queue_7__2__4_, data_queue_7__2__3_, data_queue_7__2__2_, 
        data_queue_7__2__1_, data_queue_7__2__0_}), .PRODUCT({N7543, N7542, 
        N7541, N7540, N7539, N7538, N7537, N7536, N7535, N7534, N7533, N7532, 
        N7531, N7530, N7529, N7528}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_4 r1052 ( .A({
        n19485, n19483, n19480, n19477, n19474, n19471, n19468, n19465}), .B({
        data_queue_7__3__7_, data_queue_7__3__6_, data_queue_7__3__5_, 
        data_queue_7__3__4_, data_queue_7__3__3_, data_queue_7__3__2_, 
        data_queue_7__3__1_, data_queue_7__3__0_}), .PRODUCT({N7622, N7621, 
        N7620, N7619, N7618, N7617, N7616, N7615, N7614, N7613, N7612, N7611, 
        N7610, N7609, N7608, N7607}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_3 r1054 ( .A({
        n19461, n19459, n19456, n19453, n19450, n19447, n19444, n19441}), .B({
        data_queue_7__4__7_, data_queue_7__4__6_, data_queue_7__4__5_, 
        data_queue_7__4__4_, data_queue_7__4__3_, data_queue_7__4__2_, 
        data_queue_7__4__1_, data_queue_7__4__0_}), .PRODUCT({N7711, N7710, 
        N7709, N7708, N7707, N7706, N7705, N7704, N7703, N7702, N7701, N7700, 
        N7699, N7698, N7697, N7696}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_2 r1056 ( .A({
        n19437, n19435, n19432, n19429, n19426, n19423, n19420, n19417}), .B({
        data_queue_7__5__7_, data_queue_7__5__6_, data_queue_7__5__5_, 
        data_queue_7__5__4_, data_queue_7__5__3_, data_queue_7__5__2_, 
        data_queue_7__5__1_, data_queue_7__5__0_}), .PRODUCT({N7790, N7789, 
        N7788, N7787, N7786, N7785, N7784, N7783, N7782, N7781, N7780, N7779, 
        N7778, N7777, N7776, N7775}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_1 r1058 ( .A({
        n19413, n19411, n19408, n19405, n19402, n19399, n19396, n19393}), .B({
        data_queue_7__6__7_, data_queue_7__6__6_, data_queue_7__6__5_, 
        data_queue_7__6__4_, data_queue_7__6__3_, data_queue_7__6__2_, 
        data_queue_7__6__1_, data_queue_7__6__0_}), .PRODUCT({N7879, N7878, 
        N7877, N7876, N7875, N7874, N7873, N7872, N7871, N7870, N7869, N7868, 
        N7867, N7866, N7865, N7864}) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_DW02_mult_0 r1063 ( .A({
        n19389, n19387, n19384, n19381, n19378, n19375, n19372, n19369}), .B({
        n19582, n19579, n19576, n19573, n19570, n19567, n19564, n19561}), 
        .PRODUCT({N7961, N7960, N7959, N7958, N7957, N7956, N7955, N7954, 
        N7953, N7952, N7951, N7950, N7949, N7948, N7947, N7946}) );
  DFF_X1 matrix_mul_2D_reg_7__7__8_ ( .D(n17058), .CK(clk), .Q(
        matrix_mul_2D_7__7__8_), .QN(n2874) );
  DFF_X1 matrix_mul_2D_reg_7__7__7_ ( .D(n17063), .CK(clk), .Q(
        matrix_mul_2D_7__7__7_), .QN(n2875) );
  DFF_X1 matrix_mul_2D_reg_7__7__6_ ( .D(n17043), .CK(clk), .Q(
        matrix_mul_2D_7__7__6_), .QN(n2876) );
  DFF_X1 matrix_mul_2D_reg_7__7__5_ ( .D(n17048), .CK(clk), .Q(
        matrix_mul_2D_7__7__5_), .QN(n2877) );
  DFF_X1 matrix_mul_2D_reg_7__7__4_ ( .D(n17053), .CK(clk), .Q(
        matrix_mul_2D_7__7__4_), .QN(n2878) );
  DFF_X1 matrix_mul_2D_reg_7__7__3_ ( .D(n17028), .CK(clk), .Q(
        matrix_mul_2D_7__7__3_), .QN(n2879) );
  DFF_X1 matrix_mul_2D_reg_7__7__2_ ( .D(n17033), .CK(clk), .Q(
        matrix_mul_2D_7__7__2_), .QN(n2880) );
  DFF_X1 matrix_mul_2D_reg_7__7__1_ ( .D(n17038), .CK(clk), .Q(
        matrix_mul_2D_7__7__1_), .QN(n2881) );
  DFF_X1 matrix_mul_2D_reg_7__7__0_ ( .D(n17014), .CK(clk), .Q(
        matrix_mul_2D_7__7__0_), .QN(n2882) );
  DFF_X1 matrix_mul_2D_reg_7__7__14_ ( .D(n17018), .CK(clk), .Q(
        matrix_mul_2D_7__7__14_), .QN(n28680) );
  DFF_X1 matrix_mul_2D_reg_7__7__13_ ( .D(n17023), .CK(clk), .Q(
        matrix_mul_2D_7__7__13_), .QN(n2869) );
  DFF_X1 matrix_mul_2D_reg_7__7__12_ ( .D(n17009), .CK(clk), .Q(
        matrix_mul_2D_7__7__12_), .QN(n2870) );
  DFF_X1 matrix_mul_2D_reg_7__7__11_ ( .D(n16792), .CK(clk), .Q(
        matrix_mul_2D_7__7__11_), .QN(n2871) );
  DFF_X1 matrix_mul_2D_reg_7__7__10_ ( .D(n16777), .CK(clk), .Q(
        matrix_mul_2D_7__7__10_), .QN(n2872) );
  DFF_X1 matrix_mul_2D_reg_7__7__9_ ( .D(n16782), .CK(clk), .Q(
        matrix_mul_2D_7__7__9_), .QN(n2873) );
  DFF_X1 matrix_mul_2D_reg_0__0__14_ ( .D(n16797), .CK(clk), .Q(
        matrix_mul_2D_0__0__14_), .QN(n1845) );
  DFF_X1 matrix_mul_2D_reg_0__0__13_ ( .D(n16802), .CK(clk), .Q(
        matrix_mul_2D_0__0__13_), .QN(n1846) );
  DFF_X1 matrix_mul_2D_reg_0__0__12_ ( .D(n16787), .CK(clk), .Q(
        matrix_mul_2D_0__0__12_), .QN(n1847) );
  DFF_X1 matrix_mul_2D_reg_0__0__11_ ( .D(n16812), .CK(clk), .Q(
        matrix_mul_2D_0__0__11_), .QN(n1848) );
  DFF_X1 matrix_mul_2D_reg_0__0__10_ ( .D(n16807), .CK(clk), .Q(
        matrix_mul_2D_0__0__10_), .QN(n1849) );
  DFF_X1 matrix_mul_2D_reg_0__0__9_ ( .D(n16827), .CK(clk), .Q(
        matrix_mul_2D_0__0__9_), .QN(n1850) );
  DFF_X1 matrix_mul_2D_reg_0__0__8_ ( .D(n16822), .CK(clk), .Q(
        matrix_mul_2D_0__0__8_), .QN(n1851) );
  DFF_X1 matrix_mul_2D_reg_0__0__7_ ( .D(n16817), .CK(clk), .Q(
        matrix_mul_2D_0__0__7_), .QN(n1852) );
  DFF_X1 matrix_mul_2D_reg_0__0__6_ ( .D(n16842), .CK(clk), .Q(
        matrix_mul_2D_0__0__6_), .QN(n1853) );
  DFF_X1 matrix_mul_2D_reg_0__0__5_ ( .D(n16847), .CK(clk), .Q(
        matrix_mul_2D_0__0__5_), .QN(n1854) );
  DFF_X1 matrix_mul_2D_reg_0__0__4_ ( .D(n16832), .CK(clk), .Q(
        matrix_mul_2D_0__0__4_), .QN(n1855) );
  DFF_X1 matrix_mul_2D_reg_0__0__3_ ( .D(n16857), .CK(clk), .Q(
        matrix_mul_2D_0__0__3_), .QN(n1856) );
  DFF_X1 matrix_mul_2D_reg_0__0__2_ ( .D(n16862), .CK(clk), .Q(
        matrix_mul_2D_0__0__2_), .QN(n1857) );
  DFF_X1 matrix_mul_2D_reg_0__0__1_ ( .D(n16837), .CK(clk), .Q(
        matrix_mul_2D_0__0__1_), .QN(n1858) );
  DFF_X1 matrix_mul_2D_reg_0__0__0_ ( .D(n16872), .CK(clk), .Q(
        matrix_mul_2D_0__0__0_), .QN(n1859) );
  DFF_X1 matrix_mul_2D_reg_7__6__7_ ( .D(n16876), .CK(clk), .Q(
        matrix_mul_2D_7__6__7_), .QN(n28600) );
  DFF_X1 matrix_mul_2D_reg_7__6__6_ ( .D(n16852), .CK(clk), .Q(
        matrix_mul_2D_7__6__6_), .QN(n28610) );
  DFF_X1 matrix_mul_2D_reg_7__6__2_ ( .D(n16885), .CK(clk), .Q(
        matrix_mul_2D_7__6__2_), .QN(n28650) );
  DFF_X1 matrix_mul_2D_reg_6__7__5_ ( .D(n16890), .CK(clk), .Q(
        matrix_mul_2D_6__7__5_), .QN(n274500) );
  DFF_X1 matrix_mul_2D_reg_6__7__3_ ( .D(n16867), .CK(clk), .Q(
        matrix_mul_2D_6__7__3_), .QN(n274700) );
  DFF_X1 matrix_mul_2D_reg_7__6__5_ ( .D(n16900), .CK(clk), .Q(
        matrix_mul_2D_7__6__5_), .QN(n28620) );
  DFF_X1 matrix_mul_2D_reg_6__7__2_ ( .D(n16905), .CK(clk), .Q(
        matrix_mul_2D_6__7__2_), .QN(n274800) );
  DFF_X1 matrix_mul_2D_reg_6__7__0_ ( .D(n16881), .CK(clk), .Q(
        matrix_mul_2D_6__7__0_), .QN(n2750) );
  DFF_X1 matrix_mul_2D_reg_6__7__8_ ( .D(n16915), .CK(clk), .Q(
        matrix_mul_2D_6__7__8_), .QN(n274200) );
  DFF_X1 matrix_mul_2D_reg_7__6__14_ ( .D(n16920), .CK(clk), .Q(
        matrix_mul_2D_7__6__14_), .QN(n28530) );
  DFF_X1 matrix_mul_2D_reg_7__6__9_ ( .D(n16895), .CK(clk), .Q(
        matrix_mul_2D_7__6__9_), .QN(n28580) );
  DFF_X1 matrix_mul_2D_reg_7__6__1_ ( .D(n16930), .CK(clk), .Q(
        matrix_mul_2D_7__6__1_), .QN(n28660) );
  DFF_X1 matrix_mul_2D_reg_6__7__12_ ( .D(n16935), .CK(clk), .Q(
        matrix_mul_2D_6__7__12_), .QN(n273800) );
  DFF_X1 matrix_mul_2D_reg_6__7__11_ ( .D(n16910), .CK(clk), .Q(
        matrix_mul_2D_6__7__11_), .QN(n273900) );
  DFF_X1 matrix_mul_2D_reg_7__6__8_ ( .D(n16945), .CK(clk), .Q(
        matrix_mul_2D_7__6__8_), .QN(n28590) );
  DFF_X1 matrix_mul_2D_reg_6__7__9_ ( .D(n16950), .CK(clk), .Q(
        matrix_mul_2D_6__7__9_), .QN(n274100) );
  DFF_X1 matrix_mul_2D_reg_6__7__1_ ( .D(n16925), .CK(clk), .Q(
        matrix_mul_2D_6__7__1_), .QN(n2749) );
  DFF_X1 matrix_mul_2D_reg_7__6__4_ ( .D(n16959), .CK(clk), .Q(
        matrix_mul_2D_7__6__4_), .QN(n28630) );
  DFF_X1 matrix_mul_2D_reg_6__7__7_ ( .D(n16964), .CK(clk), .Q(
        matrix_mul_2D_6__7__7_), .QN(n274300) );
  DFF_X1 matrix_mul_2D_reg_7__6__3_ ( .D(n16940), .CK(clk), .Q(
        matrix_mul_2D_7__6__3_), .QN(n28640) );
  DFF_X1 matrix_mul_2D_reg_6__7__6_ ( .D(n16974), .CK(clk), .Q(
        matrix_mul_2D_6__7__6_), .QN(n274400) );
  DFF_X1 matrix_mul_2D_reg_6__7__4_ ( .D(n16979), .CK(clk), .Q(
        matrix_mul_2D_6__7__4_), .QN(n274600) );
  DFF_X1 matrix_mul_2D_reg_7__6__0_ ( .D(n16955), .CK(clk), .Q(
        matrix_mul_2D_7__6__0_), .QN(n28670) );
  DFF_X1 matrix_mul_2D_reg_7__6__13_ ( .D(n16989), .CK(clk), .Q(
        matrix_mul_2D_7__6__13_), .QN(n28540) );
  DFF_X1 matrix_mul_2D_reg_7__6__11_ ( .D(n16994), .CK(clk), .Q(
        matrix_mul_2D_7__6__11_), .QN(n28560) );
  DFF_X1 matrix_mul_2D_reg_6__7__14_ ( .D(n16969), .CK(clk), .Q(
        matrix_mul_2D_6__7__14_), .QN(n273600) );
  DFF_X1 matrix_mul_2D_reg_6__7__10_ ( .D(n16999), .CK(clk), .Q(
        matrix_mul_2D_6__7__10_), .QN(n274000) );
  DFF_X1 matrix_mul_2D_reg_7__6__12_ ( .D(n17004), .CK(clk), .Q(
        matrix_mul_2D_7__6__12_), .QN(n28550) );
  DFF_X1 matrix_mul_2D_reg_7__6__10_ ( .D(n16984), .CK(clk), .Q(
        matrix_mul_2D_7__6__10_), .QN(n28570) );
  BUF_X1 U3 ( .A(n18863), .Z(n1) );
  BUF_X1 U4 ( .A(n18862), .Z(n2) );
  BUF_X1 U5 ( .A(n24374), .Z(n67) );
  BUF_X1 U6 ( .A(n18678), .Z(n68) );
  BUF_X1 U7 ( .A(n18667), .Z(n69) );
  BUF_X1 U8 ( .A(n18666), .Z(n70) );
  BUF_X1 U9 ( .A(n24129), .Z(n71) );
  BUF_X1 U10 ( .A(n24135), .Z(n72) );
  BUF_X1 U11 ( .A(n20684), .Z(n73) );
  BUF_X1 U12 ( .A(n20676), .Z(n74) );
  BUF_X1 U13 ( .A(n24850), .Z(n75) );
  BUF_X1 U14 ( .A(n20668), .Z(n76) );
  BUF_X1 U15 ( .A(n20667), .Z(n77) );
  BUF_X1 U16 ( .A(n20659), .Z(n78) );
  BUF_X1 U17 ( .A(n20652), .Z(n79) );
  BUF_X1 U18 ( .A(n26812), .Z(n80) );
  BUF_X1 U19 ( .A(n26811), .Z(n81) );
  BUF_X1 U20 ( .A(n26816), .Z(n82) );
  BUF_X1 U21 ( .A(n26815), .Z(n83) );
  BUF_X1 U22 ( .A(n268201), .Z(n84) );
  BUF_X1 U23 ( .A(n26819), .Z(n85) );
  BUF_X1 U24 ( .A(n26824), .Z(n86) );
  BUF_X1 U25 ( .A(n26823), .Z(n87) );
  BUF_X1 U26 ( .A(n26828), .Z(n88) );
  BUF_X1 U27 ( .A(n26827), .Z(n89) );
  BUF_X1 U28 ( .A(n26832), .Z(n90) );
  BUF_X1 U29 ( .A(n26831), .Z(n91) );
  BUF_X1 U30 ( .A(n26836), .Z(n92) );
  BUF_X1 U31 ( .A(n26835), .Z(n93) );
  BUF_X1 U32 ( .A(n268401), .Z(n94) );
  BUF_X1 U33 ( .A(n26839), .Z(n95) );
  BUF_X1 U34 ( .A(n26857), .Z(n96) );
  BUF_X1 U35 ( .A(n26858), .Z(n97) );
  BUF_X1 U36 ( .A(n26865), .Z(n98) );
  BUF_X1 U37 ( .A(n26888), .Z(n99) );
  BUF_X1 U38 ( .A(n26896), .Z(n100) );
  BUF_X1 U39 ( .A(n26892), .Z(n101) );
  BUF_X1 U40 ( .A(n269001), .Z(n102) );
  BUF_X1 U41 ( .A(n23960), .Z(n103) );
  BUF_X1 U42 ( .A(n23929), .Z(n104) );
  BUF_X1 U43 ( .A(n23930), .Z(n105) );
  BUF_X1 U44 ( .A(n23923), .Z(n106) );
  BUF_X1 U45 ( .A(n23924), .Z(n107) );
  BUF_X1 U46 ( .A(n23917), .Z(n108) );
  BUF_X1 U47 ( .A(n23918), .Z(n109) );
  BUF_X1 U48 ( .A(n23911), .Z(n110) );
  BUF_X1 U49 ( .A(n23912), .Z(n111) );
  BUF_X1 U50 ( .A(n23905), .Z(n112) );
  BUF_X1 U51 ( .A(n23906), .Z(n113) );
  BUF_X1 U52 ( .A(n23899), .Z(n114) );
  BUF_X1 U53 ( .A(n23900), .Z(n115) );
  BUF_X1 U54 ( .A(n23893), .Z(n116) );
  BUF_X1 U55 ( .A(n23894), .Z(n117) );
  BUF_X1 U56 ( .A(n23888), .Z(n118) );
  BUF_X1 U57 ( .A(n23887), .Z(n119) );
  BUF_X1 U58 ( .A(n23881), .Z(n120) );
  BUF_X1 U59 ( .A(n23882), .Z(n121) );
  BUF_X1 U60 ( .A(n23875), .Z(n122) );
  BUF_X1 U61 ( .A(n23876), .Z(n123) );
  BUF_X1 U62 ( .A(n23869), .Z(n124) );
  BUF_X1 U63 ( .A(n23870), .Z(n125) );
  BUF_X1 U64 ( .A(n23863), .Z(n126) );
  BUF_X1 U65 ( .A(n23864), .Z(n127) );
  BUF_X1 U66 ( .A(n23857), .Z(n128) );
  BUF_X1 U67 ( .A(n23858), .Z(n129) );
  BUF_X1 U68 ( .A(n23851), .Z(n130) );
  BUF_X1 U69 ( .A(n23852), .Z(n131) );
  BUF_X1 U70 ( .A(n23845), .Z(n132) );
  BUF_X1 U71 ( .A(n23846), .Z(n133) );
  BUF_X1 U72 ( .A(n23840), .Z(n134) );
  BUF_X1 U73 ( .A(n23839), .Z(n135) );
  BUF_X1 U74 ( .A(n23834), .Z(n136) );
  BUF_X1 U75 ( .A(n23833), .Z(n137) );
  BUF_X1 U76 ( .A(n23827), .Z(n138) );
  BUF_X1 U77 ( .A(n23828), .Z(n139) );
  BUF_X1 U78 ( .A(n23822), .Z(n140) );
  BUF_X1 U79 ( .A(n23821), .Z(n141) );
  BUF_X1 U80 ( .A(n23815), .Z(n142) );
  BUF_X1 U81 ( .A(n23816), .Z(n143) );
  BUF_X1 U82 ( .A(n23809), .Z(n144) );
  BUF_X1 U83 ( .A(n23810), .Z(n145) );
  BUF_X1 U84 ( .A(n23803), .Z(n146) );
  BUF_X1 U85 ( .A(n23804), .Z(n147) );
  BUF_X1 U86 ( .A(n23798), .Z(n148) );
  BUF_X1 U87 ( .A(n23797), .Z(n149) );
  BUF_X1 U88 ( .A(n23791), .Z(n150) );
  BUF_X1 U89 ( .A(n23792), .Z(n151) );
  BUF_X1 U90 ( .A(n23785), .Z(n152) );
  BUF_X1 U91 ( .A(n23786), .Z(n153) );
  BUF_X1 U92 ( .A(n23780), .Z(n154) );
  BUF_X1 U93 ( .A(n23779), .Z(n155) );
  BUF_X1 U94 ( .A(n23774), .Z(n156) );
  BUF_X1 U95 ( .A(n23773), .Z(n157) );
  BUF_X1 U96 ( .A(n23767), .Z(n158) );
  BUF_X1 U97 ( .A(n23768), .Z(n159) );
  BUF_X1 U98 ( .A(n23761), .Z(n160) );
  BUF_X1 U99 ( .A(n23762), .Z(n161) );
  BUF_X1 U100 ( .A(n23755), .Z(n162) );
  BUF_X1 U101 ( .A(n23756), .Z(n163) );
  BUF_X1 U102 ( .A(n23750), .Z(n164) );
  BUF_X1 U103 ( .A(n23749), .Z(n165) );
  BUF_X1 U104 ( .A(n23743), .Z(n166) );
  BUF_X1 U105 ( .A(n23744), .Z(n167) );
  BUF_X1 U106 ( .A(n23635), .Z(n168) );
  BUF_X1 U107 ( .A(n23636), .Z(n169) );
  BUF_X1 U108 ( .A(n23635), .Z(n170) );
  BUF_X1 U109 ( .A(n23633), .Z(n171) );
  BUF_X1 U110 ( .A(n23634), .Z(n172) );
  BUF_X1 U111 ( .A(n23633), .Z(n173) );
  BUF_X1 U112 ( .A(n23631), .Z(n174) );
  BUF_X1 U113 ( .A(n23632), .Z(n175) );
  BUF_X1 U114 ( .A(n23631), .Z(n176) );
  BUF_X1 U115 ( .A(n23629), .Z(n177) );
  BUF_X1 U116 ( .A(n23629), .Z(n178) );
  BUF_X1 U117 ( .A(n23630), .Z(n179) );
  BUF_X1 U118 ( .A(n23627), .Z(n180) );
  BUF_X1 U119 ( .A(n23628), .Z(n181) );
  BUF_X1 U120 ( .A(n23627), .Z(n182) );
  BUF_X1 U121 ( .A(n23625), .Z(n183) );
  BUF_X1 U122 ( .A(n23626), .Z(n184) );
  BUF_X1 U123 ( .A(n23625), .Z(n185) );
  BUF_X1 U124 ( .A(n23623), .Z(n186) );
  BUF_X1 U125 ( .A(n23624), .Z(n187) );
  BUF_X1 U126 ( .A(n23623), .Z(n188) );
  BUF_X1 U127 ( .A(n23621), .Z(n189) );
  BUF_X1 U128 ( .A(n23621), .Z(n190) );
  BUF_X1 U129 ( .A(n23622), .Z(n191) );
  BUF_X1 U130 ( .A(n23619), .Z(n192) );
  BUF_X1 U131 ( .A(n23620), .Z(n193) );
  BUF_X1 U132 ( .A(n23619), .Z(n194) );
  BUF_X1 U133 ( .A(n23617), .Z(n195) );
  BUF_X1 U134 ( .A(n23618), .Z(n196) );
  BUF_X1 U135 ( .A(n23617), .Z(n197) );
  BUF_X1 U200 ( .A(n23615), .Z(n198) );
  BUF_X1 U201 ( .A(n23616), .Z(n199) );
  BUF_X1 U202 ( .A(n23615), .Z(n200) );
  BUF_X1 U203 ( .A(n23613), .Z(n201) );
  BUF_X1 U204 ( .A(n23613), .Z(n202) );
  BUF_X1 U205 ( .A(n23614), .Z(n203) );
  BUF_X1 U206 ( .A(n23611), .Z(n204) );
  BUF_X1 U207 ( .A(n23612), .Z(n205) );
  BUF_X1 U208 ( .A(n23611), .Z(n206) );
  BUF_X1 U209 ( .A(n23609), .Z(n207) );
  BUF_X1 U210 ( .A(n23610), .Z(n208) );
  BUF_X1 U211 ( .A(n23609), .Z(n209) );
  BUF_X1 U212 ( .A(n23607), .Z(n210) );
  BUF_X1 U213 ( .A(n23608), .Z(n211) );
  BUF_X1 U214 ( .A(n23607), .Z(n212) );
  BUF_X1 U215 ( .A(n23605), .Z(n213) );
  BUF_X1 U216 ( .A(n23605), .Z(n214) );
  BUF_X1 U217 ( .A(n23606), .Z(n215) );
  BUF_X1 U218 ( .A(n23588), .Z(n216) );
  BUF_X1 U219 ( .A(n23580), .Z(n217) );
  BUF_X1 U220 ( .A(n23580), .Z(n218) );
  BUF_X1 U221 ( .A(n23581), .Z(n219) );
  BUF_X1 U222 ( .A(n23578), .Z(n220) );
  BUF_X1 U223 ( .A(n23579), .Z(n221) );
  BUF_X1 U224 ( .A(n23578), .Z(n222) );
  BUF_X1 U225 ( .A(n23577), .Z(n223) );
  BUF_X1 U226 ( .A(n23576), .Z(n224) );
  BUF_X1 U227 ( .A(n23576), .Z(n225) );
  BUF_X1 U228 ( .A(n23574), .Z(n226) );
  BUF_X1 U229 ( .A(n23575), .Z(n227) );
  BUF_X1 U230 ( .A(n23574), .Z(n228) );
  BUF_X1 U231 ( .A(n23572), .Z(n229) );
  BUF_X1 U232 ( .A(n23573), .Z(n230) );
  BUF_X1 U233 ( .A(n23572), .Z(n231) );
  BUF_X1 U234 ( .A(n23570), .Z(n232) );
  BUF_X1 U235 ( .A(n23571), .Z(n233) );
  BUF_X1 U236 ( .A(n23570), .Z(n234) );
  BUF_X1 U237 ( .A(n23568), .Z(n235) );
  BUF_X1 U238 ( .A(n23568), .Z(n236) );
  BUF_X1 U239 ( .A(n23569), .Z(n237) );
  BUF_X1 U240 ( .A(n23566), .Z(n238) );
  BUF_X1 U241 ( .A(n23567), .Z(n239) );
  BUF_X1 U242 ( .A(n23566), .Z(n240) );
  BUF_X1 U243 ( .A(n23565), .Z(n241) );
  BUF_X1 U244 ( .A(n23564), .Z(n242) );
  BUF_X1 U245 ( .A(n23564), .Z(n243) );
  BUF_X1 U246 ( .A(n24375), .Z(n244) );
  BUF_X1 U247 ( .A(n23561), .Z(n245) );
  BUF_X1 U248 ( .A(n23561), .Z(n246) );
  BUF_X1 U249 ( .A(n23558), .Z(n247) );
  BUF_X1 U250 ( .A(n23558), .Z(n248) );
  BUF_X1 U251 ( .A(n24376), .Z(n249) );
  BUF_X1 U252 ( .A(n24376), .Z(n250) );
  BUF_X1 U253 ( .A(n23556), .Z(n251) );
  BUF_X1 U254 ( .A(n23556), .Z(n252) );
  BUF_X1 U255 ( .A(n23553), .Z(n253) );
  BUF_X1 U256 ( .A(n23553), .Z(n254) );
  BUF_X1 U257 ( .A(n23551), .Z(n255) );
  BUF_X1 U258 ( .A(n23551), .Z(n256) );
  BUF_X1 U259 ( .A(n23550), .Z(n257) );
  BUF_X1 U260 ( .A(n23550), .Z(n258) );
  BUF_X1 U261 ( .A(n23548), .Z(n259) );
  BUF_X1 U262 ( .A(n23549), .Z(n260) );
  BUF_X1 U263 ( .A(n23548), .Z(n261) );
  BUF_X1 U264 ( .A(n23546), .Z(n262) );
  BUF_X1 U265 ( .A(n23547), .Z(n263) );
  BUF_X1 U266 ( .A(n23546), .Z(n264) );
  BUF_X1 U267 ( .A(n23544), .Z(n265) );
  BUF_X1 U268 ( .A(n23545), .Z(n266) );
  BUF_X1 U269 ( .A(n23544), .Z(n267) );
  BUF_X1 U270 ( .A(n23542), .Z(n268) );
  BUF_X1 U271 ( .A(n23542), .Z(n269) );
  BUF_X1 U272 ( .A(n23543), .Z(n270) );
  BUF_X1 U273 ( .A(n23541), .Z(n271) );
  BUF_X1 U274 ( .A(n23540), .Z(n272) );
  BUF_X1 U275 ( .A(n23540), .Z(n273) );
  BUF_X1 U276 ( .A(n23538), .Z(n274) );
  BUF_X1 U277 ( .A(n23539), .Z(n275) );
  BUF_X1 U278 ( .A(n23538), .Z(n276) );
  BUF_X1 U279 ( .A(n23536), .Z(n277) );
  BUF_X1 U280 ( .A(n23537), .Z(n278) );
  BUF_X1 U281 ( .A(n23536), .Z(n279) );
  BUF_X1 U282 ( .A(n23534), .Z(n280) );
  BUF_X1 U283 ( .A(n23535), .Z(n281) );
  BUF_X1 U284 ( .A(n23534), .Z(n282) );
  BUF_X1 U285 ( .A(n23532), .Z(n283) );
  BUF_X1 U286 ( .A(n23533), .Z(n284) );
  BUF_X1 U287 ( .A(n23532), .Z(n285) );
  BUF_X1 U288 ( .A(n23530), .Z(n286) );
  BUF_X1 U289 ( .A(n23530), .Z(n287) );
  BUF_X1 U290 ( .A(n23531), .Z(n288) );
  BUF_X1 U291 ( .A(n23529), .Z(n289) );
  BUF_X1 U292 ( .A(n23528), .Z(n290) );
  BUF_X1 U293 ( .A(n23528), .Z(n291) );
  BUF_X1 U294 ( .A(n23526), .Z(n292) );
  BUF_X1 U295 ( .A(n23527), .Z(n293) );
  BUF_X1 U296 ( .A(n23526), .Z(n294) );
  BUF_X1 U297 ( .A(n23524), .Z(n295) );
  BUF_X1 U298 ( .A(n23525), .Z(n296) );
  BUF_X1 U299 ( .A(n23524), .Z(n297) );
  BUF_X1 U300 ( .A(n23522), .Z(n298) );
  BUF_X1 U301 ( .A(n23523), .Z(n299) );
  BUF_X1 U302 ( .A(n23522), .Z(n300) );
  BUF_X1 U303 ( .A(n23520), .Z(n301) );
  BUF_X1 U304 ( .A(n23521), .Z(n302) );
  BUF_X1 U305 ( .A(n23520), .Z(n303) );
  BUF_X1 U306 ( .A(n23518), .Z(n304) );
  BUF_X1 U307 ( .A(n23518), .Z(n305) );
  BUF_X1 U308 ( .A(n23519), .Z(n306) );
  BUF_X1 U309 ( .A(n23517), .Z(n307) );
  BUF_X1 U310 ( .A(n23516), .Z(n308) );
  BUF_X1 U311 ( .A(n23516), .Z(n309) );
  BUF_X1 U312 ( .A(n23514), .Z(n310) );
  BUF_X1 U313 ( .A(n23515), .Z(n311) );
  BUF_X1 U314 ( .A(n23514), .Z(n312) );
  BUF_X1 U315 ( .A(n23512), .Z(n313) );
  BUF_X1 U316 ( .A(n23513), .Z(n314) );
  BUF_X1 U317 ( .A(n23512), .Z(n315) );
  BUF_X1 U318 ( .A(n23510), .Z(n316) );
  BUF_X1 U319 ( .A(n23511), .Z(n317) );
  BUF_X1 U320 ( .A(n23510), .Z(n318) );
  BUF_X1 U321 ( .A(n23508), .Z(n319) );
  BUF_X1 U322 ( .A(n23509), .Z(n320) );
  BUF_X1 U323 ( .A(n23508), .Z(n321) );
  BUF_X1 U324 ( .A(n23506), .Z(n322) );
  BUF_X1 U325 ( .A(n23507), .Z(n323) );
  BUF_X1 U326 ( .A(n23506), .Z(n324) );
  BUF_X1 U327 ( .A(n23505), .Z(n325) );
  BUF_X1 U328 ( .A(n23504), .Z(n326) );
  BUF_X1 U329 ( .A(n23504), .Z(n327) );
  BUF_X1 U330 ( .A(n23502), .Z(n328) );
  BUF_X1 U331 ( .A(n23503), .Z(n329) );
  BUF_X1 U332 ( .A(n23502), .Z(n330) );
  BUF_X1 U333 ( .A(n23500), .Z(n331) );
  BUF_X1 U334 ( .A(n23501), .Z(n332) );
  BUF_X1 U335 ( .A(n23500), .Z(n333) );
  BUF_X1 U336 ( .A(n23374), .Z(n334) );
  BUF_X1 U337 ( .A(n23375), .Z(n335) );
  BUF_X1 U338 ( .A(n23372), .Z(n336) );
  BUF_X1 U339 ( .A(n23373), .Z(n337) );
  BUF_X1 U340 ( .A(n23370), .Z(n338) );
  BUF_X1 U341 ( .A(n23371), .Z(n339) );
  BUF_X1 U342 ( .A(n23368), .Z(n340) );
  BUF_X1 U343 ( .A(n23369), .Z(n341) );
  BUF_X1 U344 ( .A(n23366), .Z(n342) );
  BUF_X1 U345 ( .A(n23367), .Z(n343) );
  BUF_X1 U346 ( .A(n23364), .Z(n344) );
  BUF_X1 U347 ( .A(n23365), .Z(n345) );
  BUF_X1 U348 ( .A(n23362), .Z(n346) );
  BUF_X1 U349 ( .A(n23363), .Z(n347) );
  BUF_X1 U350 ( .A(n23360), .Z(n348) );
  BUF_X1 U351 ( .A(n23361), .Z(n349) );
  BUF_X1 U352 ( .A(n23358), .Z(n350) );
  BUF_X1 U353 ( .A(n23359), .Z(n351) );
  BUF_X1 U354 ( .A(n23356), .Z(n352) );
  BUF_X1 U355 ( .A(n23357), .Z(n353) );
  BUF_X1 U356 ( .A(n23354), .Z(n354) );
  BUF_X1 U357 ( .A(n23355), .Z(n355) );
  BUF_X1 U358 ( .A(n23352), .Z(n356) );
  BUF_X1 U359 ( .A(n23353), .Z(n357) );
  BUF_X1 U360 ( .A(n23350), .Z(n358) );
  BUF_X1 U361 ( .A(n23351), .Z(n359) );
  BUF_X1 U362 ( .A(n23348), .Z(n360) );
  BUF_X1 U363 ( .A(n23349), .Z(n361) );
  BUF_X1 U364 ( .A(n23346), .Z(n362) );
  BUF_X1 U365 ( .A(n23347), .Z(n363) );
  BUF_X1 U366 ( .A(n23344), .Z(n364) );
  BUF_X1 U367 ( .A(n23345), .Z(n365) );
  BUF_X1 U368 ( .A(n23330), .Z(n366) );
  BUF_X1 U369 ( .A(n23331), .Z(n367) );
  BUF_X1 U370 ( .A(n23328), .Z(n368) );
  BUF_X1 U371 ( .A(n23329), .Z(n369) );
  BUF_X1 U372 ( .A(n23326), .Z(n370) );
  BUF_X1 U373 ( .A(n23327), .Z(n371) );
  BUF_X1 U374 ( .A(n23324), .Z(n372) );
  BUF_X1 U375 ( .A(n23325), .Z(n373) );
  BUF_X1 U376 ( .A(n23322), .Z(n374) );
  BUF_X1 U377 ( .A(n23323), .Z(n375) );
  BUF_X1 U378 ( .A(n23320), .Z(n376) );
  BUF_X1 U379 ( .A(n23321), .Z(n377) );
  BUF_X1 U380 ( .A(n23318), .Z(n378) );
  BUF_X1 U381 ( .A(n23319), .Z(n379) );
  BUF_X1 U382 ( .A(n23316), .Z(n380) );
  BUF_X1 U383 ( .A(n23317), .Z(n381) );
  BUF_X1 U384 ( .A(n23314), .Z(n382) );
  BUF_X1 U385 ( .A(n23315), .Z(n383) );
  BUF_X1 U386 ( .A(n23312), .Z(n384) );
  BUF_X1 U387 ( .A(n23313), .Z(n385) );
  BUF_X1 U388 ( .A(n23310), .Z(n386) );
  BUF_X1 U389 ( .A(n23311), .Z(n387) );
  BUF_X1 U390 ( .A(n23308), .Z(n388) );
  BUF_X1 U391 ( .A(n23309), .Z(n389) );
  BUF_X1 U392 ( .A(n23306), .Z(n390) );
  BUF_X1 U393 ( .A(n23307), .Z(n391) );
  BUF_X1 U394 ( .A(n23304), .Z(n392) );
  BUF_X1 U395 ( .A(n23305), .Z(n393) );
  BUF_X1 U396 ( .A(n23300), .Z(n394) );
  BUF_X1 U397 ( .A(n26159), .Z(n395) );
  BUF_X1 U398 ( .A(n25062), .Z(n396) );
  BUF_X1 U399 ( .A(n19015), .Z(n397) );
  BUF_X1 U400 ( .A(n19014), .Z(n398) );
  BUF_X1 U401 ( .A(n19013), .Z(n399) );
  BUF_X1 U402 ( .A(n25055), .Z(n400) );
  BUF_X1 U403 ( .A(n25053), .Z(n401) );
  BUF_X1 U404 ( .A(n19012), .Z(n402) );
  BUF_X1 U405 ( .A(n19011), .Z(n403) );
  BUF_X1 U406 ( .A(n19010), .Z(n404) );
  BUF_X1 U407 ( .A(n19009), .Z(n405) );
  BUF_X1 U408 ( .A(n25047), .Z(n406) );
  BUF_X1 U409 ( .A(n25045), .Z(n407) );
  BUF_X1 U410 ( .A(n19008), .Z(n408) );
  BUF_X1 U411 ( .A(n19007), .Z(n409) );
  BUF_X1 U412 ( .A(n19006), .Z(n410) );
  BUF_X1 U413 ( .A(n19005), .Z(n411) );
  BUF_X1 U414 ( .A(n25039), .Z(n412) );
  BUF_X1 U415 ( .A(n25037), .Z(n413) );
  BUF_X1 U416 ( .A(n19004), .Z(n414) );
  BUF_X1 U417 ( .A(n19003), .Z(n415) );
  BUF_X1 U418 ( .A(n19002), .Z(n416) );
  BUF_X1 U419 ( .A(n25030), .Z(n417) );
  BUF_X1 U420 ( .A(n18999), .Z(n418) );
  BUF_X1 U421 ( .A(n18998), .Z(n419) );
  BUF_X1 U422 ( .A(n18997), .Z(n420) );
  BUF_X1 U423 ( .A(n18996), .Z(n421) );
  BUF_X1 U424 ( .A(n18995), .Z(n422) );
  BUF_X1 U425 ( .A(n18994), .Z(n423) );
  BUF_X1 U426 ( .A(n18993), .Z(n424) );
  BUF_X1 U427 ( .A(n18992), .Z(n425) );
  BUF_X1 U428 ( .A(n18991), .Z(n426) );
  BUF_X1 U429 ( .A(n71), .Z(n427) );
  BUF_X1 U430 ( .A(n72), .Z(n428) );
  BUF_X1 U431 ( .A(n73), .Z(n429) );
  BUF_X1 U432 ( .A(n18979), .Z(n430) );
  BUF_X1 U433 ( .A(n18978), .Z(n431) );
  BUF_X1 U434 ( .A(n74), .Z(n432) );
  BUF_X1 U435 ( .A(n75), .Z(n433) );
  BUF_X1 U436 ( .A(n18976), .Z(n434) );
  BUF_X1 U437 ( .A(n76), .Z(n435) );
  BUF_X1 U438 ( .A(n18974), .Z(n436) );
  BUF_X1 U439 ( .A(n77), .Z(n437) );
  BUF_X1 U440 ( .A(n18973), .Z(n438) );
  BUF_X1 U441 ( .A(n18971), .Z(n439) );
  BUF_X1 U442 ( .A(n78), .Z(n440) );
  BUF_X1 U443 ( .A(n79), .Z(n441) );
  BUF_X1 U444 ( .A(n18969), .Z(n442) );
  BUF_X1 U445 ( .A(n18968), .Z(n443) );
  BUF_X1 U446 ( .A(n17091), .Z(n444) );
  BUF_X1 U447 ( .A(n18965), .Z(n445) );
  BUF_X1 U448 ( .A(n17092), .Z(n446) );
  BUF_X1 U449 ( .A(n18963), .Z(n447) );
  BUF_X1 U450 ( .A(n17093), .Z(n448) );
  BUF_X1 U451 ( .A(n18962), .Z(n449) );
  BUF_X1 U452 ( .A(n18960), .Z(n450) );
  BUF_X1 U453 ( .A(n17094), .Z(n451) );
  BUF_X1 U454 ( .A(cycle_num[0]), .Z(n452) );
  BUF_X1 U455 ( .A(cycle_num[6]), .Z(n453) );
  BUF_X1 U456 ( .A(cycle_num[4]), .Z(n454) );
  BUF_X1 U457 ( .A(cycle_num[1]), .Z(n455) );
  BUF_X1 U458 ( .A(n875), .Z(n456) );
  BUF_X1 U459 ( .A(n548), .Z(n457) );
  BUF_X1 U460 ( .A(n545), .Z(n458) );
  BUF_X1 U461 ( .A(n540), .Z(n459) );
  BUF_X1 U462 ( .A(n538), .Z(n460) );
  INV_X1 U463 ( .A(matrix_index[5]), .ZN(n461) );
  INV_X1 U464 ( .A(n461), .ZN(n462) );
  INV_X1 U465 ( .A(n461), .ZN(n463) );
  BUF_X1 U466 ( .A(cycle_num[8]), .Z(n464) );
  BUF_X1 U467 ( .A(cycle_num[8]), .Z(n465) );
  BUF_X1 U468 ( .A(cycle_num[2]), .Z(n466) );
  BUF_X1 U469 ( .A(cycle_num[2]), .Z(n467) );
  BUF_X1 U470 ( .A(matrix_index[0]), .Z(n881) );
  INV_X1 U471 ( .A(n881), .ZN(n468) );
  INV_X1 U472 ( .A(n881), .ZN(n469) );
  INV_X1 U473 ( .A(matrix_index[1]), .ZN(n470) );
  INV_X1 U474 ( .A(n873), .ZN(n471) );
  INV_X1 U475 ( .A(n868), .ZN(n472) );
  INV_X1 U476 ( .A(n863), .ZN(n473) );
  INV_X1 U477 ( .A(n858), .ZN(n474) );
  INV_X1 U478 ( .A(n853), .ZN(n475) );
  INV_X1 U479 ( .A(n848), .ZN(n476) );
  INV_X1 U480 ( .A(n843), .ZN(n477) );
  INV_X1 U481 ( .A(n838), .ZN(n478) );
  INV_X1 U482 ( .A(n833), .ZN(n479) );
  INV_X1 U483 ( .A(n828), .ZN(n480) );
  INV_X1 U484 ( .A(n823), .ZN(n481) );
  INV_X1 U485 ( .A(n818), .ZN(n482) );
  INV_X1 U486 ( .A(n813), .ZN(n483) );
  INV_X1 U487 ( .A(n808), .ZN(n484) );
  INV_X1 U488 ( .A(n803), .ZN(n485) );
  INV_X1 U489 ( .A(n798), .ZN(n486) );
  INV_X1 U490 ( .A(n793), .ZN(n487) );
  INV_X1 U491 ( .A(n788), .ZN(n488) );
  INV_X1 U492 ( .A(n783), .ZN(n489) );
  INV_X1 U493 ( .A(n778), .ZN(n490) );
  INV_X1 U494 ( .A(n773), .ZN(n491) );
  INV_X1 U495 ( .A(n768), .ZN(n492) );
  INV_X1 U496 ( .A(n763), .ZN(n493) );
  INV_X1 U497 ( .A(n758), .ZN(n494) );
  INV_X1 U498 ( .A(n753), .ZN(n495) );
  INV_X1 U499 ( .A(n748), .ZN(n496) );
  INV_X1 U500 ( .A(n743), .ZN(n497) );
  INV_X1 U501 ( .A(n738), .ZN(n498) );
  INV_X1 U502 ( .A(n733), .ZN(n499) );
  INV_X1 U503 ( .A(n728), .ZN(n500) );
  INV_X1 U504 ( .A(n723), .ZN(n501) );
  INV_X1 U505 ( .A(n718), .ZN(n502) );
  INV_X1 U506 ( .A(n713), .ZN(n503) );
  INV_X1 U507 ( .A(n708), .ZN(n504) );
  INV_X1 U508 ( .A(n703), .ZN(n505) );
  INV_X1 U509 ( .A(n698), .ZN(n506) );
  INV_X1 U510 ( .A(n693), .ZN(n507) );
  INV_X1 U511 ( .A(n688), .ZN(n508) );
  INV_X1 U512 ( .A(n683), .ZN(n509) );
  INV_X1 U513 ( .A(n678), .ZN(n510) );
  INV_X1 U514 ( .A(n673), .ZN(n511) );
  INV_X1 U515 ( .A(n668), .ZN(n512) );
  INV_X1 U516 ( .A(n663), .ZN(n513) );
  INV_X1 U517 ( .A(n658), .ZN(n514) );
  INV_X1 U518 ( .A(n653), .ZN(n515) );
  INV_X1 U519 ( .A(n648), .ZN(n516) );
  INV_X1 U520 ( .A(n643), .ZN(n517) );
  INV_X1 U521 ( .A(n638), .ZN(n518) );
  INV_X1 U522 ( .A(n633), .ZN(n519) );
  INV_X1 U523 ( .A(n628), .ZN(n520) );
  INV_X1 U524 ( .A(n623), .ZN(n521) );
  INV_X1 U525 ( .A(n618), .ZN(n522) );
  INV_X1 U526 ( .A(n613), .ZN(n523) );
  INV_X1 U527 ( .A(n608), .ZN(n524) );
  INV_X1 U528 ( .A(n603), .ZN(n525) );
  INV_X1 U529 ( .A(n598), .ZN(n526) );
  INV_X1 U530 ( .A(n593), .ZN(n527) );
  INV_X1 U531 ( .A(n588), .ZN(n528) );
  INV_X1 U532 ( .A(n583), .ZN(n529) );
  INV_X1 U533 ( .A(n578), .ZN(n530) );
  INV_X1 U534 ( .A(n573), .ZN(n531) );
  INV_X1 U535 ( .A(n568), .ZN(n532) );
  INV_X1 U536 ( .A(n563), .ZN(n533) );
  INV_X1 U537 ( .A(n558), .ZN(n534) );
  INV_X1 U538 ( .A(matrix_index[3]), .ZN(n535) );
  INV_X1 U539 ( .A(n535), .ZN(n536) );
  INV_X1 U540 ( .A(n535), .ZN(n537) );
  BUF_X1 U541 ( .A(cycle_num[7]), .Z(n538) );
  BUF_X1 U542 ( .A(cycle_num[7]), .Z(n539) );
  BUF_X1 U543 ( .A(cycle_num[5]), .Z(n540) );
  BUF_X1 U544 ( .A(cycle_num[5]), .Z(n541) );
  INV_X1 U545 ( .A(n27300), .ZN(n542) );
  INV_X1 U546 ( .A(n27303), .ZN(n543) );
  INV_X1 U547 ( .A(matrix_index[4]), .ZN(n544) );
  INV_X1 U548 ( .A(n544), .ZN(n545) );
  INV_X1 U549 ( .A(n544), .ZN(n546) );
  INV_X1 U550 ( .A(matrix_index[2]), .ZN(n547) );
  INV_X1 U551 ( .A(n547), .ZN(n548) );
  INV_X1 U552 ( .A(n547), .ZN(n549) );
  INV_X1 U553 ( .A(cycle_num[3]), .ZN(n550) );
  INV_X1 U554 ( .A(n27301), .ZN(n551) );
  INV_X1 U555 ( .A(n550), .ZN(n552) );
  INV_X1 U556 ( .A(n550), .ZN(n553) );
  INV_X1 U557 ( .A(N2574), .ZN(n554) );
  INV_X1 U558 ( .A(n554), .ZN(n555) );
  INV_X1 U559 ( .A(n534), .ZN(n556) );
  INV_X1 U560 ( .A(n534), .ZN(n557) );
  INV_X1 U561 ( .A(n554), .ZN(n558) );
  INV_X1 U562 ( .A(N2656), .ZN(n559) );
  INV_X1 U563 ( .A(n559), .ZN(n560) );
  INV_X1 U564 ( .A(n533), .ZN(n561) );
  INV_X1 U565 ( .A(n533), .ZN(n562) );
  INV_X1 U566 ( .A(n559), .ZN(n563) );
  INV_X1 U567 ( .A(N2748), .ZN(n564) );
  INV_X1 U568 ( .A(n564), .ZN(n565) );
  INV_X1 U569 ( .A(n532), .ZN(n566) );
  INV_X1 U570 ( .A(n532), .ZN(n567) );
  INV_X1 U571 ( .A(n564), .ZN(n568) );
  INV_X1 U572 ( .A(N2830), .ZN(n569) );
  INV_X1 U573 ( .A(n569), .ZN(n570) );
  INV_X1 U574 ( .A(n531), .ZN(n571) );
  INV_X1 U575 ( .A(n531), .ZN(n572) );
  INV_X1 U576 ( .A(n569), .ZN(n573) );
  INV_X1 U577 ( .A(N2922), .ZN(n574) );
  INV_X1 U578 ( .A(n574), .ZN(n575) );
  INV_X1 U579 ( .A(n530), .ZN(n576) );
  INV_X1 U580 ( .A(n530), .ZN(n577) );
  INV_X1 U581 ( .A(n574), .ZN(n578) );
  INV_X1 U582 ( .A(N3004), .ZN(n579) );
  INV_X1 U583 ( .A(n579), .ZN(n580) );
  INV_X1 U584 ( .A(n529), .ZN(n581) );
  INV_X1 U585 ( .A(n529), .ZN(n582) );
  INV_X1 U586 ( .A(n579), .ZN(n583) );
  INV_X1 U587 ( .A(N3096), .ZN(n584) );
  INV_X1 U588 ( .A(n584), .ZN(n585) );
  INV_X1 U589 ( .A(n528), .ZN(n586) );
  INV_X1 U590 ( .A(n528), .ZN(n587) );
  INV_X1 U591 ( .A(n584), .ZN(n588) );
  INV_X1 U592 ( .A(N3178), .ZN(n589) );
  INV_X1 U593 ( .A(n589), .ZN(n590) );
  INV_X1 U594 ( .A(n527), .ZN(n591) );
  INV_X1 U595 ( .A(n527), .ZN(n592) );
  INV_X1 U596 ( .A(n589), .ZN(n593) );
  INV_X1 U597 ( .A(N3267), .ZN(n594) );
  INV_X1 U598 ( .A(n594), .ZN(n595) );
  INV_X1 U599 ( .A(n526), .ZN(n596) );
  INV_X1 U600 ( .A(n526), .ZN(n597) );
  INV_X1 U601 ( .A(n594), .ZN(n598) );
  INV_X1 U602 ( .A(N3346), .ZN(n599) );
  INV_X1 U603 ( .A(n599), .ZN(n600) );
  INV_X1 U604 ( .A(n525), .ZN(n601) );
  INV_X1 U605 ( .A(n525), .ZN(n602) );
  INV_X1 U606 ( .A(n599), .ZN(n603) );
  INV_X1 U607 ( .A(N3435), .ZN(n604) );
  INV_X1 U608 ( .A(n604), .ZN(n605) );
  INV_X1 U609 ( .A(n524), .ZN(n606) );
  INV_X1 U610 ( .A(n524), .ZN(n607) );
  INV_X1 U611 ( .A(n604), .ZN(n608) );
  INV_X1 U612 ( .A(N3514), .ZN(n609) );
  INV_X1 U613 ( .A(n609), .ZN(n610) );
  INV_X1 U614 ( .A(n523), .ZN(n611) );
  INV_X1 U615 ( .A(n523), .ZN(n612) );
  INV_X1 U616 ( .A(n609), .ZN(n613) );
  INV_X1 U617 ( .A(N3603), .ZN(n614) );
  INV_X1 U618 ( .A(n614), .ZN(n615) );
  INV_X1 U619 ( .A(n522), .ZN(n616) );
  INV_X1 U620 ( .A(n522), .ZN(n617) );
  INV_X1 U621 ( .A(n614), .ZN(n618) );
  INV_X1 U622 ( .A(N3682), .ZN(n619) );
  INV_X1 U623 ( .A(n619), .ZN(n620) );
  INV_X1 U624 ( .A(n521), .ZN(n621) );
  INV_X1 U625 ( .A(n521), .ZN(n622) );
  INV_X1 U626 ( .A(n619), .ZN(n623) );
  INV_X1 U627 ( .A(N3771), .ZN(n624) );
  INV_X1 U628 ( .A(n624), .ZN(n625) );
  INV_X1 U629 ( .A(n520), .ZN(n626) );
  INV_X1 U630 ( .A(n520), .ZN(n627) );
  INV_X1 U631 ( .A(n624), .ZN(n628) );
  INV_X1 U632 ( .A(N3853), .ZN(n629) );
  INV_X1 U633 ( .A(n629), .ZN(n630) );
  INV_X1 U634 ( .A(n519), .ZN(n631) );
  INV_X1 U635 ( .A(n519), .ZN(n632) );
  INV_X1 U636 ( .A(n629), .ZN(n633) );
  INV_X1 U637 ( .A(N3942), .ZN(n634) );
  INV_X1 U638 ( .A(n634), .ZN(n635) );
  INV_X1 U639 ( .A(n518), .ZN(n636) );
  INV_X1 U640 ( .A(n518), .ZN(n637) );
  INV_X1 U641 ( .A(n634), .ZN(n638) );
  INV_X1 U642 ( .A(N4021), .ZN(n639) );
  INV_X1 U643 ( .A(n639), .ZN(n640) );
  INV_X1 U644 ( .A(n517), .ZN(n641) );
  INV_X1 U645 ( .A(n517), .ZN(n642) );
  INV_X1 U646 ( .A(n639), .ZN(n643) );
  INV_X1 U647 ( .A(N4110), .ZN(n644) );
  INV_X1 U648 ( .A(n644), .ZN(n645) );
  INV_X1 U649 ( .A(n516), .ZN(n646) );
  INV_X1 U650 ( .A(n516), .ZN(n647) );
  INV_X1 U651 ( .A(n644), .ZN(n648) );
  INV_X1 U652 ( .A(N4189), .ZN(n649) );
  INV_X1 U653 ( .A(n649), .ZN(n650) );
  INV_X1 U654 ( .A(n515), .ZN(n651) );
  INV_X1 U655 ( .A(n515), .ZN(n652) );
  INV_X1 U656 ( .A(n649), .ZN(n653) );
  INV_X1 U657 ( .A(N4278), .ZN(n654) );
  INV_X1 U658 ( .A(n654), .ZN(n655) );
  INV_X1 U659 ( .A(n514), .ZN(n656) );
  INV_X1 U660 ( .A(n514), .ZN(n657) );
  INV_X1 U661 ( .A(n654), .ZN(n658) );
  INV_X1 U662 ( .A(N4357), .ZN(n659) );
  INV_X1 U663 ( .A(n659), .ZN(n660) );
  INV_X1 U664 ( .A(n513), .ZN(n661) );
  INV_X1 U665 ( .A(n513), .ZN(n662) );
  INV_X1 U666 ( .A(n659), .ZN(n663) );
  INV_X1 U667 ( .A(N4446), .ZN(n664) );
  INV_X1 U668 ( .A(n664), .ZN(n665) );
  INV_X1 U669 ( .A(n512), .ZN(n666) );
  INV_X1 U670 ( .A(n512), .ZN(n667) );
  INV_X1 U671 ( .A(n664), .ZN(n668) );
  INV_X1 U672 ( .A(N4528), .ZN(n669) );
  INV_X1 U673 ( .A(n669), .ZN(n670) );
  INV_X1 U674 ( .A(n511), .ZN(n671) );
  INV_X1 U675 ( .A(n511), .ZN(n672) );
  INV_X1 U676 ( .A(n669), .ZN(n673) );
  INV_X1 U677 ( .A(N4628), .ZN(n674) );
  INV_X1 U678 ( .A(n674), .ZN(n675) );
  INV_X1 U679 ( .A(n510), .ZN(n676) );
  INV_X1 U680 ( .A(n510), .ZN(n677) );
  INV_X1 U681 ( .A(n674), .ZN(n678) );
  INV_X1 U682 ( .A(N4710), .ZN(n679) );
  INV_X1 U683 ( .A(n679), .ZN(n680) );
  INV_X1 U684 ( .A(n509), .ZN(n681) );
  INV_X1 U685 ( .A(n509), .ZN(n682) );
  INV_X1 U686 ( .A(n679), .ZN(n683) );
  INV_X1 U687 ( .A(N4802), .ZN(n684) );
  INV_X1 U688 ( .A(n684), .ZN(n685) );
  INV_X1 U689 ( .A(n508), .ZN(n686) );
  INV_X1 U690 ( .A(n508), .ZN(n687) );
  INV_X1 U691 ( .A(n684), .ZN(n688) );
  INV_X1 U692 ( .A(N4884), .ZN(n689) );
  INV_X1 U693 ( .A(n689), .ZN(n690) );
  INV_X1 U694 ( .A(n507), .ZN(n691) );
  INV_X1 U695 ( .A(n507), .ZN(n692) );
  INV_X1 U696 ( .A(n689), .ZN(n693) );
  INV_X1 U697 ( .A(N4976), .ZN(n694) );
  INV_X1 U698 ( .A(n694), .ZN(n695) );
  INV_X1 U699 ( .A(n506), .ZN(n696) );
  INV_X1 U700 ( .A(n506), .ZN(n697) );
  INV_X1 U701 ( .A(n694), .ZN(n698) );
  INV_X1 U702 ( .A(N5058), .ZN(n699) );
  INV_X1 U703 ( .A(n699), .ZN(n700) );
  INV_X1 U704 ( .A(n505), .ZN(n701) );
  INV_X1 U705 ( .A(n505), .ZN(n702) );
  INV_X1 U706 ( .A(n699), .ZN(n703) );
  INV_X1 U707 ( .A(N5150), .ZN(n704) );
  INV_X1 U708 ( .A(n704), .ZN(n705) );
  INV_X1 U709 ( .A(n504), .ZN(n706) );
  INV_X1 U710 ( .A(n504), .ZN(n707) );
  INV_X1 U711 ( .A(n704), .ZN(n708) );
  INV_X1 U712 ( .A(N5232), .ZN(n709) );
  INV_X1 U713 ( .A(n709), .ZN(n710) );
  INV_X1 U714 ( .A(n503), .ZN(n711) );
  INV_X1 U715 ( .A(n503), .ZN(n712) );
  INV_X1 U716 ( .A(n709), .ZN(n713) );
  INV_X1 U717 ( .A(N5321), .ZN(n714) );
  INV_X1 U718 ( .A(n714), .ZN(n715) );
  INV_X1 U719 ( .A(n502), .ZN(n716) );
  INV_X1 U720 ( .A(n502), .ZN(n717) );
  INV_X1 U721 ( .A(n714), .ZN(n718) );
  INV_X1 U722 ( .A(N5400), .ZN(n719) );
  INV_X1 U723 ( .A(n719), .ZN(n720) );
  INV_X1 U724 ( .A(n501), .ZN(n721) );
  INV_X1 U725 ( .A(n501), .ZN(n722) );
  INV_X1 U726 ( .A(n719), .ZN(n723) );
  INV_X1 U727 ( .A(N5489), .ZN(n724) );
  INV_X1 U728 ( .A(n724), .ZN(n725) );
  INV_X1 U729 ( .A(n500), .ZN(n726) );
  INV_X1 U730 ( .A(n500), .ZN(n727) );
  INV_X1 U731 ( .A(n724), .ZN(n728) );
  INV_X1 U732 ( .A(N5568), .ZN(n729) );
  INV_X1 U733 ( .A(n729), .ZN(n730) );
  INV_X1 U734 ( .A(n499), .ZN(n731) );
  INV_X1 U735 ( .A(n499), .ZN(n732) );
  INV_X1 U736 ( .A(n729), .ZN(n733) );
  INV_X1 U737 ( .A(N5657), .ZN(n734) );
  INV_X1 U738 ( .A(n734), .ZN(n735) );
  INV_X1 U739 ( .A(n498), .ZN(n736) );
  INV_X1 U740 ( .A(n498), .ZN(n737) );
  INV_X1 U741 ( .A(n734), .ZN(n738) );
  INV_X1 U742 ( .A(N5736), .ZN(n739) );
  INV_X1 U743 ( .A(n739), .ZN(n740) );
  INV_X1 U744 ( .A(n497), .ZN(n741) );
  INV_X1 U745 ( .A(n497), .ZN(n742) );
  INV_X1 U746 ( .A(n739), .ZN(n743) );
  INV_X1 U747 ( .A(N5825), .ZN(n744) );
  INV_X1 U748 ( .A(n744), .ZN(n745) );
  INV_X1 U749 ( .A(n496), .ZN(n746) );
  INV_X1 U750 ( .A(n496), .ZN(n747) );
  INV_X1 U751 ( .A(n744), .ZN(n748) );
  INV_X1 U752 ( .A(N5907), .ZN(n749) );
  INV_X1 U753 ( .A(n749), .ZN(n750) );
  INV_X1 U754 ( .A(n495), .ZN(n751) );
  INV_X1 U755 ( .A(n495), .ZN(n752) );
  INV_X1 U756 ( .A(n749), .ZN(n753) );
  INV_X1 U757 ( .A(N5996), .ZN(n754) );
  INV_X1 U758 ( .A(n754), .ZN(n755) );
  INV_X1 U759 ( .A(n494), .ZN(n756) );
  INV_X1 U760 ( .A(n494), .ZN(n757) );
  INV_X1 U761 ( .A(n754), .ZN(n758) );
  INV_X1 U762 ( .A(N6075), .ZN(n759) );
  INV_X1 U763 ( .A(n759), .ZN(n760) );
  INV_X1 U764 ( .A(n493), .ZN(n761) );
  INV_X1 U765 ( .A(n493), .ZN(n762) );
  INV_X1 U766 ( .A(n759), .ZN(n763) );
  INV_X1 U767 ( .A(N6164), .ZN(n764) );
  INV_X1 U768 ( .A(n764), .ZN(n765) );
  INV_X1 U769 ( .A(n492), .ZN(n766) );
  INV_X1 U770 ( .A(n492), .ZN(n767) );
  INV_X1 U771 ( .A(n764), .ZN(n768) );
  INV_X1 U772 ( .A(N6243), .ZN(n769) );
  INV_X1 U773 ( .A(n769), .ZN(n770) );
  INV_X1 U774 ( .A(n491), .ZN(n771) );
  INV_X1 U775 ( .A(n491), .ZN(n772) );
  INV_X1 U776 ( .A(n769), .ZN(n773) );
  INV_X1 U777 ( .A(N6332), .ZN(n774) );
  INV_X1 U778 ( .A(n774), .ZN(n775) );
  INV_X1 U779 ( .A(n490), .ZN(n776) );
  INV_X1 U780 ( .A(n490), .ZN(n777) );
  INV_X1 U781 ( .A(n774), .ZN(n778) );
  INV_X1 U782 ( .A(N6411), .ZN(n779) );
  INV_X1 U783 ( .A(n779), .ZN(n780) );
  INV_X1 U784 ( .A(n489), .ZN(n781) );
  INV_X1 U785 ( .A(n489), .ZN(n782) );
  INV_X1 U786 ( .A(n779), .ZN(n783) );
  INV_X1 U787 ( .A(N6500), .ZN(n784) );
  INV_X1 U788 ( .A(n784), .ZN(n785) );
  INV_X1 U789 ( .A(n488), .ZN(n786) );
  INV_X1 U790 ( .A(n488), .ZN(n787) );
  INV_X1 U791 ( .A(n784), .ZN(n788) );
  INV_X1 U792 ( .A(N6582), .ZN(n789) );
  INV_X1 U793 ( .A(n789), .ZN(n790) );
  INV_X1 U794 ( .A(n487), .ZN(n791) );
  INV_X1 U795 ( .A(n487), .ZN(n792) );
  INV_X1 U796 ( .A(n789), .ZN(n793) );
  INV_X1 U797 ( .A(N6682), .ZN(n794) );
  INV_X1 U798 ( .A(n794), .ZN(n795) );
  INV_X1 U799 ( .A(n486), .ZN(n796) );
  INV_X1 U800 ( .A(n486), .ZN(n797) );
  INV_X1 U801 ( .A(n794), .ZN(n798) );
  INV_X1 U802 ( .A(N6764), .ZN(n799) );
  INV_X1 U803 ( .A(n799), .ZN(n800) );
  INV_X1 U804 ( .A(n485), .ZN(n801) );
  INV_X1 U805 ( .A(n485), .ZN(n802) );
  INV_X1 U806 ( .A(n799), .ZN(n803) );
  INV_X1 U807 ( .A(N6856), .ZN(n804) );
  INV_X1 U808 ( .A(n804), .ZN(n805) );
  INV_X1 U809 ( .A(n484), .ZN(n806) );
  INV_X1 U810 ( .A(n484), .ZN(n807) );
  INV_X1 U811 ( .A(n804), .ZN(n808) );
  INV_X1 U812 ( .A(N6938), .ZN(n809) );
  INV_X1 U813 ( .A(n809), .ZN(n810) );
  INV_X1 U814 ( .A(n483), .ZN(n811) );
  INV_X1 U815 ( .A(n483), .ZN(n812) );
  INV_X1 U816 ( .A(n809), .ZN(n813) );
  INV_X1 U817 ( .A(N7030), .ZN(n814) );
  INV_X1 U818 ( .A(n814), .ZN(n815) );
  INV_X1 U819 ( .A(n482), .ZN(n816) );
  INV_X1 U820 ( .A(n482), .ZN(n817) );
  INV_X1 U821 ( .A(n814), .ZN(n818) );
  INV_X1 U822 ( .A(N7112), .ZN(n819) );
  INV_X1 U823 ( .A(n819), .ZN(n820) );
  INV_X1 U824 ( .A(n481), .ZN(n821) );
  INV_X1 U825 ( .A(n481), .ZN(n822) );
  INV_X1 U826 ( .A(n819), .ZN(n823) );
  INV_X1 U827 ( .A(N7204), .ZN(n824) );
  INV_X1 U828 ( .A(n824), .ZN(n825) );
  INV_X1 U829 ( .A(n480), .ZN(n826) );
  INV_X1 U830 ( .A(n480), .ZN(n827) );
  INV_X1 U831 ( .A(n824), .ZN(n828) );
  INV_X1 U832 ( .A(N7286), .ZN(n829) );
  INV_X1 U833 ( .A(n829), .ZN(n830) );
  INV_X1 U834 ( .A(n479), .ZN(n831) );
  INV_X1 U835 ( .A(n479), .ZN(n832) );
  INV_X1 U836 ( .A(n829), .ZN(n833) );
  INV_X1 U837 ( .A(N7375), .ZN(n834) );
  INV_X1 U838 ( .A(n834), .ZN(n835) );
  INV_X1 U839 ( .A(n478), .ZN(n836) );
  INV_X1 U840 ( .A(n478), .ZN(n837) );
  INV_X1 U841 ( .A(n834), .ZN(n838) );
  INV_X1 U842 ( .A(N7454), .ZN(n839) );
  INV_X1 U843 ( .A(n839), .ZN(n840) );
  INV_X1 U844 ( .A(n477), .ZN(n841) );
  INV_X1 U845 ( .A(n477), .ZN(n842) );
  INV_X1 U846 ( .A(n839), .ZN(n843) );
  INV_X1 U847 ( .A(N7543), .ZN(n844) );
  INV_X1 U848 ( .A(n844), .ZN(n845) );
  INV_X1 U849 ( .A(n476), .ZN(n846) );
  INV_X1 U850 ( .A(n476), .ZN(n847) );
  INV_X1 U851 ( .A(n844), .ZN(n848) );
  INV_X1 U852 ( .A(N7622), .ZN(n849) );
  INV_X1 U853 ( .A(n849), .ZN(n850) );
  INV_X1 U854 ( .A(n475), .ZN(n851) );
  INV_X1 U855 ( .A(n475), .ZN(n852) );
  INV_X1 U856 ( .A(n849), .ZN(n853) );
  INV_X1 U857 ( .A(N7711), .ZN(n854) );
  INV_X1 U858 ( .A(n854), .ZN(n855) );
  INV_X1 U859 ( .A(n474), .ZN(n856) );
  INV_X1 U860 ( .A(n474), .ZN(n857) );
  INV_X1 U861 ( .A(n854), .ZN(n858) );
  INV_X1 U862 ( .A(N7790), .ZN(n859) );
  INV_X1 U863 ( .A(n859), .ZN(n860) );
  INV_X1 U864 ( .A(n473), .ZN(n861) );
  INV_X1 U865 ( .A(n473), .ZN(n862) );
  INV_X1 U866 ( .A(n859), .ZN(n863) );
  INV_X1 U867 ( .A(N7879), .ZN(n864) );
  INV_X1 U868 ( .A(n864), .ZN(n865) );
  INV_X1 U869 ( .A(n472), .ZN(n866) );
  INV_X1 U870 ( .A(n472), .ZN(n867) );
  INV_X1 U871 ( .A(n864), .ZN(n868) );
  INV_X1 U872 ( .A(N7961), .ZN(n869) );
  INV_X1 U873 ( .A(n869), .ZN(n870) );
  INV_X1 U874 ( .A(n471), .ZN(n871) );
  INV_X1 U875 ( .A(n471), .ZN(n872) );
  INV_X1 U876 ( .A(n869), .ZN(n873) );
  INV_X1 U877 ( .A(cycle_num[0]), .ZN(n874) );
  INV_X1 U878 ( .A(n874), .ZN(n875) );
  INV_X1 U879 ( .A(n874), .ZN(n876) );
  INV_X1 U880 ( .A(n470), .ZN(n877) );
  INV_X1 U881 ( .A(n25664), .ZN(n878) );
  INV_X1 U882 ( .A(n470), .ZN(n879) );
  INV_X1 U883 ( .A(n25663), .ZN(n880) );
  INV_X1 U884 ( .A(n468), .ZN(n882) );
  INV_X1 U885 ( .A(n469), .ZN(n883) );
  INV_X1 U886 ( .A(n468), .ZN(n884) );
  INV_X1 U887 ( .A(n469), .ZN(n885) );
  BUF_X1 U888 ( .A(n277201), .Z(n886) );
  BUF_X1 U889 ( .A(n27721), .Z(n887) );
  BUF_X1 U890 ( .A(n27722), .Z(n888) );
  BUF_X1 U891 ( .A(n27723), .Z(n889) );
  BUF_X1 U892 ( .A(n27724), .Z(n890) );
  BUF_X1 U893 ( .A(n27725), .Z(n891) );
  BUF_X1 U894 ( .A(n27714), .Z(n892) );
  BUF_X1 U895 ( .A(n27715), .Z(n893) );
  BUF_X1 U896 ( .A(n27716), .Z(n894) );
  BUF_X1 U897 ( .A(n27717), .Z(n895) );
  BUF_X1 U898 ( .A(n27718), .Z(n896) );
  BUF_X1 U899 ( .A(n27719), .Z(n897) );
  BUF_X1 U900 ( .A(n27708), .Z(n898) );
  BUF_X1 U901 ( .A(n27709), .Z(n899) );
  BUF_X1 U902 ( .A(n277101), .Z(n900) );
  BUF_X1 U903 ( .A(n27711), .Z(n901) );
  BUF_X1 U904 ( .A(n27712), .Z(n902) );
  BUF_X1 U905 ( .A(n27713), .Z(n903) );
  BUF_X1 U906 ( .A(n907), .Z(n904) );
  INV_X1 U907 ( .A(matrix_mul_2D_7__5__14_), .ZN(n905) );
  INV_X1 U908 ( .A(n6341), .ZN(n906) );
  INV_X1 U909 ( .A(n906), .ZN(n907) );
  BUF_X1 U910 ( .A(n911), .Z(n908) );
  INV_X1 U911 ( .A(matrix_mul_2D_7__5__13_), .ZN(n909) );
  INV_X1 U912 ( .A(n6342), .ZN(n910) );
  INV_X1 U913 ( .A(n910), .ZN(n911) );
  BUF_X1 U914 ( .A(n915), .Z(n912) );
  INV_X1 U915 ( .A(matrix_mul_2D_7__5__12_), .ZN(n913) );
  INV_X1 U916 ( .A(n6343), .ZN(n914) );
  INV_X1 U917 ( .A(n914), .ZN(n915) );
  BUF_X1 U918 ( .A(n919), .Z(n916) );
  INV_X1 U919 ( .A(matrix_mul_2D_7__5__11_), .ZN(n917) );
  INV_X1 U920 ( .A(n6344), .ZN(n918) );
  INV_X1 U921 ( .A(n918), .ZN(n919) );
  BUF_X1 U922 ( .A(n923), .Z(n920) );
  INV_X1 U923 ( .A(matrix_mul_2D_7__5__10_), .ZN(n921) );
  INV_X1 U924 ( .A(n6345), .ZN(n922) );
  INV_X1 U925 ( .A(n922), .ZN(n923) );
  BUF_X1 U926 ( .A(n927), .Z(n924) );
  INV_X1 U927 ( .A(matrix_mul_2D_7__5__9_), .ZN(n925) );
  INV_X1 U928 ( .A(n6346), .ZN(n926) );
  INV_X1 U929 ( .A(n926), .ZN(n927) );
  BUF_X1 U930 ( .A(n931), .Z(n928) );
  INV_X1 U931 ( .A(matrix_mul_2D_7__5__8_), .ZN(n929) );
  INV_X1 U932 ( .A(n6347), .ZN(n930) );
  INV_X1 U933 ( .A(n930), .ZN(n931) );
  BUF_X1 U934 ( .A(n935), .Z(n932) );
  INV_X1 U935 ( .A(matrix_mul_2D_7__5__7_), .ZN(n933) );
  INV_X1 U936 ( .A(n6348), .ZN(n934) );
  INV_X1 U937 ( .A(n934), .ZN(n935) );
  BUF_X1 U938 ( .A(n939), .Z(n936) );
  INV_X1 U939 ( .A(matrix_mul_2D_7__5__6_), .ZN(n937) );
  INV_X1 U940 ( .A(n6349), .ZN(n938) );
  INV_X1 U941 ( .A(n938), .ZN(n939) );
  BUF_X1 U942 ( .A(n943), .Z(n940) );
  INV_X1 U943 ( .A(matrix_mul_2D_7__5__5_), .ZN(n941) );
  INV_X1 U944 ( .A(n63500), .ZN(n942) );
  INV_X1 U945 ( .A(n942), .ZN(n943) );
  BUF_X1 U946 ( .A(n947), .Z(n944) );
  INV_X1 U947 ( .A(matrix_mul_2D_7__5__4_), .ZN(n945) );
  INV_X1 U948 ( .A(n63510), .ZN(n946) );
  INV_X1 U949 ( .A(n946), .ZN(n947) );
  BUF_X1 U950 ( .A(n1922), .Z(n948) );
  INV_X1 U951 ( .A(matrix_mul_2D_7__5__3_), .ZN(n1920) );
  INV_X1 U952 ( .A(n63520), .ZN(n1921) );
  INV_X1 U953 ( .A(n1921), .ZN(n1922) );
  BUF_X1 U954 ( .A(n2205), .Z(n1923) );
  INV_X1 U955 ( .A(matrix_mul_2D_7__5__2_), .ZN(n1924) );
  INV_X1 U956 ( .A(n63530), .ZN(n1925) );
  INV_X1 U957 ( .A(n1925), .ZN(n2205) );
  BUF_X1 U958 ( .A(n2209), .Z(n2206) );
  INV_X1 U959 ( .A(matrix_mul_2D_7__5__1_), .ZN(n2207) );
  INV_X1 U960 ( .A(n63540), .ZN(n2208) );
  INV_X1 U961 ( .A(n2208), .ZN(n2209) );
  BUF_X1 U962 ( .A(n2289), .Z(n2210) );
  INV_X1 U963 ( .A(n28520), .ZN(n2286) );
  INV_X1 U964 ( .A(n2286), .ZN(n2287) );
  INV_X1 U965 ( .A(n63550), .ZN(n2288) );
  INV_X1 U966 ( .A(n2288), .ZN(n2289) );
  BUF_X1 U967 ( .A(n27702), .Z(n2290) );
  BUF_X1 U968 ( .A(n27703), .Z(n2291) );
  BUF_X1 U969 ( .A(n27704), .Z(n2427) );
  BUF_X1 U970 ( .A(n27705), .Z(n2428) );
  BUF_X1 U971 ( .A(n27706), .Z(n2429) );
  BUF_X1 U972 ( .A(n27707), .Z(n2430) );
  BUF_X1 U973 ( .A(n2554), .Z(n2431) );
  INV_X1 U974 ( .A(matrix_mul_2D_7__4__14_), .ZN(n2432) );
  INV_X1 U975 ( .A(n63260), .ZN(n2553) );
  INV_X1 U976 ( .A(n2553), .ZN(n2554) );
  BUF_X1 U977 ( .A(n2558), .Z(n2555) );
  INV_X1 U978 ( .A(matrix_mul_2D_7__4__13_), .ZN(n2556) );
  INV_X1 U979 ( .A(n63270), .ZN(n2557) );
  INV_X1 U980 ( .A(n2557), .ZN(n2558) );
  BUF_X1 U981 ( .A(n265200), .Z(n264900) );
  INV_X1 U982 ( .A(matrix_mul_2D_7__4__12_), .ZN(n265000) );
  INV_X1 U983 ( .A(n63280), .ZN(n265100) );
  INV_X1 U984 ( .A(n265100), .ZN(n265200) );
  BUF_X1 U985 ( .A(n268600), .Z(n265300) );
  INV_X1 U986 ( .A(matrix_mul_2D_7__4__11_), .ZN(n265400) );
  INV_X1 U987 ( .A(n63290), .ZN(n268500) );
  INV_X1 U988 ( .A(n268500), .ZN(n268600) );
  BUF_X1 U989 ( .A(n269000), .Z(n268700) );
  INV_X1 U990 ( .A(matrix_mul_2D_7__4__10_), .ZN(n268800) );
  INV_X1 U991 ( .A(n63300), .ZN(n268900) );
  INV_X1 U992 ( .A(n268900), .ZN(n269000) );
  BUF_X1 U993 ( .A(n278400), .Z(n278100) );
  INV_X1 U994 ( .A(matrix_mul_2D_7__4__9_), .ZN(n278200) );
  INV_X1 U995 ( .A(n63310), .ZN(n278300) );
  INV_X1 U996 ( .A(n278300), .ZN(n278400) );
  BUF_X1 U997 ( .A(n28180), .Z(n278500) );
  INV_X1 U998 ( .A(matrix_mul_2D_7__4__8_), .ZN(n278600) );
  INV_X1 U999 ( .A(n63320), .ZN(n28170) );
  INV_X1 U1000 ( .A(n28170), .ZN(n28180) );
  BUF_X1 U1001 ( .A(n28220), .Z(n28190) );
  INV_X1 U1002 ( .A(matrix_mul_2D_7__4__7_), .ZN(n28200) );
  INV_X1 U1003 ( .A(n6333), .ZN(n28210) );
  INV_X1 U1004 ( .A(n28210), .ZN(n28220) );
  BUF_X1 U1005 ( .A(n2886), .Z(n2883) );
  INV_X1 U1006 ( .A(matrix_mul_2D_7__4__6_), .ZN(n2884) );
  INV_X1 U1007 ( .A(n6334), .ZN(n2885) );
  INV_X1 U1008 ( .A(n2885), .ZN(n2886) );
  BUF_X1 U1009 ( .A(n2890), .Z(n2887) );
  INV_X1 U1010 ( .A(matrix_mul_2D_7__4__5_), .ZN(n2888) );
  INV_X1 U1011 ( .A(n6335), .ZN(n2889) );
  INV_X1 U1012 ( .A(n2889), .ZN(n2890) );
  BUF_X1 U1013 ( .A(n2894), .Z(n2891) );
  INV_X1 U1014 ( .A(matrix_mul_2D_7__4__4_), .ZN(n2892) );
  INV_X1 U1015 ( .A(n6336), .ZN(n2893) );
  INV_X1 U1016 ( .A(n2893), .ZN(n2894) );
  BUF_X1 U1017 ( .A(n2898), .Z(n2895) );
  INV_X1 U1018 ( .A(matrix_mul_2D_7__4__3_), .ZN(n2896) );
  INV_X1 U1019 ( .A(n6337), .ZN(n2897) );
  INV_X1 U1020 ( .A(n2897), .ZN(n2898) );
  BUF_X1 U1021 ( .A(n2902), .Z(n2899) );
  INV_X1 U1022 ( .A(matrix_mul_2D_7__4__2_), .ZN(n2900) );
  INV_X1 U1023 ( .A(n6338), .ZN(n2901) );
  INV_X1 U1024 ( .A(n2901), .ZN(n2902) );
  BUF_X1 U1025 ( .A(n2906), .Z(n29030) );
  INV_X1 U1026 ( .A(matrix_mul_2D_7__4__1_), .ZN(n2904) );
  INV_X1 U1027 ( .A(n6339), .ZN(n2905) );
  INV_X1 U1028 ( .A(n2905), .ZN(n2906) );
  BUF_X1 U1029 ( .A(n29110), .Z(n29070) );
  INV_X1 U1030 ( .A(n2837), .ZN(n29080) );
  INV_X1 U1031 ( .A(n29080), .ZN(n29090) );
  INV_X1 U1032 ( .A(n6340), .ZN(n29100) );
  INV_X1 U1033 ( .A(n29100), .ZN(n29110) );
  BUF_X1 U1034 ( .A(n27696), .Z(n29120) );
  BUF_X1 U1035 ( .A(n27697), .Z(n29130) );
  BUF_X1 U1036 ( .A(n27698), .Z(n29140) );
  BUF_X1 U1037 ( .A(n27699), .Z(n29150) );
  BUF_X1 U1038 ( .A(n277001), .Z(n29160) );
  BUF_X1 U1039 ( .A(n27701), .Z(n29170) );
  BUF_X1 U1040 ( .A(n29210), .Z(n29180) );
  INV_X1 U1041 ( .A(matrix_mul_2D_7__3__14_), .ZN(n29190) );
  INV_X1 U1042 ( .A(n6311), .ZN(n29200) );
  INV_X1 U1043 ( .A(n29200), .ZN(n29210) );
  BUF_X1 U1044 ( .A(n2925), .Z(n29220) );
  INV_X1 U1045 ( .A(matrix_mul_2D_7__3__13_), .ZN(n2923) );
  INV_X1 U1046 ( .A(n6312), .ZN(n2924) );
  INV_X1 U1047 ( .A(n2924), .ZN(n2925) );
  BUF_X1 U1048 ( .A(n2929), .Z(n2926) );
  INV_X1 U1049 ( .A(matrix_mul_2D_7__3__12_), .ZN(n2927) );
  INV_X1 U1050 ( .A(n6313), .ZN(n2928) );
  INV_X1 U1051 ( .A(n2928), .ZN(n2929) );
  BUF_X1 U1052 ( .A(n2933), .Z(n2930) );
  INV_X1 U1053 ( .A(matrix_mul_2D_7__3__11_), .ZN(n2931) );
  INV_X1 U1054 ( .A(n6314), .ZN(n2932) );
  INV_X1 U1055 ( .A(n2932), .ZN(n2933) );
  BUF_X1 U1056 ( .A(n2937), .Z(n2934) );
  INV_X1 U1057 ( .A(matrix_mul_2D_7__3__10_), .ZN(n2935) );
  INV_X1 U1058 ( .A(n6315), .ZN(n2936) );
  INV_X1 U1059 ( .A(n2936), .ZN(n2937) );
  BUF_X1 U1060 ( .A(n29410), .Z(n2938) );
  INV_X1 U1061 ( .A(matrix_mul_2D_7__3__9_), .ZN(n2939) );
  INV_X1 U1062 ( .A(n6316), .ZN(n29400) );
  INV_X1 U1063 ( .A(n29400), .ZN(n29410) );
  BUF_X1 U1064 ( .A(n29450), .Z(n29420) );
  INV_X1 U1065 ( .A(matrix_mul_2D_7__3__8_), .ZN(n29430) );
  INV_X1 U1066 ( .A(n63170), .ZN(n29440) );
  INV_X1 U1067 ( .A(n29440), .ZN(n29450) );
  BUF_X1 U1068 ( .A(n29490), .Z(n29460) );
  INV_X1 U1069 ( .A(matrix_mul_2D_7__3__7_), .ZN(n29470) );
  INV_X1 U1070 ( .A(n63180), .ZN(n29480) );
  INV_X1 U1071 ( .A(n29480), .ZN(n29490) );
  BUF_X1 U1072 ( .A(n29530), .Z(n29500) );
  INV_X1 U1073 ( .A(matrix_mul_2D_7__3__6_), .ZN(n29510) );
  INV_X1 U1074 ( .A(n63190), .ZN(n29520) );
  INV_X1 U1075 ( .A(n29520), .ZN(n29530) );
  BUF_X1 U1076 ( .A(n29570), .Z(n29540) );
  INV_X1 U1077 ( .A(matrix_mul_2D_7__3__5_), .ZN(n29550) );
  INV_X1 U1078 ( .A(n63200), .ZN(n29560) );
  INV_X1 U1079 ( .A(n29560), .ZN(n29570) );
  BUF_X1 U1080 ( .A(n2961), .Z(n29580) );
  INV_X1 U1081 ( .A(matrix_mul_2D_7__3__4_), .ZN(n29590) );
  INV_X1 U1082 ( .A(n63210), .ZN(n29600) );
  INV_X1 U1083 ( .A(n29600), .ZN(n2961) );
  BUF_X1 U1084 ( .A(n2965), .Z(n2962) );
  INV_X1 U1085 ( .A(matrix_mul_2D_7__3__3_), .ZN(n2963) );
  INV_X1 U1086 ( .A(n63220), .ZN(n2964) );
  INV_X1 U1087 ( .A(n2964), .ZN(n2965) );
  BUF_X1 U1088 ( .A(n2969), .Z(n2966) );
  INV_X1 U1089 ( .A(matrix_mul_2D_7__3__2_), .ZN(n2967) );
  INV_X1 U1090 ( .A(n63230), .ZN(n2968) );
  INV_X1 U1091 ( .A(n2968), .ZN(n2969) );
  BUF_X1 U1092 ( .A(n2973), .Z(n2970) );
  INV_X1 U1093 ( .A(matrix_mul_2D_7__3__1_), .ZN(n2971) );
  INV_X1 U1094 ( .A(n63240), .ZN(n2972) );
  INV_X1 U1095 ( .A(n2972), .ZN(n2973) );
  BUF_X1 U1096 ( .A(n2978), .Z(n2974) );
  INV_X1 U1097 ( .A(n28160), .ZN(n2975) );
  INV_X1 U1098 ( .A(n2975), .ZN(n2976) );
  INV_X1 U1099 ( .A(n63250), .ZN(n2977) );
  INV_X1 U1100 ( .A(n2977), .ZN(n2978) );
  BUF_X1 U1101 ( .A(n276901), .Z(n2979) );
  BUF_X1 U1102 ( .A(n27691), .Z(n2980) );
  BUF_X1 U1103 ( .A(n27692), .Z(n2981) );
  BUF_X1 U1104 ( .A(n27693), .Z(n2982) );
  BUF_X1 U1105 ( .A(n27694), .Z(n2983) );
  BUF_X1 U1106 ( .A(n27695), .Z(n2984) );
  BUF_X1 U1107 ( .A(n2988), .Z(n29850) );
  INV_X1 U1108 ( .A(matrix_mul_2D_7__2__14_), .ZN(n2986) );
  INV_X1 U1109 ( .A(n6296), .ZN(n2987) );
  INV_X1 U1110 ( .A(n2987), .ZN(n2988) );
  BUF_X1 U1111 ( .A(n29920), .Z(n29890) );
  INV_X1 U1112 ( .A(matrix_mul_2D_7__2__13_), .ZN(n29900) );
  INV_X1 U1113 ( .A(n6297), .ZN(n29910) );
  INV_X1 U1114 ( .A(n29910), .ZN(n29920) );
  BUF_X1 U1115 ( .A(n29960), .Z(n29930) );
  INV_X1 U1116 ( .A(matrix_mul_2D_7__2__12_), .ZN(n29940) );
  INV_X1 U1117 ( .A(n6298), .ZN(n29950) );
  INV_X1 U1118 ( .A(n29950), .ZN(n29960) );
  BUF_X1 U1119 ( .A(n30000), .Z(n29970) );
  INV_X1 U1120 ( .A(matrix_mul_2D_7__2__11_), .ZN(n29980) );
  INV_X1 U1121 ( .A(n6299), .ZN(n29990) );
  INV_X1 U1122 ( .A(n29990), .ZN(n30000) );
  BUF_X1 U1123 ( .A(n30040), .Z(n30010) );
  INV_X1 U1124 ( .A(matrix_mul_2D_7__2__10_), .ZN(n30020) );
  INV_X1 U1125 ( .A(n6300), .ZN(n30030) );
  INV_X1 U1126 ( .A(n30030), .ZN(n30040) );
  BUF_X1 U1127 ( .A(n3008), .Z(n3005) );
  INV_X1 U1128 ( .A(matrix_mul_2D_7__2__9_), .ZN(n3006) );
  INV_X1 U1129 ( .A(n6301), .ZN(n3007) );
  INV_X1 U1130 ( .A(n3007), .ZN(n3008) );
  BUF_X1 U1131 ( .A(n3012), .Z(n3009) );
  INV_X1 U1132 ( .A(matrix_mul_2D_7__2__8_), .ZN(n3010) );
  INV_X1 U1133 ( .A(n6302), .ZN(n3011) );
  INV_X1 U1134 ( .A(n3011), .ZN(n3012) );
  BUF_X1 U1135 ( .A(n3016), .Z(n3013) );
  INV_X1 U1136 ( .A(matrix_mul_2D_7__2__7_), .ZN(n3014) );
  INV_X1 U1137 ( .A(n6303), .ZN(n3015) );
  INV_X1 U1138 ( .A(n3015), .ZN(n3016) );
  BUF_X1 U1139 ( .A(n3020), .Z(n3017) );
  INV_X1 U1140 ( .A(matrix_mul_2D_7__2__6_), .ZN(n3018) );
  INV_X1 U1141 ( .A(n6304), .ZN(n3019) );
  INV_X1 U1142 ( .A(n3019), .ZN(n3020) );
  BUF_X1 U1143 ( .A(n30240), .Z(n3021) );
  INV_X1 U1144 ( .A(matrix_mul_2D_7__2__5_), .ZN(n30220) );
  INV_X1 U1145 ( .A(n6305), .ZN(n30230) );
  INV_X1 U1146 ( .A(n30230), .ZN(n30240) );
  BUF_X1 U1147 ( .A(n30280), .Z(n30250) );
  INV_X1 U1148 ( .A(matrix_mul_2D_7__2__4_), .ZN(n30260) );
  INV_X1 U1149 ( .A(n6306), .ZN(n30270) );
  INV_X1 U1150 ( .A(n30270), .ZN(n30280) );
  BUF_X1 U1151 ( .A(n30320), .Z(n30290) );
  INV_X1 U1152 ( .A(matrix_mul_2D_7__2__3_), .ZN(n30300) );
  INV_X1 U1153 ( .A(n6307), .ZN(n30310) );
  INV_X1 U1154 ( .A(n30310), .ZN(n30320) );
  BUF_X1 U1155 ( .A(n30360), .Z(n30330) );
  INV_X1 U1156 ( .A(matrix_mul_2D_7__2__2_), .ZN(n30340) );
  INV_X1 U1157 ( .A(n6308), .ZN(n30350) );
  INV_X1 U1158 ( .A(n30350), .ZN(n30360) );
  BUF_X1 U1159 ( .A(n30400), .Z(n30370) );
  INV_X1 U1160 ( .A(matrix_mul_2D_7__2__1_), .ZN(n30380) );
  INV_X1 U1161 ( .A(n6309), .ZN(n30390) );
  INV_X1 U1162 ( .A(n30390), .ZN(n30400) );
  BUF_X1 U1163 ( .A(n3045), .Z(n30410) );
  INV_X1 U1164 ( .A(n2801), .ZN(n30420) );
  INV_X1 U1165 ( .A(n30420), .ZN(n3043) );
  INV_X1 U1166 ( .A(n6310), .ZN(n3044) );
  INV_X1 U1167 ( .A(n3044), .ZN(n3045) );
  BUF_X1 U1168 ( .A(n27684), .Z(n3046) );
  BUF_X1 U1169 ( .A(n27685), .Z(n3047) );
  BUF_X1 U1170 ( .A(n27686), .Z(n3048) );
  BUF_X1 U1171 ( .A(n27687), .Z(n3049) );
  BUF_X1 U1172 ( .A(n27688), .Z(n3050) );
  BUF_X1 U1173 ( .A(n27689), .Z(n3051) );
  BUF_X1 U1174 ( .A(n3056), .Z(n3052) );
  INV_X1 U1175 ( .A(n276600), .ZN(n3053) );
  INV_X1 U1176 ( .A(n3053), .ZN(n3054) );
  INV_X1 U1177 ( .A(n62810), .ZN(n3055) );
  INV_X1 U1178 ( .A(n3055), .ZN(n3056) );
  BUF_X1 U1179 ( .A(n3061), .Z(n3057) );
  INV_X1 U1180 ( .A(n276700), .ZN(n3058) );
  INV_X1 U1181 ( .A(n3058), .ZN(n3059) );
  INV_X1 U1182 ( .A(n6282), .ZN(n3060) );
  INV_X1 U1183 ( .A(n3060), .ZN(n3061) );
  BUF_X1 U1184 ( .A(n3066), .Z(n3062) );
  INV_X1 U1185 ( .A(n276800), .ZN(n3063) );
  INV_X1 U1186 ( .A(n3063), .ZN(n3064) );
  INV_X1 U1187 ( .A(n6283), .ZN(n3065) );
  INV_X1 U1188 ( .A(n3065), .ZN(n3066) );
  BUF_X1 U1189 ( .A(n30960), .Z(n3067) );
  INV_X1 U1190 ( .A(n276900), .ZN(n3068) );
  INV_X1 U1191 ( .A(n3068), .ZN(n3069) );
  INV_X1 U1192 ( .A(n6284), .ZN(n3071) );
  INV_X1 U1193 ( .A(n3071), .ZN(n30960) );
  BUF_X1 U1194 ( .A(n3136), .Z(n3100) );
  INV_X1 U1195 ( .A(n277000), .ZN(n3101) );
  INV_X1 U1196 ( .A(n3101), .ZN(n3110) );
  INV_X1 U1197 ( .A(n6285), .ZN(n3111) );
  INV_X1 U1198 ( .A(n3111), .ZN(n3136) );
  BUF_X1 U1199 ( .A(n3235), .Z(n3153) );
  INV_X1 U1200 ( .A(n277100), .ZN(n32030) );
  INV_X1 U1201 ( .A(n32030), .ZN(n32100) );
  INV_X1 U1202 ( .A(n6286), .ZN(n3228) );
  INV_X1 U1203 ( .A(n3228), .ZN(n3235) );
  BUF_X1 U1204 ( .A(n3442), .Z(n32530) );
  INV_X1 U1205 ( .A(n277200), .ZN(n32610) );
  INV_X1 U1206 ( .A(n32610), .ZN(n33010) );
  INV_X1 U1207 ( .A(n6287), .ZN(n34350) );
  INV_X1 U1208 ( .A(n34350), .ZN(n3442) );
  BUF_X1 U1209 ( .A(n43530), .Z(n3617) );
  INV_X1 U1210 ( .A(n277300), .ZN(n36240) );
  INV_X1 U1211 ( .A(n36240), .ZN(n38460) );
  INV_X1 U1212 ( .A(n6288), .ZN(n4171) );
  INV_X1 U1213 ( .A(n4171), .ZN(n43530) );
  BUF_X1 U1214 ( .A(n47070), .Z(n43540) );
  INV_X1 U1215 ( .A(n277400), .ZN(n43940) );
  INV_X1 U1216 ( .A(n43940), .ZN(n4568) );
  INV_X1 U1217 ( .A(n6289), .ZN(n47030) );
  INV_X1 U1218 ( .A(n47030), .ZN(n47070) );
  BUF_X1 U1219 ( .A(n4887), .Z(n47080) );
  INV_X1 U1220 ( .A(n277500), .ZN(n4722) );
  INV_X1 U1221 ( .A(n4722), .ZN(n47870) );
  INV_X1 U1222 ( .A(n6290), .ZN(n48800) );
  INV_X1 U1223 ( .A(n48800), .ZN(n4887) );
  BUF_X1 U1224 ( .A(n5201), .Z(n4888) );
  INV_X1 U1225 ( .A(n277600), .ZN(n50790) );
  INV_X1 U1226 ( .A(n50790), .ZN(n5107) );
  INV_X1 U1227 ( .A(n6291), .ZN(n51350) );
  INV_X1 U1228 ( .A(n51350), .ZN(n5201) );
  BUF_X1 U1229 ( .A(n74110), .Z(n5296) );
  INV_X1 U1230 ( .A(n277700), .ZN(n5416) );
  INV_X1 U1231 ( .A(n5416), .ZN(n5417) );
  INV_X1 U1232 ( .A(n6292), .ZN(n74100) );
  INV_X1 U1233 ( .A(n74100), .ZN(n74110) );
  BUF_X1 U1234 ( .A(n7416), .Z(n74120) );
  INV_X1 U1235 ( .A(n277800), .ZN(n74130) );
  INV_X1 U1236 ( .A(n74130), .ZN(n7414) );
  INV_X1 U1237 ( .A(n6293), .ZN(n7415) );
  INV_X1 U1238 ( .A(n7415), .ZN(n7416) );
  BUF_X1 U1239 ( .A(n7421), .Z(n7417) );
  INV_X1 U1240 ( .A(n277900), .ZN(n7418) );
  INV_X1 U1241 ( .A(n7418), .ZN(n7419) );
  INV_X1 U1242 ( .A(n6294), .ZN(n7420) );
  INV_X1 U1243 ( .A(n7420), .ZN(n7421) );
  BUF_X1 U1244 ( .A(n7425), .Z(n7422) );
  INV_X1 U1245 ( .A(matrix_mul_2D_7__1__0_), .ZN(n7423) );
  INV_X1 U1246 ( .A(n6295), .ZN(n7424) );
  INV_X1 U1247 ( .A(n7424), .ZN(n7425) );
  BUF_X1 U1248 ( .A(n27678), .Z(n7426) );
  BUF_X1 U1249 ( .A(n27679), .Z(n7427) );
  BUF_X1 U1250 ( .A(n276801), .Z(n7428) );
  BUF_X1 U1251 ( .A(n27681), .Z(n7429) );
  BUF_X1 U1252 ( .A(n27682), .Z(n7430) );
  BUF_X1 U1253 ( .A(n27683), .Z(n7431) );
  BUF_X1 U1254 ( .A(n7436), .Z(n7432) );
  INV_X1 U1255 ( .A(n2751), .ZN(n7433) );
  INV_X1 U1256 ( .A(n7433), .ZN(n7434) );
  INV_X1 U1257 ( .A(n62660), .ZN(n7435) );
  INV_X1 U1258 ( .A(n7435), .ZN(n7436) );
  BUF_X1 U1259 ( .A(n74410), .Z(n7437) );
  INV_X1 U1260 ( .A(n2752), .ZN(n7438) );
  INV_X1 U1261 ( .A(n7438), .ZN(n74390) );
  INV_X1 U1262 ( .A(n62670), .ZN(n74400) );
  INV_X1 U1263 ( .A(n74400), .ZN(n74410) );
  BUF_X1 U1264 ( .A(n74460), .Z(n74420) );
  INV_X1 U1265 ( .A(n2753), .ZN(n74430) );
  INV_X1 U1266 ( .A(n74430), .ZN(n74440) );
  INV_X1 U1267 ( .A(n62680), .ZN(n74450) );
  INV_X1 U1268 ( .A(n74450), .ZN(n74460) );
  BUF_X1 U1269 ( .A(n74510), .Z(n74470) );
  INV_X1 U1270 ( .A(n2754), .ZN(n74480) );
  INV_X1 U1271 ( .A(n74480), .ZN(n74490) );
  INV_X1 U1272 ( .A(n62690), .ZN(n74500) );
  INV_X1 U1273 ( .A(n74500), .ZN(n74510) );
  BUF_X1 U1274 ( .A(n7456), .Z(n74520) );
  INV_X1 U1275 ( .A(n2755), .ZN(n74530) );
  INV_X1 U1276 ( .A(n74530), .ZN(n74540) );
  INV_X1 U1277 ( .A(n62700), .ZN(n7455) );
  INV_X1 U1278 ( .A(n7455), .ZN(n7456) );
  BUF_X1 U1279 ( .A(n7461), .Z(n7457) );
  INV_X1 U1280 ( .A(n2756), .ZN(n7458) );
  INV_X1 U1281 ( .A(n7458), .ZN(n7459) );
  INV_X1 U1282 ( .A(n62710), .ZN(n7460) );
  INV_X1 U1283 ( .A(n7460), .ZN(n7461) );
  BUF_X1 U1284 ( .A(n7466), .Z(n7462) );
  INV_X1 U1285 ( .A(n2757), .ZN(n7463) );
  INV_X1 U1286 ( .A(n7463), .ZN(n7464) );
  INV_X1 U1287 ( .A(n62720), .ZN(n7465) );
  INV_X1 U1288 ( .A(n7465), .ZN(n7466) );
  BUF_X1 U1289 ( .A(n7471), .Z(n7467) );
  INV_X1 U1290 ( .A(n2758), .ZN(n7468) );
  INV_X1 U1291 ( .A(n7468), .ZN(n7469) );
  INV_X1 U1292 ( .A(n62730), .ZN(n7470) );
  INV_X1 U1293 ( .A(n7470), .ZN(n7471) );
  BUF_X1 U1294 ( .A(n74760), .Z(n74720) );
  INV_X1 U1295 ( .A(n2759), .ZN(n74730) );
  INV_X1 U1296 ( .A(n74730), .ZN(n74740) );
  INV_X1 U1297 ( .A(n62740), .ZN(n74750) );
  INV_X1 U1298 ( .A(n74750), .ZN(n74760) );
  BUF_X1 U1299 ( .A(n74810), .Z(n74770) );
  INV_X1 U1300 ( .A(n2760), .ZN(n74780) );
  INV_X1 U1301 ( .A(n74780), .ZN(n74790) );
  INV_X1 U1302 ( .A(n62750), .ZN(n74800) );
  INV_X1 U1303 ( .A(n74800), .ZN(n74810) );
  BUF_X1 U1304 ( .A(n74860), .Z(n74820) );
  INV_X1 U1305 ( .A(n2761), .ZN(n74830) );
  INV_X1 U1306 ( .A(n74830), .ZN(n74840) );
  INV_X1 U1307 ( .A(n62760), .ZN(n74850) );
  INV_X1 U1308 ( .A(n74850), .ZN(n74860) );
  BUF_X1 U1309 ( .A(n74910), .Z(n74870) );
  INV_X1 U1310 ( .A(n2762), .ZN(n74880) );
  INV_X1 U1311 ( .A(n74880), .ZN(n74890) );
  INV_X1 U1312 ( .A(n62770), .ZN(n74900) );
  INV_X1 U1313 ( .A(n74900), .ZN(n74910) );
  BUF_X1 U1314 ( .A(n7496), .Z(n74920) );
  INV_X1 U1315 ( .A(n2763), .ZN(n7493) );
  INV_X1 U1316 ( .A(n7493), .ZN(n7494) );
  INV_X1 U1317 ( .A(n62780), .ZN(n7495) );
  INV_X1 U1318 ( .A(n7495), .ZN(n7496) );
  BUF_X1 U1319 ( .A(n7501), .Z(n7497) );
  INV_X1 U1320 ( .A(n2764), .ZN(n7498) );
  INV_X1 U1321 ( .A(n7498), .ZN(n7499) );
  INV_X1 U1322 ( .A(n62790), .ZN(n7500) );
  INV_X1 U1323 ( .A(n7500), .ZN(n7501) );
  BUF_X1 U1324 ( .A(n7505), .Z(n7502) );
  INV_X1 U1325 ( .A(matrix_mul_2D_7__0__0_), .ZN(n7503) );
  INV_X1 U1326 ( .A(n62800), .ZN(n7504) );
  INV_X1 U1327 ( .A(n7504), .ZN(n7505) );
  BUF_X1 U1328 ( .A(n27672), .Z(n7506) );
  BUF_X1 U1329 ( .A(n27673), .Z(n7507) );
  BUF_X1 U1330 ( .A(n27674), .Z(n7508) );
  BUF_X1 U1331 ( .A(n27675), .Z(n7509) );
  BUF_X1 U1332 ( .A(n27676), .Z(n7510) );
  BUF_X1 U1333 ( .A(n27677), .Z(n7511) );
  BUF_X1 U1334 ( .A(n7516), .Z(n7512) );
  INV_X1 U1335 ( .A(n273700), .ZN(n7513) );
  INV_X1 U1336 ( .A(n7513), .ZN(n7514) );
  INV_X1 U1337 ( .A(n6252), .ZN(n7515) );
  INV_X1 U1338 ( .A(n7515), .ZN(n7516) );
  BUF_X1 U1339 ( .A(n27666), .Z(n7517) );
  BUF_X1 U1340 ( .A(n27667), .Z(n7518) );
  BUF_X1 U1341 ( .A(n27668), .Z(n7519) );
  BUF_X1 U1342 ( .A(n27669), .Z(n7520) );
  BUF_X1 U1343 ( .A(n276701), .Z(n7521) );
  BUF_X1 U1344 ( .A(n27671), .Z(n7522) );
  BUF_X1 U1345 ( .A(n7526), .Z(n7523) );
  INV_X1 U1346 ( .A(matrix_mul_2D_6__6__14_), .ZN(n7524) );
  INV_X1 U1347 ( .A(n62360), .ZN(n7525) );
  INV_X1 U1348 ( .A(n7525), .ZN(n7526) );
  BUF_X1 U1349 ( .A(n75300), .Z(n7527) );
  INV_X1 U1350 ( .A(matrix_mul_2D_6__6__13_), .ZN(n75280) );
  INV_X1 U1351 ( .A(n62370), .ZN(n75290) );
  INV_X1 U1352 ( .A(n75290), .ZN(n75300) );
  BUF_X1 U1353 ( .A(n75340), .Z(n75310) );
  INV_X1 U1354 ( .A(matrix_mul_2D_6__6__12_), .ZN(n75320) );
  INV_X1 U1355 ( .A(n62380), .ZN(n75330) );
  INV_X1 U1356 ( .A(n75330), .ZN(n75340) );
  BUF_X1 U1357 ( .A(n75380), .Z(n75350) );
  INV_X1 U1358 ( .A(matrix_mul_2D_6__6__11_), .ZN(n75360) );
  INV_X1 U1359 ( .A(n62390), .ZN(n75370) );
  INV_X1 U1360 ( .A(n75370), .ZN(n75380) );
  BUF_X1 U1361 ( .A(n75420), .Z(n75390) );
  INV_X1 U1362 ( .A(matrix_mul_2D_6__6__10_), .ZN(n75400) );
  INV_X1 U1363 ( .A(n62400), .ZN(n75410) );
  INV_X1 U1364 ( .A(n75410), .ZN(n75420) );
  BUF_X1 U1365 ( .A(n7546), .Z(n75430) );
  INV_X1 U1366 ( .A(matrix_mul_2D_6__6__9_), .ZN(n7544) );
  INV_X1 U1367 ( .A(n62410), .ZN(n7545) );
  INV_X1 U1368 ( .A(n7545), .ZN(n7546) );
  BUF_X1 U1369 ( .A(n7550), .Z(n7547) );
  INV_X1 U1370 ( .A(matrix_mul_2D_6__6__8_), .ZN(n7548) );
  INV_X1 U1371 ( .A(n62420), .ZN(n7549) );
  INV_X1 U1372 ( .A(n7549), .ZN(n7550) );
  BUF_X1 U1373 ( .A(n7554), .Z(n7551) );
  INV_X1 U1374 ( .A(matrix_mul_2D_6__6__7_), .ZN(n7552) );
  INV_X1 U1375 ( .A(n62430), .ZN(n7553) );
  INV_X1 U1376 ( .A(n7553), .ZN(n7554) );
  BUF_X1 U1377 ( .A(n7558), .Z(n7555) );
  INV_X1 U1378 ( .A(matrix_mul_2D_6__6__6_), .ZN(n7556) );
  INV_X1 U1379 ( .A(n6244), .ZN(n7557) );
  INV_X1 U1380 ( .A(n7557), .ZN(n7558) );
  BUF_X1 U1381 ( .A(n75620), .Z(n7559) );
  INV_X1 U1382 ( .A(matrix_mul_2D_6__6__5_), .ZN(n7560) );
  INV_X1 U1383 ( .A(n6245), .ZN(n75610) );
  INV_X1 U1384 ( .A(n75610), .ZN(n75620) );
  BUF_X1 U1385 ( .A(n75660), .Z(n75630) );
  INV_X1 U1386 ( .A(matrix_mul_2D_6__6__4_), .ZN(n75640) );
  INV_X1 U1387 ( .A(n6246), .ZN(n75650) );
  INV_X1 U1388 ( .A(n75650), .ZN(n75660) );
  BUF_X1 U1389 ( .A(n75700), .Z(n75670) );
  INV_X1 U1390 ( .A(matrix_mul_2D_6__6__3_), .ZN(n75680) );
  INV_X1 U1391 ( .A(n6247), .ZN(n75690) );
  INV_X1 U1392 ( .A(n75690), .ZN(n75700) );
  BUF_X1 U1393 ( .A(n75740), .Z(n75710) );
  INV_X1 U1394 ( .A(matrix_mul_2D_6__6__2_), .ZN(n75720) );
  INV_X1 U1395 ( .A(n6248), .ZN(n75730) );
  INV_X1 U1396 ( .A(n75730), .ZN(n75740) );
  BUF_X1 U1397 ( .A(n75780), .Z(n75750) );
  INV_X1 U1398 ( .A(matrix_mul_2D_6__6__1_), .ZN(n75760) );
  INV_X1 U1399 ( .A(n6249), .ZN(n75770) );
  INV_X1 U1400 ( .A(n75770), .ZN(n75780) );
  BUF_X1 U1401 ( .A(n7583), .Z(n75790) );
  INV_X1 U1402 ( .A(n273500), .ZN(n75800) );
  INV_X1 U1403 ( .A(n75800), .ZN(n75810) );
  INV_X1 U1404 ( .A(n6250), .ZN(n7582) );
  INV_X1 U1405 ( .A(n7582), .ZN(n7583) );
  BUF_X1 U1406 ( .A(n276601), .Z(n7584) );
  BUF_X1 U1407 ( .A(n27661), .Z(n7585) );
  BUF_X1 U1408 ( .A(n27662), .Z(n7586) );
  BUF_X1 U1409 ( .A(n27663), .Z(n7587) );
  BUF_X1 U1410 ( .A(n27664), .Z(n7588) );
  BUF_X1 U1411 ( .A(n27665), .Z(n7589) );
  BUF_X1 U1412 ( .A(n7594), .Z(n7590) );
  INV_X1 U1413 ( .A(n2706), .ZN(n7591) );
  INV_X1 U1414 ( .A(n7591), .ZN(n7592) );
  INV_X1 U1415 ( .A(n6221), .ZN(n7593) );
  INV_X1 U1416 ( .A(n7593), .ZN(n7594) );
  BUF_X1 U1417 ( .A(n7599), .Z(n7595) );
  INV_X1 U1418 ( .A(n2707), .ZN(n7596) );
  INV_X1 U1419 ( .A(n7596), .ZN(n7597) );
  INV_X1 U1420 ( .A(n6222), .ZN(n7598) );
  INV_X1 U1421 ( .A(n7598), .ZN(n7599) );
  BUF_X1 U1422 ( .A(n7604), .Z(n7600) );
  INV_X1 U1423 ( .A(n2708), .ZN(n7601) );
  INV_X1 U1424 ( .A(n7601), .ZN(n7602) );
  INV_X1 U1425 ( .A(n6223), .ZN(n7603) );
  INV_X1 U1426 ( .A(n7603), .ZN(n7604) );
  BUF_X1 U1427 ( .A(n76090), .Z(n7605) );
  INV_X1 U1428 ( .A(n2709), .ZN(n7606) );
  INV_X1 U1429 ( .A(n7606), .ZN(n76070) );
  INV_X1 U1430 ( .A(n6224), .ZN(n76080) );
  INV_X1 U1431 ( .A(n76080), .ZN(n76090) );
  BUF_X1 U1432 ( .A(n76140), .Z(n76100) );
  INV_X1 U1433 ( .A(n2710), .ZN(n76110) );
  INV_X1 U1434 ( .A(n76110), .ZN(n76120) );
  INV_X1 U1435 ( .A(n6225), .ZN(n76130) );
  INV_X1 U1436 ( .A(n76130), .ZN(n76140) );
  BUF_X1 U1437 ( .A(n76190), .Z(n76150) );
  INV_X1 U1438 ( .A(n2711), .ZN(n76160) );
  INV_X1 U1439 ( .A(n76160), .ZN(n76170) );
  INV_X1 U1440 ( .A(n6226), .ZN(n76180) );
  INV_X1 U1441 ( .A(n76180), .ZN(n76190) );
  BUF_X1 U1442 ( .A(n7624), .Z(n76200) );
  INV_X1 U1443 ( .A(n2712), .ZN(n76210) );
  INV_X1 U1444 ( .A(n76210), .ZN(n76220) );
  INV_X1 U1445 ( .A(n6227), .ZN(n7623) );
  INV_X1 U1446 ( .A(n7623), .ZN(n7624) );
  BUF_X1 U1447 ( .A(n7629), .Z(n7625) );
  INV_X1 U1448 ( .A(n2713), .ZN(n7626) );
  INV_X1 U1449 ( .A(n7626), .ZN(n7627) );
  INV_X1 U1450 ( .A(n62280), .ZN(n7628) );
  INV_X1 U1451 ( .A(n7628), .ZN(n7629) );
  BUF_X1 U1452 ( .A(n7634), .Z(n7630) );
  INV_X1 U1453 ( .A(n2714), .ZN(n7631) );
  INV_X1 U1454 ( .A(n7631), .ZN(n7632) );
  INV_X1 U1455 ( .A(n62290), .ZN(n7633) );
  INV_X1 U1456 ( .A(n7633), .ZN(n7634) );
  BUF_X1 U1457 ( .A(n7639), .Z(n7635) );
  INV_X1 U1458 ( .A(n2715), .ZN(n7636) );
  INV_X1 U1459 ( .A(n7636), .ZN(n7637) );
  INV_X1 U1460 ( .A(n62300), .ZN(n7638) );
  INV_X1 U1461 ( .A(n7638), .ZN(n7639) );
  BUF_X1 U1462 ( .A(n76440), .Z(n76400) );
  INV_X1 U1463 ( .A(n2716), .ZN(n76410) );
  INV_X1 U1464 ( .A(n76410), .ZN(n76420) );
  INV_X1 U1465 ( .A(n62310), .ZN(n76430) );
  INV_X1 U1466 ( .A(n76430), .ZN(n76440) );
  BUF_X1 U1467 ( .A(n76490), .Z(n76450) );
  INV_X1 U1468 ( .A(n2717), .ZN(n76460) );
  INV_X1 U1469 ( .A(n76460), .ZN(n76470) );
  INV_X1 U1470 ( .A(n62320), .ZN(n76480) );
  INV_X1 U1471 ( .A(n76480), .ZN(n76490) );
  BUF_X1 U1472 ( .A(n76540), .Z(n76500) );
  INV_X1 U1473 ( .A(n2718), .ZN(n76510) );
  INV_X1 U1474 ( .A(n76510), .ZN(n76520) );
  INV_X1 U1475 ( .A(n62330), .ZN(n76530) );
  INV_X1 U1476 ( .A(n76530), .ZN(n76540) );
  BUF_X1 U1477 ( .A(n76590), .Z(n76550) );
  INV_X1 U1478 ( .A(n2719), .ZN(n76560) );
  INV_X1 U1479 ( .A(n76560), .ZN(n76570) );
  INV_X1 U1480 ( .A(n62340), .ZN(n76580) );
  INV_X1 U1481 ( .A(n76580), .ZN(n76590) );
  BUF_X1 U1482 ( .A(n7663), .Z(n76600) );
  INV_X1 U1483 ( .A(matrix_mul_2D_6__5__0_), .ZN(n7661) );
  INV_X1 U1484 ( .A(n62350), .ZN(n7662) );
  INV_X1 U1485 ( .A(n7662), .ZN(n7663) );
  BUF_X1 U1486 ( .A(n27654), .Z(n7664) );
  BUF_X1 U1487 ( .A(n27655), .Z(n7665) );
  BUF_X1 U1488 ( .A(n27656), .Z(n7666) );
  BUF_X1 U1489 ( .A(n27657), .Z(n7667) );
  BUF_X1 U1490 ( .A(n27658), .Z(n7668) );
  BUF_X1 U1491 ( .A(n27659), .Z(n7669) );
  BUF_X1 U1492 ( .A(n7673), .Z(n7670) );
  INV_X1 U1493 ( .A(matrix_mul_2D_6__4__14_), .ZN(n7671) );
  INV_X1 U1494 ( .A(n6206), .ZN(n7672) );
  INV_X1 U1495 ( .A(n7672), .ZN(n7673) );
  BUF_X1 U1496 ( .A(n7677), .Z(n7674) );
  INV_X1 U1497 ( .A(matrix_mul_2D_6__4__13_), .ZN(n7675) );
  INV_X1 U1498 ( .A(n6207), .ZN(n7676) );
  INV_X1 U1499 ( .A(n7676), .ZN(n7677) );
  BUF_X1 U1500 ( .A(n7681), .Z(n7678) );
  INV_X1 U1501 ( .A(matrix_mul_2D_6__4__12_), .ZN(n7679) );
  INV_X1 U1502 ( .A(n6208), .ZN(n7680) );
  INV_X1 U1503 ( .A(n7680), .ZN(n7681) );
  BUF_X1 U1504 ( .A(n7685), .Z(n7682) );
  INV_X1 U1505 ( .A(matrix_mul_2D_6__4__11_), .ZN(n7683) );
  INV_X1 U1506 ( .A(n6209), .ZN(n7684) );
  INV_X1 U1507 ( .A(n7684), .ZN(n7685) );
  BUF_X1 U1508 ( .A(n7689), .Z(n7686) );
  INV_X1 U1509 ( .A(matrix_mul_2D_6__4__10_), .ZN(n7687) );
  INV_X1 U1510 ( .A(n6210), .ZN(n7688) );
  INV_X1 U1511 ( .A(n7688), .ZN(n7689) );
  BUF_X1 U1512 ( .A(n7693), .Z(n7690) );
  INV_X1 U1513 ( .A(matrix_mul_2D_6__4__9_), .ZN(n7691) );
  INV_X1 U1514 ( .A(n6211), .ZN(n7692) );
  INV_X1 U1515 ( .A(n7692), .ZN(n7693) );
  BUF_X1 U1516 ( .A(n76970), .Z(n7694) );
  INV_X1 U1517 ( .A(matrix_mul_2D_6__4__8_), .ZN(n7695) );
  INV_X1 U1518 ( .A(n6212), .ZN(n76960) );
  INV_X1 U1519 ( .A(n76960), .ZN(n76970) );
  BUF_X1 U1520 ( .A(n77010), .Z(n76980) );
  INV_X1 U1521 ( .A(matrix_mul_2D_6__4__7_), .ZN(n76990) );
  INV_X1 U1522 ( .A(n6213), .ZN(n77000) );
  INV_X1 U1523 ( .A(n77000), .ZN(n77010) );
  BUF_X1 U1524 ( .A(n77050), .Z(n77020) );
  INV_X1 U1525 ( .A(matrix_mul_2D_6__4__6_), .ZN(n77030) );
  INV_X1 U1526 ( .A(n6214), .ZN(n77040) );
  INV_X1 U1527 ( .A(n77040), .ZN(n77050) );
  BUF_X1 U1528 ( .A(n77090), .Z(n77060) );
  INV_X1 U1529 ( .A(matrix_mul_2D_6__4__5_), .ZN(n77070) );
  INV_X1 U1530 ( .A(n6215), .ZN(n77080) );
  INV_X1 U1531 ( .A(n77080), .ZN(n77090) );
  BUF_X1 U1532 ( .A(n7713), .Z(n77100) );
  INV_X1 U1533 ( .A(matrix_mul_2D_6__4__4_), .ZN(n77110) );
  INV_X1 U1534 ( .A(n6216), .ZN(n7712) );
  INV_X1 U1535 ( .A(n7712), .ZN(n7713) );
  BUF_X1 U1536 ( .A(n7717), .Z(n7714) );
  INV_X1 U1537 ( .A(matrix_mul_2D_6__4__3_), .ZN(n7715) );
  INV_X1 U1538 ( .A(n6217), .ZN(n7716) );
  INV_X1 U1539 ( .A(n7716), .ZN(n7717) );
  BUF_X1 U1540 ( .A(n7721), .Z(n7718) );
  INV_X1 U1541 ( .A(matrix_mul_2D_6__4__2_), .ZN(n7719) );
  INV_X1 U1542 ( .A(n6218), .ZN(n7720) );
  INV_X1 U1543 ( .A(n7720), .ZN(n7721) );
  BUF_X1 U1544 ( .A(n7725), .Z(n7722) );
  INV_X1 U1545 ( .A(matrix_mul_2D_6__4__1_), .ZN(n7723) );
  INV_X1 U1546 ( .A(n6219), .ZN(n7724) );
  INV_X1 U1547 ( .A(n7724), .ZN(n7725) );
  BUF_X1 U1548 ( .A(n77300), .Z(n7726) );
  INV_X1 U1549 ( .A(n2705), .ZN(n7727) );
  INV_X1 U1550 ( .A(n7727), .ZN(n7728) );
  INV_X1 U1551 ( .A(n6220), .ZN(n77290) );
  INV_X1 U1552 ( .A(n77290), .ZN(n77300) );
  BUF_X1 U1553 ( .A(n27648), .Z(n77310) );
  BUF_X1 U1554 ( .A(n27649), .Z(n77320) );
  BUF_X1 U1555 ( .A(n27650), .Z(n77330) );
  BUF_X1 U1556 ( .A(n27651), .Z(n77340) );
  BUF_X1 U1557 ( .A(n27652), .Z(n77350) );
  BUF_X1 U1558 ( .A(n27653), .Z(n77360) );
  BUF_X1 U1559 ( .A(n77400), .Z(n77370) );
  INV_X1 U1560 ( .A(matrix_mul_2D_6__3__14_), .ZN(n77380) );
  INV_X1 U1561 ( .A(n61910), .ZN(n77390) );
  INV_X1 U1562 ( .A(n77390), .ZN(n77400) );
  BUF_X1 U1563 ( .A(n77440), .Z(n77410) );
  INV_X1 U1564 ( .A(matrix_mul_2D_6__3__13_), .ZN(n77420) );
  INV_X1 U1565 ( .A(n61920), .ZN(n77430) );
  INV_X1 U1566 ( .A(n77430), .ZN(n77440) );
  BUF_X1 U1567 ( .A(n77480), .Z(n77450) );
  INV_X1 U1568 ( .A(matrix_mul_2D_6__3__12_), .ZN(n77460) );
  INV_X1 U1569 ( .A(n61930), .ZN(n77470) );
  INV_X1 U1570 ( .A(n77470), .ZN(n77480) );
  BUF_X1 U1571 ( .A(n7752), .Z(n77490) );
  INV_X1 U1572 ( .A(matrix_mul_2D_6__3__11_), .ZN(n7750) );
  INV_X1 U1573 ( .A(n61940), .ZN(n7751) );
  INV_X1 U1574 ( .A(n7751), .ZN(n7752) );
  BUF_X1 U1575 ( .A(n7756), .Z(n7753) );
  INV_X1 U1576 ( .A(matrix_mul_2D_6__3__10_), .ZN(n7754) );
  INV_X1 U1577 ( .A(n61950), .ZN(n7755) );
  INV_X1 U1578 ( .A(n7755), .ZN(n7756) );
  BUF_X1 U1579 ( .A(n7760), .Z(n7757) );
  INV_X1 U1580 ( .A(matrix_mul_2D_6__3__9_), .ZN(n7758) );
  INV_X1 U1581 ( .A(n61960), .ZN(n7759) );
  INV_X1 U1582 ( .A(n7759), .ZN(n7760) );
  BUF_X1 U1583 ( .A(n7764), .Z(n7761) );
  INV_X1 U1584 ( .A(matrix_mul_2D_6__3__8_), .ZN(n7762) );
  INV_X1 U1585 ( .A(n61970), .ZN(n7763) );
  INV_X1 U1586 ( .A(n7763), .ZN(n7764) );
  BUF_X1 U1587 ( .A(n7768), .Z(n7765) );
  INV_X1 U1588 ( .A(matrix_mul_2D_6__3__7_), .ZN(n7766) );
  INV_X1 U1589 ( .A(n61980), .ZN(n7767) );
  INV_X1 U1590 ( .A(n7767), .ZN(n7768) );
  BUF_X1 U1591 ( .A(n7772), .Z(n7769) );
  INV_X1 U1592 ( .A(matrix_mul_2D_6__3__6_), .ZN(n7770) );
  INV_X1 U1593 ( .A(n61990), .ZN(n7771) );
  INV_X1 U1594 ( .A(n7771), .ZN(n7772) );
  BUF_X1 U1595 ( .A(n77760), .Z(n7773) );
  INV_X1 U1596 ( .A(matrix_mul_2D_6__3__5_), .ZN(n7774) );
  INV_X1 U1597 ( .A(n62000), .ZN(n77750) );
  INV_X1 U1598 ( .A(n77750), .ZN(n77760) );
  BUF_X1 U1599 ( .A(n77800), .Z(n77770) );
  INV_X1 U1600 ( .A(matrix_mul_2D_6__3__4_), .ZN(n77780) );
  INV_X1 U1601 ( .A(n62010), .ZN(n77790) );
  INV_X1 U1602 ( .A(n77790), .ZN(n77800) );
  BUF_X1 U1603 ( .A(n77840), .Z(n77810) );
  INV_X1 U1604 ( .A(matrix_mul_2D_6__3__3_), .ZN(n77820) );
  INV_X1 U1605 ( .A(n62020), .ZN(n77830) );
  INV_X1 U1606 ( .A(n77830), .ZN(n77840) );
  BUF_X1 U1607 ( .A(n77880), .Z(n77850) );
  INV_X1 U1608 ( .A(matrix_mul_2D_6__3__2_), .ZN(n77860) );
  INV_X1 U1609 ( .A(n6203), .ZN(n77870) );
  INV_X1 U1610 ( .A(n77870), .ZN(n77880) );
  BUF_X1 U1611 ( .A(n7792), .Z(n77890) );
  INV_X1 U1612 ( .A(matrix_mul_2D_6__3__1_), .ZN(n77900) );
  INV_X1 U1613 ( .A(n6204), .ZN(n7791) );
  INV_X1 U1614 ( .A(n7791), .ZN(n7792) );
  BUF_X1 U1615 ( .A(n7797), .Z(n7793) );
  INV_X1 U1616 ( .A(n268400), .ZN(n7794) );
  INV_X1 U1617 ( .A(n7794), .ZN(n7795) );
  INV_X1 U1618 ( .A(n6205), .ZN(n7796) );
  INV_X1 U1619 ( .A(n7796), .ZN(n7797) );
  BUF_X1 U1620 ( .A(n27642), .Z(n7798) );
  BUF_X1 U1621 ( .A(n27643), .Z(n7799) );
  BUF_X1 U1622 ( .A(n27644), .Z(n7800) );
  BUF_X1 U1623 ( .A(n27645), .Z(n7801) );
  BUF_X1 U1624 ( .A(n27646), .Z(n7802) );
  BUF_X1 U1625 ( .A(n27647), .Z(n7803) );
  BUF_X1 U1626 ( .A(n7807), .Z(n7804) );
  INV_X1 U1627 ( .A(matrix_mul_2D_6__2__14_), .ZN(n7805) );
  INV_X1 U1628 ( .A(n6176), .ZN(n7806) );
  INV_X1 U1629 ( .A(n7806), .ZN(n7807) );
  BUF_X1 U1630 ( .A(n78110), .Z(n78080) );
  INV_X1 U1631 ( .A(matrix_mul_2D_6__2__13_), .ZN(n78090) );
  INV_X1 U1632 ( .A(n6177), .ZN(n78100) );
  INV_X1 U1633 ( .A(n78100), .ZN(n78110) );
  BUF_X1 U1634 ( .A(n78150), .Z(n78120) );
  INV_X1 U1635 ( .A(matrix_mul_2D_6__2__12_), .ZN(n78130) );
  INV_X1 U1636 ( .A(n6178), .ZN(n78140) );
  INV_X1 U1637 ( .A(n78140), .ZN(n78150) );
  BUF_X1 U1638 ( .A(n78190), .Z(n78160) );
  INV_X1 U1639 ( .A(matrix_mul_2D_6__2__11_), .ZN(n78170) );
  INV_X1 U1640 ( .A(n6179), .ZN(n78180) );
  INV_X1 U1641 ( .A(n78180), .ZN(n78190) );
  BUF_X1 U1642 ( .A(n78230), .Z(n78200) );
  INV_X1 U1643 ( .A(matrix_mul_2D_6__2__10_), .ZN(n78210) );
  INV_X1 U1644 ( .A(n6180), .ZN(n78220) );
  INV_X1 U1645 ( .A(n78220), .ZN(n78230) );
  BUF_X1 U1646 ( .A(n78270), .Z(n78240) );
  INV_X1 U1647 ( .A(matrix_mul_2D_6__2__9_), .ZN(n78250) );
  INV_X1 U1648 ( .A(n6181), .ZN(n78260) );
  INV_X1 U1649 ( .A(n78260), .ZN(n78270) );
  BUF_X1 U1650 ( .A(n7831), .Z(n78280) );
  INV_X1 U1651 ( .A(matrix_mul_2D_6__2__8_), .ZN(n7829) );
  INV_X1 U1652 ( .A(n61820), .ZN(n7830) );
  INV_X1 U1653 ( .A(n7830), .ZN(n7831) );
  BUF_X1 U1654 ( .A(n7835), .Z(n7832) );
  INV_X1 U1655 ( .A(matrix_mul_2D_6__2__7_), .ZN(n7833) );
  INV_X1 U1656 ( .A(n61830), .ZN(n7834) );
  INV_X1 U1657 ( .A(n7834), .ZN(n7835) );
  BUF_X1 U1658 ( .A(n7839), .Z(n7836) );
  INV_X1 U1659 ( .A(matrix_mul_2D_6__2__6_), .ZN(n7837) );
  INV_X1 U1660 ( .A(n61840), .ZN(n7838) );
  INV_X1 U1661 ( .A(n7838), .ZN(n7839) );
  BUF_X1 U1662 ( .A(n7843), .Z(n7840) );
  INV_X1 U1663 ( .A(matrix_mul_2D_6__2__5_), .ZN(n7841) );
  INV_X1 U1664 ( .A(n61850), .ZN(n7842) );
  INV_X1 U1665 ( .A(n7842), .ZN(n7843) );
  BUF_X1 U1666 ( .A(n7847), .Z(n7844) );
  INV_X1 U1667 ( .A(matrix_mul_2D_6__2__4_), .ZN(n7845) );
  INV_X1 U1668 ( .A(n61860), .ZN(n7846) );
  INV_X1 U1669 ( .A(n7846), .ZN(n7847) );
  BUF_X1 U1670 ( .A(n7851), .Z(n7848) );
  INV_X1 U1671 ( .A(matrix_mul_2D_6__2__3_), .ZN(n7849) );
  INV_X1 U1672 ( .A(n61870), .ZN(n7850) );
  INV_X1 U1673 ( .A(n7850), .ZN(n7851) );
  BUF_X1 U1674 ( .A(n7855), .Z(n7852) );
  INV_X1 U1675 ( .A(matrix_mul_2D_6__2__2_), .ZN(n7853) );
  INV_X1 U1676 ( .A(n61880), .ZN(n7854) );
  INV_X1 U1677 ( .A(n7854), .ZN(n7855) );
  BUF_X1 U1678 ( .A(n7859), .Z(n7856) );
  INV_X1 U1679 ( .A(matrix_mul_2D_6__2__1_), .ZN(n7857) );
  INV_X1 U1680 ( .A(n61890), .ZN(n7858) );
  INV_X1 U1681 ( .A(n7858), .ZN(n7859) );
  BUF_X1 U1682 ( .A(n78640), .Z(n7860) );
  INV_X1 U1683 ( .A(n2669), .ZN(n7861) );
  INV_X1 U1684 ( .A(n7861), .ZN(n7862) );
  INV_X1 U1685 ( .A(n61900), .ZN(n7863) );
  INV_X1 U1686 ( .A(n7863), .ZN(n78640) );
  BUF_X1 U1687 ( .A(n27636), .Z(n78650) );
  BUF_X1 U1688 ( .A(n27637), .Z(n78660) );
  BUF_X1 U1689 ( .A(n27638), .Z(n78670) );
  BUF_X1 U1690 ( .A(n27639), .Z(n78680) );
  BUF_X1 U1691 ( .A(n27640), .Z(n78690) );
  BUF_X1 U1692 ( .A(n27641), .Z(n78700) );
  BUF_X1 U1693 ( .A(n78750), .Z(n78710) );
  INV_X1 U1694 ( .A(n2634), .ZN(n78720) );
  INV_X1 U1695 ( .A(n78720), .ZN(n78730) );
  INV_X1 U1696 ( .A(n61610), .ZN(n78740) );
  INV_X1 U1697 ( .A(n78740), .ZN(n78750) );
  BUF_X1 U1698 ( .A(n7880), .Z(n78760) );
  INV_X1 U1699 ( .A(n2635), .ZN(n78770) );
  INV_X1 U1700 ( .A(n78770), .ZN(n78780) );
  INV_X1 U1701 ( .A(n61620), .ZN(n78790) );
  INV_X1 U1702 ( .A(n78790), .ZN(n7880) );
  BUF_X1 U1703 ( .A(n7885), .Z(n7881) );
  INV_X1 U1704 ( .A(n2636), .ZN(n7882) );
  INV_X1 U1705 ( .A(n7882), .ZN(n7883) );
  INV_X1 U1706 ( .A(n61630), .ZN(n7884) );
  INV_X1 U1707 ( .A(n7884), .ZN(n7885) );
  BUF_X1 U1708 ( .A(n7890), .Z(n7886) );
  INV_X1 U1709 ( .A(n263700), .ZN(n7887) );
  INV_X1 U1710 ( .A(n7887), .ZN(n7888) );
  INV_X1 U1711 ( .A(n61640), .ZN(n7889) );
  INV_X1 U1712 ( .A(n7889), .ZN(n7890) );
  BUF_X1 U1713 ( .A(n7895), .Z(n7891) );
  INV_X1 U1714 ( .A(n2638), .ZN(n7892) );
  INV_X1 U1715 ( .A(n7892), .ZN(n7893) );
  INV_X1 U1716 ( .A(n6165), .ZN(n7894) );
  INV_X1 U1717 ( .A(n7894), .ZN(n7895) );
  BUF_X1 U1718 ( .A(n79000), .Z(n7896) );
  INV_X1 U1719 ( .A(n2639), .ZN(n78970) );
  INV_X1 U1720 ( .A(n78970), .ZN(n78980) );
  INV_X1 U1721 ( .A(n6166), .ZN(n78990) );
  INV_X1 U1722 ( .A(n78990), .ZN(n79000) );
  BUF_X1 U1723 ( .A(n79050), .Z(n79010) );
  INV_X1 U1724 ( .A(n2640), .ZN(n79020) );
  INV_X1 U1725 ( .A(n79020), .ZN(n79030) );
  INV_X1 U1726 ( .A(n6167), .ZN(n79040) );
  INV_X1 U1727 ( .A(n79040), .ZN(n79050) );
  BUF_X1 U1728 ( .A(n79100), .Z(n79060) );
  INV_X1 U1729 ( .A(n264100), .ZN(n79070) );
  INV_X1 U1730 ( .A(n79070), .ZN(n79080) );
  INV_X1 U1731 ( .A(n6168), .ZN(n79090) );
  INV_X1 U1732 ( .A(n79090), .ZN(n79100) );
  BUF_X1 U1733 ( .A(n79150), .Z(n79110) );
  INV_X1 U1734 ( .A(n264200), .ZN(n79120) );
  INV_X1 U1735 ( .A(n79120), .ZN(n79130) );
  INV_X1 U1736 ( .A(n6169), .ZN(n79140) );
  INV_X1 U1737 ( .A(n79140), .ZN(n79150) );
  BUF_X1 U1738 ( .A(n7920), .Z(n79160) );
  INV_X1 U1739 ( .A(n264300), .ZN(n79170) );
  INV_X1 U1740 ( .A(n79170), .ZN(n7918) );
  INV_X1 U1741 ( .A(n6170), .ZN(n7919) );
  INV_X1 U1742 ( .A(n7919), .ZN(n7920) );
  BUF_X1 U1743 ( .A(n7925), .Z(n7921) );
  INV_X1 U1744 ( .A(n264400), .ZN(n7922) );
  INV_X1 U1745 ( .A(n7922), .ZN(n7923) );
  INV_X1 U1746 ( .A(n6171), .ZN(n7924) );
  INV_X1 U1747 ( .A(n7924), .ZN(n7925) );
  BUF_X1 U1748 ( .A(n7930), .Z(n7926) );
  INV_X1 U1749 ( .A(n264500), .ZN(n7927) );
  INV_X1 U1750 ( .A(n7927), .ZN(n7928) );
  INV_X1 U1751 ( .A(n6172), .ZN(n7929) );
  INV_X1 U1752 ( .A(n7929), .ZN(n7930) );
  BUF_X1 U1753 ( .A(n7935), .Z(n7931) );
  INV_X1 U1754 ( .A(n264600), .ZN(n7932) );
  INV_X1 U1755 ( .A(n7932), .ZN(n7933) );
  INV_X1 U1756 ( .A(n6173), .ZN(n7934) );
  INV_X1 U1757 ( .A(n7934), .ZN(n7935) );
  BUF_X1 U1758 ( .A(n7940), .Z(n7936) );
  INV_X1 U1759 ( .A(n264700), .ZN(n7937) );
  INV_X1 U1760 ( .A(n7937), .ZN(n7938) );
  INV_X1 U1761 ( .A(n6174), .ZN(n7939) );
  INV_X1 U1762 ( .A(n7939), .ZN(n7940) );
  BUF_X1 U1763 ( .A(n7944), .Z(n7941) );
  INV_X1 U1764 ( .A(matrix_mul_2D_6__1__0_), .ZN(n79420) );
  INV_X1 U1765 ( .A(n6175), .ZN(n7943) );
  INV_X1 U1766 ( .A(n7943), .ZN(n7944) );
  BUF_X1 U1767 ( .A(n27630), .Z(n7945) );
  BUF_X1 U1768 ( .A(n27631), .Z(n79460) );
  BUF_X1 U1769 ( .A(n27632), .Z(n79470) );
  BUF_X1 U1770 ( .A(n27633), .Z(n79480) );
  BUF_X1 U1771 ( .A(n27634), .Z(n79490) );
  BUF_X1 U1772 ( .A(n27635), .Z(n79500) );
  BUF_X1 U1773 ( .A(n79550), .Z(n79510) );
  INV_X1 U1774 ( .A(n2619), .ZN(n79520) );
  INV_X1 U1775 ( .A(n79520), .ZN(n79530) );
  INV_X1 U1776 ( .A(n6146), .ZN(n79540) );
  INV_X1 U1777 ( .A(n79540), .ZN(n79550) );
  BUF_X1 U1778 ( .A(n79600), .Z(n79560) );
  INV_X1 U1779 ( .A(n2620), .ZN(n79570) );
  INV_X1 U1780 ( .A(n79570), .ZN(n79580) );
  INV_X1 U1781 ( .A(n6147), .ZN(n79590) );
  INV_X1 U1782 ( .A(n79590), .ZN(n79600) );
  BUF_X1 U1783 ( .A(n7965), .Z(n79610) );
  INV_X1 U1784 ( .A(n2621), .ZN(n7962) );
  INV_X1 U1785 ( .A(n7962), .ZN(n7963) );
  INV_X1 U1786 ( .A(n6148), .ZN(n7964) );
  INV_X1 U1787 ( .A(n7964), .ZN(n7965) );
  BUF_X1 U1788 ( .A(n7970), .Z(n7966) );
  INV_X1 U1789 ( .A(n2622), .ZN(n7967) );
  INV_X1 U1790 ( .A(n7967), .ZN(n7968) );
  INV_X1 U1791 ( .A(n61490), .ZN(n7969) );
  INV_X1 U1792 ( .A(n7969), .ZN(n7970) );
  BUF_X1 U1793 ( .A(n7975), .Z(n7971) );
  INV_X1 U1794 ( .A(n2623), .ZN(n7972) );
  INV_X1 U1795 ( .A(n7972), .ZN(n7973) );
  INV_X1 U1796 ( .A(n61500), .ZN(n7974) );
  INV_X1 U1797 ( .A(n7974), .ZN(n7975) );
  BUF_X1 U1798 ( .A(n79800), .Z(n7976) );
  INV_X1 U1799 ( .A(n2624), .ZN(n7977) );
  INV_X1 U1800 ( .A(n7977), .ZN(n7978) );
  INV_X1 U1801 ( .A(n61510), .ZN(n79790) );
  INV_X1 U1802 ( .A(n79790), .ZN(n79800) );
  BUF_X1 U1803 ( .A(n79850), .Z(n79810) );
  INV_X1 U1804 ( .A(n2625), .ZN(n79820) );
  INV_X1 U1805 ( .A(n79820), .ZN(n79830) );
  INV_X1 U1806 ( .A(n61520), .ZN(n79840) );
  INV_X1 U1807 ( .A(n79840), .ZN(n79850) );
  BUF_X1 U1808 ( .A(n79900), .Z(n79860) );
  INV_X1 U1809 ( .A(n2626), .ZN(n79870) );
  INV_X1 U1810 ( .A(n79870), .ZN(n79880) );
  INV_X1 U1811 ( .A(n61530), .ZN(n79890) );
  INV_X1 U1812 ( .A(n79890), .ZN(n79900) );
  BUF_X1 U1813 ( .A(n79950), .Z(n79910) );
  INV_X1 U1814 ( .A(n2627), .ZN(n79920) );
  INV_X1 U1815 ( .A(n79920), .ZN(n79930) );
  INV_X1 U1816 ( .A(n61540), .ZN(n79940) );
  INV_X1 U1817 ( .A(n79940), .ZN(n79950) );
  BUF_X1 U1818 ( .A(n8000), .Z(n79960) );
  INV_X1 U1819 ( .A(n2628), .ZN(n79970) );
  INV_X1 U1820 ( .A(n79970), .ZN(n79980) );
  INV_X1 U1821 ( .A(n61550), .ZN(n79990) );
  INV_X1 U1822 ( .A(n79990), .ZN(n8000) );
  BUF_X1 U1823 ( .A(n8005), .Z(n8001) );
  INV_X1 U1824 ( .A(n2629), .ZN(n8002) );
  INV_X1 U1825 ( .A(n8002), .ZN(n8003) );
  INV_X1 U1826 ( .A(n61560), .ZN(n8004) );
  INV_X1 U1827 ( .A(n8004), .ZN(n8005) );
  BUF_X1 U1828 ( .A(n8010), .Z(n8006) );
  INV_X1 U1829 ( .A(n2630), .ZN(n8007) );
  INV_X1 U1830 ( .A(n8007), .ZN(n8008) );
  INV_X1 U1831 ( .A(n61570), .ZN(n8009) );
  INV_X1 U1832 ( .A(n8009), .ZN(n8010) );
  BUF_X1 U1833 ( .A(n8015), .Z(n8011) );
  INV_X1 U1834 ( .A(n2631), .ZN(n8012) );
  INV_X1 U1835 ( .A(n8012), .ZN(n8013) );
  INV_X1 U1836 ( .A(n61580), .ZN(n8014) );
  INV_X1 U1837 ( .A(n8014), .ZN(n8015) );
  BUF_X1 U1838 ( .A(n8020), .Z(n8016) );
  INV_X1 U1839 ( .A(n2632), .ZN(n8017) );
  INV_X1 U1840 ( .A(n8017), .ZN(n8018) );
  INV_X1 U1841 ( .A(n61590), .ZN(n8019) );
  INV_X1 U1842 ( .A(n8019), .ZN(n8020) );
  BUF_X1 U1843 ( .A(n8024), .Z(n8021) );
  INV_X1 U1844 ( .A(matrix_mul_2D_6__0__0_), .ZN(n8022) );
  INV_X1 U1845 ( .A(n61600), .ZN(n8023) );
  INV_X1 U1846 ( .A(n8023), .ZN(n8024) );
  BUF_X1 U1847 ( .A(n27624), .Z(n8025) );
  BUF_X1 U1848 ( .A(n27625), .Z(n8026) );
  BUF_X1 U1849 ( .A(n27626), .Z(n8027) );
  BUF_X1 U1850 ( .A(n27627), .Z(n8028) );
  BUF_X1 U1851 ( .A(n27628), .Z(n8029) );
  BUF_X1 U1852 ( .A(n27629), .Z(n8030) );
  BUF_X1 U1853 ( .A(n8035), .Z(n8031) );
  INV_X1 U1854 ( .A(n260400), .ZN(n8032) );
  INV_X1 U1855 ( .A(n8032), .ZN(n8033) );
  INV_X1 U1856 ( .A(n6131), .ZN(n8034) );
  INV_X1 U1857 ( .A(n8034), .ZN(n8035) );
  BUF_X1 U1858 ( .A(n8040), .Z(n8036) );
  INV_X1 U1859 ( .A(n260500), .ZN(n8037) );
  INV_X1 U1860 ( .A(n8037), .ZN(n8038) );
  INV_X1 U1861 ( .A(n6132), .ZN(n8039) );
  INV_X1 U1862 ( .A(n8039), .ZN(n8040) );
  BUF_X1 U1863 ( .A(n8045), .Z(n8041) );
  INV_X1 U1864 ( .A(n260600), .ZN(n8042) );
  INV_X1 U1865 ( .A(n8042), .ZN(n8043) );
  INV_X1 U1866 ( .A(n6133), .ZN(n8044) );
  INV_X1 U1867 ( .A(n8044), .ZN(n8045) );
  BUF_X1 U1868 ( .A(n8050), .Z(n8046) );
  INV_X1 U1869 ( .A(n260700), .ZN(n8047) );
  INV_X1 U1870 ( .A(n8047), .ZN(n8048) );
  INV_X1 U1871 ( .A(n6134), .ZN(n8049) );
  INV_X1 U1872 ( .A(n8049), .ZN(n8050) );
  BUF_X1 U1873 ( .A(n8055), .Z(n8051) );
  INV_X1 U1874 ( .A(n260800), .ZN(n8052) );
  INV_X1 U1875 ( .A(n8052), .ZN(n8053) );
  INV_X1 U1876 ( .A(n6135), .ZN(n8054) );
  INV_X1 U1877 ( .A(n8054), .ZN(n8055) );
  BUF_X1 U1878 ( .A(n8060), .Z(n8056) );
  INV_X1 U1879 ( .A(n260900), .ZN(n8057) );
  INV_X1 U1880 ( .A(n8057), .ZN(n8058) );
  INV_X1 U1881 ( .A(n6136), .ZN(n8059) );
  INV_X1 U1882 ( .A(n8059), .ZN(n8060) );
  BUF_X1 U1883 ( .A(n8065), .Z(n8061) );
  INV_X1 U1884 ( .A(n261000), .ZN(n8062) );
  INV_X1 U1885 ( .A(n8062), .ZN(n8063) );
  INV_X1 U1886 ( .A(n6137), .ZN(n8064) );
  INV_X1 U1887 ( .A(n8064), .ZN(n8065) );
  BUF_X1 U1888 ( .A(n8070), .Z(n8066) );
  INV_X1 U1889 ( .A(n261100), .ZN(n8067) );
  INV_X1 U1890 ( .A(n8067), .ZN(n8068) );
  INV_X1 U1891 ( .A(n6138), .ZN(n8069) );
  INV_X1 U1892 ( .A(n8069), .ZN(n8070) );
  BUF_X1 U1893 ( .A(n8075), .Z(n8071) );
  INV_X1 U1894 ( .A(n261200), .ZN(n8072) );
  INV_X1 U1895 ( .A(n8072), .ZN(n8073) );
  INV_X1 U1896 ( .A(n6139), .ZN(n8074) );
  INV_X1 U1897 ( .A(n8074), .ZN(n8075) );
  BUF_X1 U1898 ( .A(n8080), .Z(n8076) );
  INV_X1 U1899 ( .A(n2613), .ZN(n8077) );
  INV_X1 U1900 ( .A(n8077), .ZN(n8078) );
  INV_X1 U1901 ( .A(n6140), .ZN(n8079) );
  INV_X1 U1902 ( .A(n8079), .ZN(n8080) );
  BUF_X1 U1903 ( .A(n8085), .Z(n8081) );
  INV_X1 U1904 ( .A(n2614), .ZN(n8082) );
  INV_X1 U1905 ( .A(n8082), .ZN(n8083) );
  INV_X1 U1906 ( .A(n6141), .ZN(n8084) );
  INV_X1 U1907 ( .A(n8084), .ZN(n8085) );
  BUF_X1 U1908 ( .A(n8090), .Z(n8086) );
  INV_X1 U1909 ( .A(n2615), .ZN(n8087) );
  INV_X1 U1910 ( .A(n8087), .ZN(n8088) );
  INV_X1 U1911 ( .A(n6142), .ZN(n8089) );
  INV_X1 U1912 ( .A(n8089), .ZN(n8090) );
  BUF_X1 U1913 ( .A(n8095), .Z(n8091) );
  INV_X1 U1914 ( .A(n2616), .ZN(n8092) );
  INV_X1 U1915 ( .A(n8092), .ZN(n8093) );
  INV_X1 U1916 ( .A(n6143), .ZN(n8094) );
  INV_X1 U1917 ( .A(n8094), .ZN(n8095) );
  BUF_X1 U1918 ( .A(n8100), .Z(n8096) );
  INV_X1 U1919 ( .A(n2617), .ZN(n8097) );
  INV_X1 U1920 ( .A(n8097), .ZN(n8098) );
  INV_X1 U1921 ( .A(n6144), .ZN(n8099) );
  INV_X1 U1922 ( .A(n8099), .ZN(n8100) );
  BUF_X1 U1923 ( .A(n8104), .Z(n8101) );
  INV_X1 U1924 ( .A(matrix_mul_2D_5__7__0_), .ZN(n8102) );
  INV_X1 U1925 ( .A(n6145), .ZN(n8103) );
  INV_X1 U1926 ( .A(n8103), .ZN(n8104) );
  BUF_X1 U1927 ( .A(n27618), .Z(n8105) );
  BUF_X1 U1928 ( .A(n27619), .Z(n8106) );
  BUF_X1 U1929 ( .A(n27620), .Z(n8107) );
  BUF_X1 U1930 ( .A(n27621), .Z(n8108) );
  BUF_X1 U1931 ( .A(n27622), .Z(n8109) );
  BUF_X1 U1932 ( .A(n27623), .Z(n8110) );
  BUF_X1 U1933 ( .A(n8115), .Z(n8111) );
  INV_X1 U1934 ( .A(n2589), .ZN(n8112) );
  INV_X1 U1935 ( .A(n8112), .ZN(n8113) );
  INV_X1 U1936 ( .A(n6116), .ZN(n8114) );
  INV_X1 U1937 ( .A(n8114), .ZN(n8115) );
  BUF_X1 U1938 ( .A(n8120), .Z(n8116) );
  INV_X1 U1939 ( .A(n2590), .ZN(n8117) );
  INV_X1 U1940 ( .A(n8117), .ZN(n8118) );
  INV_X1 U1941 ( .A(n6117), .ZN(n8119) );
  INV_X1 U1942 ( .A(n8119), .ZN(n8120) );
  BUF_X1 U1943 ( .A(n8125), .Z(n8121) );
  INV_X1 U1944 ( .A(n2591), .ZN(n8122) );
  INV_X1 U1945 ( .A(n8122), .ZN(n8123) );
  INV_X1 U1946 ( .A(n6118), .ZN(n8124) );
  INV_X1 U1947 ( .A(n8124), .ZN(n8125) );
  BUF_X1 U1948 ( .A(n8130), .Z(n8126) );
  INV_X1 U1949 ( .A(n259200), .ZN(n8127) );
  INV_X1 U1950 ( .A(n8127), .ZN(n8128) );
  INV_X1 U1951 ( .A(n6119), .ZN(n8129) );
  INV_X1 U1952 ( .A(n8129), .ZN(n8130) );
  BUF_X1 U1953 ( .A(n8135), .Z(n8131) );
  INV_X1 U1954 ( .A(n259300), .ZN(n8132) );
  INV_X1 U1955 ( .A(n8132), .ZN(n8133) );
  INV_X1 U1956 ( .A(n6120), .ZN(n8134) );
  INV_X1 U1957 ( .A(n8134), .ZN(n8135) );
  BUF_X1 U1958 ( .A(n8140), .Z(n8136) );
  INV_X1 U1959 ( .A(n259400), .ZN(n8137) );
  INV_X1 U1960 ( .A(n8137), .ZN(n8138) );
  INV_X1 U1961 ( .A(n6121), .ZN(n8139) );
  INV_X1 U1962 ( .A(n8139), .ZN(n8140) );
  BUF_X1 U1963 ( .A(n8145), .Z(n8141) );
  INV_X1 U1964 ( .A(n259500), .ZN(n8142) );
  INV_X1 U1965 ( .A(n8142), .ZN(n8143) );
  INV_X1 U1966 ( .A(n6122), .ZN(n8144) );
  INV_X1 U1967 ( .A(n8144), .ZN(n8145) );
  BUF_X1 U1968 ( .A(n8150), .Z(n8146) );
  INV_X1 U1969 ( .A(n259600), .ZN(n8147) );
  INV_X1 U1970 ( .A(n8147), .ZN(n8148) );
  INV_X1 U1971 ( .A(n6123), .ZN(n8149) );
  INV_X1 U1972 ( .A(n8149), .ZN(n8150) );
  BUF_X1 U1973 ( .A(n8155), .Z(n8151) );
  INV_X1 U1974 ( .A(n259700), .ZN(n8152) );
  INV_X1 U1975 ( .A(n8152), .ZN(n8153) );
  INV_X1 U1976 ( .A(n6124), .ZN(n8154) );
  INV_X1 U1977 ( .A(n8154), .ZN(n8155) );
  BUF_X1 U1978 ( .A(n8160), .Z(n8156) );
  INV_X1 U1979 ( .A(n259800), .ZN(n8157) );
  INV_X1 U1980 ( .A(n8157), .ZN(n8158) );
  INV_X1 U1981 ( .A(n6125), .ZN(n8159) );
  INV_X1 U1982 ( .A(n8159), .ZN(n8160) );
  BUF_X1 U1983 ( .A(n8165), .Z(n8161) );
  INV_X1 U1984 ( .A(n259900), .ZN(n8162) );
  INV_X1 U1985 ( .A(n8162), .ZN(n8163) );
  INV_X1 U1986 ( .A(n6126), .ZN(n8164) );
  INV_X1 U1987 ( .A(n8164), .ZN(n8165) );
  BUF_X1 U1988 ( .A(n8170), .Z(n8166) );
  INV_X1 U1989 ( .A(n260000), .ZN(n8167) );
  INV_X1 U1990 ( .A(n8167), .ZN(n8168) );
  INV_X1 U1991 ( .A(n6127), .ZN(n8169) );
  INV_X1 U1992 ( .A(n8169), .ZN(n8170) );
  BUF_X1 U1993 ( .A(n8175), .Z(n8171) );
  INV_X1 U1994 ( .A(n260100), .ZN(n8172) );
  INV_X1 U1995 ( .A(n8172), .ZN(n8173) );
  INV_X1 U1996 ( .A(n6128), .ZN(n8174) );
  INV_X1 U1997 ( .A(n8174), .ZN(n8175) );
  BUF_X1 U1998 ( .A(n8180), .Z(n8176) );
  INV_X1 U1999 ( .A(n260200), .ZN(n8177) );
  INV_X1 U2000 ( .A(n8177), .ZN(n8178) );
  INV_X1 U2001 ( .A(n6129), .ZN(n8179) );
  INV_X1 U2002 ( .A(n8179), .ZN(n8180) );
  BUF_X1 U2003 ( .A(n8184), .Z(n8181) );
  INV_X1 U2004 ( .A(matrix_mul_2D_5__6__0_), .ZN(n8182) );
  INV_X1 U2005 ( .A(n6130), .ZN(n8183) );
  INV_X1 U2006 ( .A(n8183), .ZN(n8184) );
  BUF_X1 U2007 ( .A(n27612), .Z(n8185) );
  BUF_X1 U2008 ( .A(n27613), .Z(n8186) );
  BUF_X1 U2009 ( .A(n27614), .Z(n8187) );
  BUF_X1 U2010 ( .A(n27615), .Z(n8188) );
  BUF_X1 U2011 ( .A(n27616), .Z(n8189) );
  BUF_X1 U2012 ( .A(n27617), .Z(n8190) );
  BUF_X1 U2013 ( .A(n8194), .Z(n8191) );
  INV_X1 U2014 ( .A(matrix_mul_2D_5__5__14_), .ZN(n8192) );
  INV_X1 U2015 ( .A(n61010), .ZN(n8193) );
  INV_X1 U2016 ( .A(n8193), .ZN(n8194) );
  BUF_X1 U2017 ( .A(n8198), .Z(n8195) );
  INV_X1 U2018 ( .A(matrix_mul_2D_5__5__13_), .ZN(n8196) );
  INV_X1 U2019 ( .A(n61020), .ZN(n8197) );
  INV_X1 U2020 ( .A(n8197), .ZN(n8198) );
  BUF_X1 U2021 ( .A(n8202), .Z(n8199) );
  INV_X1 U2022 ( .A(matrix_mul_2D_5__5__12_), .ZN(n8200) );
  INV_X1 U2023 ( .A(n61030), .ZN(n8201) );
  INV_X1 U2024 ( .A(n8201), .ZN(n8202) );
  BUF_X1 U2025 ( .A(n8206), .Z(n8203) );
  INV_X1 U2026 ( .A(matrix_mul_2D_5__5__11_), .ZN(n8204) );
  INV_X1 U2027 ( .A(n61040), .ZN(n8205) );
  INV_X1 U2028 ( .A(n8205), .ZN(n8206) );
  BUF_X1 U2029 ( .A(n8210), .Z(n8207) );
  INV_X1 U2030 ( .A(matrix_mul_2D_5__5__10_), .ZN(n8208) );
  INV_X1 U2031 ( .A(n61050), .ZN(n8209) );
  INV_X1 U2032 ( .A(n8209), .ZN(n8210) );
  BUF_X1 U2033 ( .A(n8214), .Z(n8211) );
  INV_X1 U2034 ( .A(matrix_mul_2D_5__5__9_), .ZN(n8212) );
  INV_X1 U2035 ( .A(n61060), .ZN(n8213) );
  INV_X1 U2036 ( .A(n8213), .ZN(n8214) );
  BUF_X1 U2037 ( .A(n8218), .Z(n8215) );
  INV_X1 U2038 ( .A(matrix_mul_2D_5__5__8_), .ZN(n8216) );
  INV_X1 U2039 ( .A(n61070), .ZN(n8217) );
  INV_X1 U2040 ( .A(n8217), .ZN(n8218) );
  BUF_X1 U2041 ( .A(n8222), .Z(n8219) );
  INV_X1 U2042 ( .A(matrix_mul_2D_5__5__7_), .ZN(n8220) );
  INV_X1 U2043 ( .A(n61080), .ZN(n8221) );
  INV_X1 U2044 ( .A(n8221), .ZN(n8222) );
  BUF_X1 U2045 ( .A(n8226), .Z(n8223) );
  INV_X1 U2046 ( .A(matrix_mul_2D_5__5__6_), .ZN(n8224) );
  INV_X1 U2047 ( .A(n61090), .ZN(n8225) );
  INV_X1 U2048 ( .A(n8225), .ZN(n8226) );
  BUF_X1 U2049 ( .A(n8230), .Z(n8227) );
  INV_X1 U2050 ( .A(matrix_mul_2D_5__5__5_), .ZN(n8228) );
  INV_X1 U2051 ( .A(n61100), .ZN(n8229) );
  INV_X1 U2052 ( .A(n8229), .ZN(n8230) );
  BUF_X1 U2053 ( .A(n8234), .Z(n8231) );
  INV_X1 U2054 ( .A(matrix_mul_2D_5__5__4_), .ZN(n8232) );
  INV_X1 U2055 ( .A(n61110), .ZN(n8233) );
  INV_X1 U2056 ( .A(n8233), .ZN(n8234) );
  BUF_X1 U2057 ( .A(n8238), .Z(n8235) );
  INV_X1 U2058 ( .A(matrix_mul_2D_5__5__3_), .ZN(n8236) );
  INV_X1 U2059 ( .A(n61120), .ZN(n8237) );
  INV_X1 U2060 ( .A(n8237), .ZN(n8238) );
  BUF_X1 U2061 ( .A(n8242), .Z(n8239) );
  INV_X1 U2062 ( .A(matrix_mul_2D_5__5__2_), .ZN(n8240) );
  INV_X1 U2063 ( .A(n61130), .ZN(n8241) );
  INV_X1 U2064 ( .A(n8241), .ZN(n8242) );
  BUF_X1 U2065 ( .A(n8246), .Z(n8243) );
  INV_X1 U2066 ( .A(matrix_mul_2D_5__5__1_), .ZN(n8244) );
  INV_X1 U2067 ( .A(n6114), .ZN(n8245) );
  INV_X1 U2068 ( .A(n8245), .ZN(n8246) );
  BUF_X1 U2069 ( .A(n8251), .Z(n8247) );
  INV_X1 U2070 ( .A(n2588), .ZN(n8248) );
  INV_X1 U2071 ( .A(n8248), .ZN(n8249) );
  INV_X1 U2072 ( .A(n6115), .ZN(n8250) );
  INV_X1 U2073 ( .A(n8250), .ZN(n8251) );
  BUF_X1 U2074 ( .A(n27606), .Z(n8252) );
  BUF_X1 U2075 ( .A(n27607), .Z(n8253) );
  BUF_X1 U2076 ( .A(n27608), .Z(n8254) );
  BUF_X1 U2077 ( .A(n27609), .Z(n8255) );
  BUF_X1 U2078 ( .A(n27610), .Z(n8256) );
  BUF_X1 U2079 ( .A(n27611), .Z(n8257) );
  BUF_X1 U2080 ( .A(n8261), .Z(n8258) );
  INV_X1 U2081 ( .A(matrix_mul_2D_5__4__14_), .ZN(n8259) );
  INV_X1 U2082 ( .A(n6086), .ZN(n8260) );
  INV_X1 U2083 ( .A(n8260), .ZN(n8261) );
  BUF_X1 U2084 ( .A(n8265), .Z(n8262) );
  INV_X1 U2085 ( .A(matrix_mul_2D_5__4__13_), .ZN(n8263) );
  INV_X1 U2086 ( .A(n6087), .ZN(n8264) );
  INV_X1 U2087 ( .A(n8264), .ZN(n8265) );
  BUF_X1 U2088 ( .A(n8269), .Z(n8266) );
  INV_X1 U2089 ( .A(matrix_mul_2D_5__4__12_), .ZN(n8267) );
  INV_X1 U2090 ( .A(n6088), .ZN(n8268) );
  INV_X1 U2091 ( .A(n8268), .ZN(n8269) );
  BUF_X1 U2092 ( .A(n8273), .Z(n8270) );
  INV_X1 U2093 ( .A(matrix_mul_2D_5__4__11_), .ZN(n8271) );
  INV_X1 U2094 ( .A(n6089), .ZN(n8272) );
  INV_X1 U2095 ( .A(n8272), .ZN(n8273) );
  BUF_X1 U2096 ( .A(n8277), .Z(n8274) );
  INV_X1 U2097 ( .A(matrix_mul_2D_5__4__10_), .ZN(n8275) );
  INV_X1 U2098 ( .A(n6090), .ZN(n8276) );
  INV_X1 U2099 ( .A(n8276), .ZN(n8277) );
  BUF_X1 U2100 ( .A(n8281), .Z(n8278) );
  INV_X1 U2101 ( .A(matrix_mul_2D_5__4__9_), .ZN(n8279) );
  INV_X1 U2102 ( .A(n6091), .ZN(n8280) );
  INV_X1 U2103 ( .A(n8280), .ZN(n8281) );
  BUF_X1 U2104 ( .A(n8285), .Z(n8282) );
  INV_X1 U2105 ( .A(matrix_mul_2D_5__4__8_), .ZN(n8283) );
  INV_X1 U2106 ( .A(n6092), .ZN(n8284) );
  INV_X1 U2107 ( .A(n8284), .ZN(n8285) );
  BUF_X1 U2108 ( .A(n8289), .Z(n8286) );
  INV_X1 U2109 ( .A(matrix_mul_2D_5__4__7_), .ZN(n8287) );
  INV_X1 U2110 ( .A(n60930), .ZN(n8288) );
  INV_X1 U2111 ( .A(n8288), .ZN(n8289) );
  BUF_X1 U2112 ( .A(n8293), .Z(n8290) );
  INV_X1 U2113 ( .A(matrix_mul_2D_5__4__6_), .ZN(n8291) );
  INV_X1 U2114 ( .A(n60940), .ZN(n8292) );
  INV_X1 U2115 ( .A(n8292), .ZN(n8293) );
  BUF_X1 U2116 ( .A(n8297), .Z(n8294) );
  INV_X1 U2117 ( .A(matrix_mul_2D_5__4__5_), .ZN(n8295) );
  INV_X1 U2118 ( .A(n60950), .ZN(n8296) );
  INV_X1 U2119 ( .A(n8296), .ZN(n8297) );
  BUF_X1 U2120 ( .A(n8301), .Z(n8298) );
  INV_X1 U2121 ( .A(matrix_mul_2D_5__4__4_), .ZN(n8299) );
  INV_X1 U2122 ( .A(n60960), .ZN(n8300) );
  INV_X1 U2123 ( .A(n8300), .ZN(n8301) );
  BUF_X1 U2124 ( .A(n8305), .Z(n8302) );
  INV_X1 U2125 ( .A(matrix_mul_2D_5__4__3_), .ZN(n8303) );
  INV_X1 U2126 ( .A(n60970), .ZN(n8304) );
  INV_X1 U2127 ( .A(n8304), .ZN(n8305) );
  BUF_X1 U2128 ( .A(n8309), .Z(n8306) );
  INV_X1 U2129 ( .A(matrix_mul_2D_5__4__2_), .ZN(n8307) );
  INV_X1 U2130 ( .A(n60980), .ZN(n8308) );
  INV_X1 U2131 ( .A(n8308), .ZN(n8309) );
  BUF_X1 U2132 ( .A(n8313), .Z(n8310) );
  INV_X1 U2133 ( .A(matrix_mul_2D_5__4__1_), .ZN(n8311) );
  INV_X1 U2134 ( .A(n60990), .ZN(n8312) );
  INV_X1 U2135 ( .A(n8312), .ZN(n8313) );
  BUF_X1 U2136 ( .A(n8318), .Z(n8314) );
  INV_X1 U2137 ( .A(n257300), .ZN(n8315) );
  INV_X1 U2138 ( .A(n8315), .ZN(n8316) );
  INV_X1 U2139 ( .A(n61000), .ZN(n8317) );
  INV_X1 U2140 ( .A(n8317), .ZN(n8318) );
  BUF_X1 U2141 ( .A(n27600), .Z(n8319) );
  BUF_X1 U2142 ( .A(n27601), .Z(n8320) );
  BUF_X1 U2143 ( .A(n27602), .Z(n8321) );
  BUF_X1 U2144 ( .A(n27603), .Z(n8322) );
  BUF_X1 U2145 ( .A(n27604), .Z(n8323) );
  BUF_X1 U2146 ( .A(n27605), .Z(n8324) );
  BUF_X1 U2147 ( .A(n8329), .Z(n8325) );
  INV_X1 U2148 ( .A(n2538), .ZN(n8326) );
  INV_X1 U2149 ( .A(n8326), .ZN(n8327) );
  INV_X1 U2150 ( .A(n60710), .ZN(n8328) );
  INV_X1 U2151 ( .A(n8328), .ZN(n8329) );
  BUF_X1 U2152 ( .A(n8334), .Z(n8330) );
  INV_X1 U2153 ( .A(n2539), .ZN(n8331) );
  INV_X1 U2154 ( .A(n8331), .ZN(n8332) );
  INV_X1 U2155 ( .A(n60720), .ZN(n8333) );
  INV_X1 U2156 ( .A(n8333), .ZN(n8334) );
  BUF_X1 U2157 ( .A(n8339), .Z(n8335) );
  INV_X1 U2158 ( .A(n2540), .ZN(n8336) );
  INV_X1 U2159 ( .A(n8336), .ZN(n8337) );
  INV_X1 U2160 ( .A(n60730), .ZN(n8338) );
  INV_X1 U2161 ( .A(n8338), .ZN(n8339) );
  BUF_X1 U2162 ( .A(n8344), .Z(n8340) );
  INV_X1 U2163 ( .A(n2541), .ZN(n8341) );
  INV_X1 U2164 ( .A(n8341), .ZN(n8342) );
  INV_X1 U2165 ( .A(n60740), .ZN(n8343) );
  INV_X1 U2166 ( .A(n8343), .ZN(n8344) );
  BUF_X1 U2167 ( .A(n8349), .Z(n8345) );
  INV_X1 U2168 ( .A(n2542), .ZN(n8346) );
  INV_X1 U2169 ( .A(n8346), .ZN(n8347) );
  INV_X1 U2170 ( .A(n60750), .ZN(n8348) );
  INV_X1 U2171 ( .A(n8348), .ZN(n8349) );
  BUF_X1 U2172 ( .A(n8354), .Z(n8350) );
  INV_X1 U2173 ( .A(n2543), .ZN(n8351) );
  INV_X1 U2174 ( .A(n8351), .ZN(n8352) );
  INV_X1 U2175 ( .A(n6076), .ZN(n8353) );
  INV_X1 U2176 ( .A(n8353), .ZN(n8354) );
  BUF_X1 U2177 ( .A(n8359), .Z(n8355) );
  INV_X1 U2178 ( .A(n2544), .ZN(n8356) );
  INV_X1 U2179 ( .A(n8356), .ZN(n8357) );
  INV_X1 U2180 ( .A(n6077), .ZN(n8358) );
  INV_X1 U2181 ( .A(n8358), .ZN(n8359) );
  BUF_X1 U2182 ( .A(n8364), .Z(n8360) );
  INV_X1 U2183 ( .A(n2545), .ZN(n8361) );
  INV_X1 U2184 ( .A(n8361), .ZN(n8362) );
  INV_X1 U2185 ( .A(n6078), .ZN(n8363) );
  INV_X1 U2186 ( .A(n8363), .ZN(n8364) );
  BUF_X1 U2187 ( .A(n8369), .Z(n8365) );
  INV_X1 U2188 ( .A(n2546), .ZN(n8366) );
  INV_X1 U2189 ( .A(n8366), .ZN(n8367) );
  INV_X1 U2190 ( .A(n6079), .ZN(n8368) );
  INV_X1 U2191 ( .A(n8368), .ZN(n8369) );
  BUF_X1 U2192 ( .A(n8374), .Z(n8370) );
  INV_X1 U2193 ( .A(n2547), .ZN(n8371) );
  INV_X1 U2194 ( .A(n8371), .ZN(n8372) );
  INV_X1 U2195 ( .A(n6080), .ZN(n8373) );
  INV_X1 U2196 ( .A(n8373), .ZN(n8374) );
  BUF_X1 U2197 ( .A(n8379), .Z(n8375) );
  INV_X1 U2198 ( .A(n2548), .ZN(n8376) );
  INV_X1 U2199 ( .A(n8376), .ZN(n8377) );
  INV_X1 U2200 ( .A(n6081), .ZN(n8378) );
  INV_X1 U2201 ( .A(n8378), .ZN(n8379) );
  BUF_X1 U2202 ( .A(n8384), .Z(n8380) );
  INV_X1 U2203 ( .A(n2549), .ZN(n8381) );
  INV_X1 U2204 ( .A(n8381), .ZN(n8382) );
  INV_X1 U2205 ( .A(n6082), .ZN(n8383) );
  INV_X1 U2206 ( .A(n8383), .ZN(n8384) );
  BUF_X1 U2207 ( .A(n8389), .Z(n8385) );
  INV_X1 U2208 ( .A(n2550), .ZN(n8386) );
  INV_X1 U2209 ( .A(n8386), .ZN(n8387) );
  INV_X1 U2210 ( .A(n6083), .ZN(n8388) );
  INV_X1 U2211 ( .A(n8388), .ZN(n8389) );
  BUF_X1 U2212 ( .A(n8394), .Z(n8390) );
  INV_X1 U2213 ( .A(n2551), .ZN(n8391) );
  INV_X1 U2214 ( .A(n8391), .ZN(n8392) );
  INV_X1 U2215 ( .A(n6084), .ZN(n8393) );
  INV_X1 U2216 ( .A(n8393), .ZN(n8394) );
  BUF_X1 U2217 ( .A(n8398), .Z(n8395) );
  INV_X1 U2218 ( .A(matrix_mul_2D_5__3__0_), .ZN(n8396) );
  INV_X1 U2219 ( .A(n6085), .ZN(n8397) );
  INV_X1 U2220 ( .A(n8397), .ZN(n8398) );
  BUF_X1 U2221 ( .A(n27594), .Z(n8399) );
  BUF_X1 U2222 ( .A(n27595), .Z(n8400) );
  BUF_X1 U2223 ( .A(n27596), .Z(n8401) );
  BUF_X1 U2224 ( .A(n27597), .Z(n8402) );
  BUF_X1 U2225 ( .A(n27598), .Z(n8403) );
  BUF_X1 U2226 ( .A(n27599), .Z(n8404) );
  BUF_X1 U2227 ( .A(n8409), .Z(n8405) );
  INV_X1 U2228 ( .A(n2523), .ZN(n8406) );
  INV_X1 U2229 ( .A(n8406), .ZN(n8407) );
  INV_X1 U2230 ( .A(n6056), .ZN(n8408) );
  INV_X1 U2231 ( .A(n8408), .ZN(n8409) );
  BUF_X1 U2232 ( .A(n8414), .Z(n8410) );
  INV_X1 U2233 ( .A(n2524), .ZN(n8411) );
  INV_X1 U2234 ( .A(n8411), .ZN(n8412) );
  INV_X1 U2235 ( .A(n6057), .ZN(n8413) );
  INV_X1 U2236 ( .A(n8413), .ZN(n8414) );
  BUF_X1 U2237 ( .A(n8419), .Z(n8415) );
  INV_X1 U2238 ( .A(n2525), .ZN(n8416) );
  INV_X1 U2239 ( .A(n8416), .ZN(n8417) );
  INV_X1 U2240 ( .A(n6058), .ZN(n8418) );
  INV_X1 U2241 ( .A(n8418), .ZN(n8419) );
  BUF_X1 U2242 ( .A(n8424), .Z(n8420) );
  INV_X1 U2243 ( .A(n2526), .ZN(n8421) );
  INV_X1 U2244 ( .A(n8421), .ZN(n8422) );
  INV_X1 U2245 ( .A(n6059), .ZN(n8423) );
  INV_X1 U2246 ( .A(n8423), .ZN(n8424) );
  BUF_X1 U2247 ( .A(n8429), .Z(n8425) );
  INV_X1 U2248 ( .A(n2527), .ZN(n8426) );
  INV_X1 U2249 ( .A(n8426), .ZN(n8427) );
  INV_X1 U2250 ( .A(n60600), .ZN(n8428) );
  INV_X1 U2251 ( .A(n8428), .ZN(n8429) );
  BUF_X1 U2252 ( .A(n8434), .Z(n8430) );
  INV_X1 U2253 ( .A(n2528), .ZN(n8431) );
  INV_X1 U2254 ( .A(n8431), .ZN(n8432) );
  INV_X1 U2255 ( .A(n60610), .ZN(n8433) );
  INV_X1 U2256 ( .A(n8433), .ZN(n8434) );
  BUF_X1 U2257 ( .A(n8439), .Z(n8435) );
  INV_X1 U2258 ( .A(n2529), .ZN(n8436) );
  INV_X1 U2259 ( .A(n8436), .ZN(n8437) );
  INV_X1 U2260 ( .A(n60620), .ZN(n8438) );
  INV_X1 U2261 ( .A(n8438), .ZN(n8439) );
  BUF_X1 U2262 ( .A(n8444), .Z(n8440) );
  INV_X1 U2263 ( .A(n2530), .ZN(n8441) );
  INV_X1 U2264 ( .A(n8441), .ZN(n8442) );
  INV_X1 U2265 ( .A(n60630), .ZN(n8443) );
  INV_X1 U2266 ( .A(n8443), .ZN(n8444) );
  BUF_X1 U2267 ( .A(n8449), .Z(n8445) );
  INV_X1 U2268 ( .A(n2531), .ZN(n8446) );
  INV_X1 U2269 ( .A(n8446), .ZN(n8447) );
  INV_X1 U2270 ( .A(n60640), .ZN(n8448) );
  INV_X1 U2271 ( .A(n8448), .ZN(n8449) );
  BUF_X1 U2272 ( .A(n8454), .Z(n8450) );
  INV_X1 U2273 ( .A(n2532), .ZN(n8451) );
  INV_X1 U2274 ( .A(n8451), .ZN(n8452) );
  INV_X1 U2275 ( .A(n60650), .ZN(n8453) );
  INV_X1 U2276 ( .A(n8453), .ZN(n8454) );
  BUF_X1 U2277 ( .A(n8459), .Z(n8455) );
  INV_X1 U2278 ( .A(n2533), .ZN(n8456) );
  INV_X1 U2279 ( .A(n8456), .ZN(n8457) );
  INV_X1 U2280 ( .A(n60660), .ZN(n8458) );
  INV_X1 U2281 ( .A(n8458), .ZN(n8459) );
  BUF_X1 U2282 ( .A(n8464), .Z(n8460) );
  INV_X1 U2283 ( .A(n2534), .ZN(n8461) );
  INV_X1 U2284 ( .A(n8461), .ZN(n8462) );
  INV_X1 U2285 ( .A(n60670), .ZN(n8463) );
  INV_X1 U2286 ( .A(n8463), .ZN(n8464) );
  BUF_X1 U2287 ( .A(n8469), .Z(n8465) );
  INV_X1 U2288 ( .A(n2535), .ZN(n8466) );
  INV_X1 U2289 ( .A(n8466), .ZN(n8467) );
  INV_X1 U2290 ( .A(n60680), .ZN(n8468) );
  INV_X1 U2291 ( .A(n8468), .ZN(n8469) );
  BUF_X1 U2292 ( .A(n8474), .Z(n8470) );
  INV_X1 U2293 ( .A(n2536), .ZN(n8471) );
  INV_X1 U2294 ( .A(n8471), .ZN(n8472) );
  INV_X1 U2295 ( .A(n60690), .ZN(n8473) );
  INV_X1 U2296 ( .A(n8473), .ZN(n8474) );
  BUF_X1 U2297 ( .A(n8478), .Z(n8475) );
  INV_X1 U2298 ( .A(matrix_mul_2D_5__2__0_), .ZN(n8476) );
  INV_X1 U2299 ( .A(n60700), .ZN(n8477) );
  INV_X1 U2300 ( .A(n8477), .ZN(n8478) );
  BUF_X1 U2301 ( .A(n27588), .Z(n8479) );
  BUF_X1 U2302 ( .A(n27589), .Z(n8480) );
  BUF_X1 U2303 ( .A(n27590), .Z(n8481) );
  BUF_X1 U2304 ( .A(n27591), .Z(n8482) );
  BUF_X1 U2305 ( .A(n27592), .Z(n8483) );
  BUF_X1 U2306 ( .A(n27593), .Z(n8484) );
  BUF_X1 U2307 ( .A(n8489), .Z(n8485) );
  INV_X1 U2308 ( .A(n2508), .ZN(n8486) );
  INV_X1 U2309 ( .A(n8486), .ZN(n8487) );
  INV_X1 U2310 ( .A(n6041), .ZN(n8488) );
  INV_X1 U2311 ( .A(n8488), .ZN(n8489) );
  BUF_X1 U2312 ( .A(n8494), .Z(n8490) );
  INV_X1 U2313 ( .A(n2509), .ZN(n8491) );
  INV_X1 U2314 ( .A(n8491), .ZN(n8492) );
  INV_X1 U2315 ( .A(n6042), .ZN(n8493) );
  INV_X1 U2316 ( .A(n8493), .ZN(n8494) );
  BUF_X1 U2317 ( .A(n8499), .Z(n8495) );
  INV_X1 U2318 ( .A(n2510), .ZN(n8496) );
  INV_X1 U2319 ( .A(n8496), .ZN(n8497) );
  INV_X1 U2320 ( .A(n6043), .ZN(n8498) );
  INV_X1 U2321 ( .A(n8498), .ZN(n8499) );
  BUF_X1 U2322 ( .A(n8504), .Z(n8500) );
  INV_X1 U2323 ( .A(n2511), .ZN(n8501) );
  INV_X1 U2324 ( .A(n8501), .ZN(n8502) );
  INV_X1 U2325 ( .A(n6044), .ZN(n8503) );
  INV_X1 U2326 ( .A(n8503), .ZN(n8504) );
  BUF_X1 U2327 ( .A(n8509), .Z(n8505) );
  INV_X1 U2328 ( .A(n2512), .ZN(n8506) );
  INV_X1 U2329 ( .A(n8506), .ZN(n8507) );
  INV_X1 U2330 ( .A(n6045), .ZN(n8508) );
  INV_X1 U2331 ( .A(n8508), .ZN(n8509) );
  BUF_X1 U2332 ( .A(n8514), .Z(n8510) );
  INV_X1 U2333 ( .A(n2513), .ZN(n8511) );
  INV_X1 U2334 ( .A(n8511), .ZN(n8512) );
  INV_X1 U2335 ( .A(n6046), .ZN(n8513) );
  INV_X1 U2336 ( .A(n8513), .ZN(n8514) );
  BUF_X1 U2337 ( .A(n8519), .Z(n8515) );
  INV_X1 U2338 ( .A(n2514), .ZN(n8516) );
  INV_X1 U2339 ( .A(n8516), .ZN(n8517) );
  INV_X1 U2340 ( .A(n6047), .ZN(n8518) );
  INV_X1 U2341 ( .A(n8518), .ZN(n8519) );
  BUF_X1 U2342 ( .A(n8524), .Z(n8520) );
  INV_X1 U2343 ( .A(n2515), .ZN(n8521) );
  INV_X1 U2344 ( .A(n8521), .ZN(n8522) );
  INV_X1 U2345 ( .A(n6048), .ZN(n8523) );
  INV_X1 U2346 ( .A(n8523), .ZN(n8524) );
  BUF_X1 U2347 ( .A(n8529), .Z(n8525) );
  INV_X1 U2348 ( .A(n2516), .ZN(n8526) );
  INV_X1 U2349 ( .A(n8526), .ZN(n8527) );
  INV_X1 U2350 ( .A(n6049), .ZN(n8528) );
  INV_X1 U2351 ( .A(n8528), .ZN(n8529) );
  BUF_X1 U2352 ( .A(n8534), .Z(n8530) );
  INV_X1 U2353 ( .A(n2517), .ZN(n8531) );
  INV_X1 U2354 ( .A(n8531), .ZN(n8532) );
  INV_X1 U2355 ( .A(n6050), .ZN(n8533) );
  INV_X1 U2356 ( .A(n8533), .ZN(n8534) );
  BUF_X1 U2357 ( .A(n8539), .Z(n8535) );
  INV_X1 U2358 ( .A(n2518), .ZN(n8536) );
  INV_X1 U2359 ( .A(n8536), .ZN(n8537) );
  INV_X1 U2360 ( .A(n6051), .ZN(n8538) );
  INV_X1 U2361 ( .A(n8538), .ZN(n8539) );
  BUF_X1 U2362 ( .A(n8544), .Z(n8540) );
  INV_X1 U2363 ( .A(n2519), .ZN(n8541) );
  INV_X1 U2364 ( .A(n8541), .ZN(n8542) );
  INV_X1 U2365 ( .A(n6052), .ZN(n8543) );
  INV_X1 U2366 ( .A(n8543), .ZN(n8544) );
  BUF_X1 U2367 ( .A(n8549), .Z(n8545) );
  INV_X1 U2368 ( .A(n2520), .ZN(n8546) );
  INV_X1 U2369 ( .A(n8546), .ZN(n8547) );
  INV_X1 U2370 ( .A(n6053), .ZN(n8548) );
  INV_X1 U2371 ( .A(n8548), .ZN(n8549) );
  BUF_X1 U2372 ( .A(n8554), .Z(n8550) );
  INV_X1 U2373 ( .A(n2521), .ZN(n8551) );
  INV_X1 U2374 ( .A(n8551), .ZN(n8552) );
  INV_X1 U2375 ( .A(n6054), .ZN(n8553) );
  INV_X1 U2376 ( .A(n8553), .ZN(n8554) );
  BUF_X1 U2377 ( .A(n8558), .Z(n8555) );
  INV_X1 U2378 ( .A(matrix_mul_2D_5__1__0_), .ZN(n8556) );
  INV_X1 U2379 ( .A(n6055), .ZN(n8557) );
  INV_X1 U2380 ( .A(n8557), .ZN(n8558) );
  BUF_X1 U2381 ( .A(n27582), .Z(n8559) );
  BUF_X1 U2382 ( .A(n27583), .Z(n8560) );
  BUF_X1 U2383 ( .A(n27584), .Z(n8561) );
  BUF_X1 U2384 ( .A(n27585), .Z(n8562) );
  BUF_X1 U2385 ( .A(n27586), .Z(n8563) );
  BUF_X1 U2386 ( .A(n27587), .Z(n8564) );
  BUF_X1 U2387 ( .A(n8569), .Z(n8565) );
  INV_X1 U2388 ( .A(n2493), .ZN(n8566) );
  INV_X1 U2389 ( .A(n8566), .ZN(n8567) );
  INV_X1 U2390 ( .A(n60260), .ZN(n8568) );
  INV_X1 U2391 ( .A(n8568), .ZN(n8569) );
  BUF_X1 U2392 ( .A(n8574), .Z(n8570) );
  INV_X1 U2393 ( .A(n2494), .ZN(n8571) );
  INV_X1 U2394 ( .A(n8571), .ZN(n8572) );
  INV_X1 U2395 ( .A(n60270), .ZN(n8573) );
  INV_X1 U2396 ( .A(n8573), .ZN(n8574) );
  BUF_X1 U2397 ( .A(n8579), .Z(n8575) );
  INV_X1 U2398 ( .A(n2495), .ZN(n8576) );
  INV_X1 U2399 ( .A(n8576), .ZN(n8577) );
  INV_X1 U2400 ( .A(n60280), .ZN(n8578) );
  INV_X1 U2401 ( .A(n8578), .ZN(n8579) );
  BUF_X1 U2402 ( .A(n8584), .Z(n8580) );
  INV_X1 U2403 ( .A(n2496), .ZN(n8581) );
  INV_X1 U2404 ( .A(n8581), .ZN(n8582) );
  INV_X1 U2405 ( .A(n60290), .ZN(n8583) );
  INV_X1 U2406 ( .A(n8583), .ZN(n8584) );
  BUF_X1 U2407 ( .A(n8589), .Z(n8585) );
  INV_X1 U2408 ( .A(n2497), .ZN(n8586) );
  INV_X1 U2409 ( .A(n8586), .ZN(n8587) );
  INV_X1 U2410 ( .A(n60300), .ZN(n8588) );
  INV_X1 U2411 ( .A(n8588), .ZN(n8589) );
  BUF_X1 U2412 ( .A(n8594), .Z(n8590) );
  INV_X1 U2413 ( .A(n2498), .ZN(n8591) );
  INV_X1 U2414 ( .A(n8591), .ZN(n8592) );
  INV_X1 U2415 ( .A(n60310), .ZN(n8593) );
  INV_X1 U2416 ( .A(n8593), .ZN(n8594) );
  BUF_X1 U2417 ( .A(n8599), .Z(n8595) );
  INV_X1 U2418 ( .A(n2499), .ZN(n8596) );
  INV_X1 U2419 ( .A(n8596), .ZN(n8597) );
  INV_X1 U2420 ( .A(n60320), .ZN(n8598) );
  INV_X1 U2421 ( .A(n8598), .ZN(n8599) );
  BUF_X1 U2422 ( .A(n8604), .Z(n8600) );
  INV_X1 U2423 ( .A(n2500), .ZN(n8601) );
  INV_X1 U2424 ( .A(n8601), .ZN(n8602) );
  INV_X1 U2425 ( .A(n60330), .ZN(n8603) );
  INV_X1 U2426 ( .A(n8603), .ZN(n8604) );
  BUF_X1 U2427 ( .A(n8609), .Z(n8605) );
  INV_X1 U2428 ( .A(n2501), .ZN(n8606) );
  INV_X1 U2429 ( .A(n8606), .ZN(n8607) );
  INV_X1 U2430 ( .A(n60340), .ZN(n8608) );
  INV_X1 U2431 ( .A(n8608), .ZN(n8609) );
  BUF_X1 U2432 ( .A(n8614), .Z(n8610) );
  INV_X1 U2433 ( .A(n2502), .ZN(n8611) );
  INV_X1 U2434 ( .A(n8611), .ZN(n8612) );
  INV_X1 U2435 ( .A(n6035), .ZN(n8613) );
  INV_X1 U2436 ( .A(n8613), .ZN(n8614) );
  BUF_X1 U2437 ( .A(n8619), .Z(n8615) );
  INV_X1 U2438 ( .A(n2503), .ZN(n8616) );
  INV_X1 U2439 ( .A(n8616), .ZN(n8617) );
  INV_X1 U2440 ( .A(n6036), .ZN(n8618) );
  INV_X1 U2441 ( .A(n8618), .ZN(n8619) );
  BUF_X1 U2442 ( .A(n8624), .Z(n8620) );
  INV_X1 U2443 ( .A(n2504), .ZN(n8621) );
  INV_X1 U2444 ( .A(n8621), .ZN(n8622) );
  INV_X1 U2445 ( .A(n6037), .ZN(n8623) );
  INV_X1 U2446 ( .A(n8623), .ZN(n8624) );
  BUF_X1 U2447 ( .A(n8629), .Z(n8625) );
  INV_X1 U2448 ( .A(n2505), .ZN(n8626) );
  INV_X1 U2449 ( .A(n8626), .ZN(n8627) );
  INV_X1 U2450 ( .A(n6038), .ZN(n8628) );
  INV_X1 U2451 ( .A(n8628), .ZN(n8629) );
  BUF_X1 U2452 ( .A(n8634), .Z(n8630) );
  INV_X1 U2453 ( .A(n2506), .ZN(n8631) );
  INV_X1 U2454 ( .A(n8631), .ZN(n8632) );
  INV_X1 U2455 ( .A(n6039), .ZN(n8633) );
  INV_X1 U2456 ( .A(n8633), .ZN(n8634) );
  BUF_X1 U2457 ( .A(n8638), .Z(n8635) );
  INV_X1 U2458 ( .A(matrix_mul_2D_5__0__0_), .ZN(n8636) );
  INV_X1 U2459 ( .A(n6040), .ZN(n8637) );
  INV_X1 U2460 ( .A(n8637), .ZN(n8638) );
  BUF_X1 U2461 ( .A(n27576), .Z(n8639) );
  BUF_X1 U2462 ( .A(n27577), .Z(n8640) );
  BUF_X1 U2463 ( .A(n27578), .Z(n8641) );
  BUF_X1 U2464 ( .A(n27579), .Z(n8642) );
  BUF_X1 U2465 ( .A(n27580), .Z(n8643) );
  BUF_X1 U2466 ( .A(n27581), .Z(n8644) );
  BUF_X1 U2467 ( .A(n8649), .Z(n8645) );
  INV_X1 U2468 ( .A(n2478), .ZN(n8646) );
  INV_X1 U2469 ( .A(n8646), .ZN(n8647) );
  INV_X1 U2470 ( .A(n6011), .ZN(n8648) );
  INV_X1 U2471 ( .A(n8648), .ZN(n8649) );
  BUF_X1 U2472 ( .A(n8654), .Z(n8650) );
  INV_X1 U2473 ( .A(n2479), .ZN(n8651) );
  INV_X1 U2474 ( .A(n8651), .ZN(n8652) );
  INV_X1 U2475 ( .A(n6012), .ZN(n8653) );
  INV_X1 U2476 ( .A(n8653), .ZN(n8654) );
  BUF_X1 U2477 ( .A(n8659), .Z(n8655) );
  INV_X1 U2478 ( .A(n2480), .ZN(n8656) );
  INV_X1 U2479 ( .A(n8656), .ZN(n8657) );
  INV_X1 U2480 ( .A(n6013), .ZN(n8658) );
  INV_X1 U2481 ( .A(n8658), .ZN(n8659) );
  BUF_X1 U2482 ( .A(n8664), .Z(n8660) );
  INV_X1 U2483 ( .A(n2481), .ZN(n8661) );
  INV_X1 U2484 ( .A(n8661), .ZN(n8662) );
  INV_X1 U2485 ( .A(n60140), .ZN(n8663) );
  INV_X1 U2486 ( .A(n8663), .ZN(n8664) );
  BUF_X1 U2487 ( .A(n8669), .Z(n8665) );
  INV_X1 U2488 ( .A(n2482), .ZN(n8666) );
  INV_X1 U2489 ( .A(n8666), .ZN(n8667) );
  INV_X1 U2490 ( .A(n60150), .ZN(n8668) );
  INV_X1 U2491 ( .A(n8668), .ZN(n8669) );
  BUF_X1 U2492 ( .A(n8674), .Z(n8670) );
  INV_X1 U2493 ( .A(n2483), .ZN(n8671) );
  INV_X1 U2494 ( .A(n8671), .ZN(n8672) );
  INV_X1 U2495 ( .A(n60160), .ZN(n8673) );
  INV_X1 U2496 ( .A(n8673), .ZN(n8674) );
  BUF_X1 U2497 ( .A(n8679), .Z(n8675) );
  INV_X1 U2498 ( .A(n2484), .ZN(n8676) );
  INV_X1 U2499 ( .A(n8676), .ZN(n8677) );
  INV_X1 U2500 ( .A(n60170), .ZN(n8678) );
  INV_X1 U2501 ( .A(n8678), .ZN(n8679) );
  BUF_X1 U2502 ( .A(n8684), .Z(n8680) );
  INV_X1 U2503 ( .A(n2485), .ZN(n8681) );
  INV_X1 U2504 ( .A(n8681), .ZN(n8682) );
  INV_X1 U2505 ( .A(n60180), .ZN(n8683) );
  INV_X1 U2506 ( .A(n8683), .ZN(n8684) );
  BUF_X1 U2507 ( .A(n8689), .Z(n8685) );
  INV_X1 U2508 ( .A(n2486), .ZN(n8686) );
  INV_X1 U2509 ( .A(n8686), .ZN(n8687) );
  INV_X1 U2510 ( .A(n60190), .ZN(n8688) );
  INV_X1 U2511 ( .A(n8688), .ZN(n8689) );
  BUF_X1 U2512 ( .A(n8694), .Z(n8690) );
  INV_X1 U2513 ( .A(n2487), .ZN(n8691) );
  INV_X1 U2514 ( .A(n8691), .ZN(n8692) );
  INV_X1 U2515 ( .A(n60200), .ZN(n8693) );
  INV_X1 U2516 ( .A(n8693), .ZN(n8694) );
  BUF_X1 U2517 ( .A(n8699), .Z(n8695) );
  INV_X1 U2518 ( .A(n2488), .ZN(n8696) );
  INV_X1 U2519 ( .A(n8696), .ZN(n8697) );
  INV_X1 U2520 ( .A(n60210), .ZN(n8698) );
  INV_X1 U2521 ( .A(n8698), .ZN(n8699) );
  BUF_X1 U2522 ( .A(n8704), .Z(n8700) );
  INV_X1 U2523 ( .A(n2489), .ZN(n8701) );
  INV_X1 U2524 ( .A(n8701), .ZN(n8702) );
  INV_X1 U2525 ( .A(n60220), .ZN(n8703) );
  INV_X1 U2526 ( .A(n8703), .ZN(n8704) );
  BUF_X1 U2527 ( .A(n8709), .Z(n8705) );
  INV_X1 U2528 ( .A(n2490), .ZN(n8706) );
  INV_X1 U2529 ( .A(n8706), .ZN(n8707) );
  INV_X1 U2530 ( .A(n60230), .ZN(n8708) );
  INV_X1 U2531 ( .A(n8708), .ZN(n8709) );
  BUF_X1 U2532 ( .A(n8714), .Z(n8710) );
  INV_X1 U2533 ( .A(n2491), .ZN(n8711) );
  INV_X1 U2534 ( .A(n8711), .ZN(n8712) );
  INV_X1 U2535 ( .A(n60240), .ZN(n8713) );
  INV_X1 U2536 ( .A(n8713), .ZN(n8714) );
  BUF_X1 U2537 ( .A(n8718), .Z(n8715) );
  INV_X1 U2538 ( .A(matrix_mul_2D_4__7__0_), .ZN(n8716) );
  INV_X1 U2539 ( .A(n60250), .ZN(n8717) );
  INV_X1 U2540 ( .A(n8717), .ZN(n8718) );
  BUF_X1 U2541 ( .A(n27570), .Z(n8719) );
  BUF_X1 U2542 ( .A(n27571), .Z(n8720) );
  BUF_X1 U2543 ( .A(n27572), .Z(n8721) );
  BUF_X1 U2544 ( .A(n27573), .Z(n8722) );
  BUF_X1 U2545 ( .A(n27574), .Z(n8723) );
  BUF_X1 U2546 ( .A(n27575), .Z(n8724) );
  BUF_X1 U2547 ( .A(n8729), .Z(n8725) );
  INV_X1 U2548 ( .A(n2463), .ZN(n8726) );
  INV_X1 U2549 ( .A(n8726), .ZN(n8727) );
  INV_X1 U2550 ( .A(n59960), .ZN(n8728) );
  INV_X1 U2551 ( .A(n8728), .ZN(n8729) );
  BUF_X1 U2552 ( .A(n8734), .Z(n8730) );
  INV_X1 U2553 ( .A(n2464), .ZN(n8731) );
  INV_X1 U2554 ( .A(n8731), .ZN(n8732) );
  INV_X1 U2555 ( .A(n5997), .ZN(n8733) );
  INV_X1 U2556 ( .A(n8733), .ZN(n8734) );
  BUF_X1 U2557 ( .A(n8739), .Z(n8735) );
  INV_X1 U2558 ( .A(n2465), .ZN(n8736) );
  INV_X1 U2559 ( .A(n8736), .ZN(n8737) );
  INV_X1 U2560 ( .A(n5998), .ZN(n8738) );
  INV_X1 U2561 ( .A(n8738), .ZN(n8739) );
  BUF_X1 U2562 ( .A(n8744), .Z(n8740) );
  INV_X1 U2563 ( .A(n2466), .ZN(n8741) );
  INV_X1 U2564 ( .A(n8741), .ZN(n8742) );
  INV_X1 U2565 ( .A(n5999), .ZN(n8743) );
  INV_X1 U2566 ( .A(n8743), .ZN(n8744) );
  BUF_X1 U2567 ( .A(n8749), .Z(n8745) );
  INV_X1 U2568 ( .A(n2467), .ZN(n8746) );
  INV_X1 U2569 ( .A(n8746), .ZN(n8747) );
  INV_X1 U2570 ( .A(n6000), .ZN(n8748) );
  INV_X1 U2571 ( .A(n8748), .ZN(n8749) );
  BUF_X1 U2572 ( .A(n8754), .Z(n8750) );
  INV_X1 U2573 ( .A(n2468), .ZN(n8751) );
  INV_X1 U2574 ( .A(n8751), .ZN(n8752) );
  INV_X1 U2575 ( .A(n6001), .ZN(n8753) );
  INV_X1 U2576 ( .A(n8753), .ZN(n8754) );
  BUF_X1 U2577 ( .A(n8759), .Z(n8755) );
  INV_X1 U2578 ( .A(n2469), .ZN(n8756) );
  INV_X1 U2579 ( .A(n8756), .ZN(n8757) );
  INV_X1 U2580 ( .A(n6002), .ZN(n8758) );
  INV_X1 U2581 ( .A(n8758), .ZN(n8759) );
  BUF_X1 U2582 ( .A(n8764), .Z(n8760) );
  INV_X1 U2583 ( .A(n2470), .ZN(n8761) );
  INV_X1 U2584 ( .A(n8761), .ZN(n8762) );
  INV_X1 U2585 ( .A(n6003), .ZN(n8763) );
  INV_X1 U2586 ( .A(n8763), .ZN(n8764) );
  BUF_X1 U2587 ( .A(n8769), .Z(n8765) );
  INV_X1 U2588 ( .A(n2471), .ZN(n8766) );
  INV_X1 U2589 ( .A(n8766), .ZN(n8767) );
  INV_X1 U2590 ( .A(n6004), .ZN(n8768) );
  INV_X1 U2591 ( .A(n8768), .ZN(n8769) );
  BUF_X1 U2592 ( .A(n8774), .Z(n8770) );
  INV_X1 U2593 ( .A(n2472), .ZN(n8771) );
  INV_X1 U2594 ( .A(n8771), .ZN(n8772) );
  INV_X1 U2595 ( .A(n6005), .ZN(n8773) );
  INV_X1 U2596 ( .A(n8773), .ZN(n8774) );
  BUF_X1 U2597 ( .A(n8779), .Z(n8775) );
  INV_X1 U2598 ( .A(n2473), .ZN(n8776) );
  INV_X1 U2599 ( .A(n8776), .ZN(n8777) );
  INV_X1 U2600 ( .A(n6006), .ZN(n8778) );
  INV_X1 U2601 ( .A(n8778), .ZN(n8779) );
  BUF_X1 U2602 ( .A(n8784), .Z(n8780) );
  INV_X1 U2603 ( .A(n2474), .ZN(n8781) );
  INV_X1 U2604 ( .A(n8781), .ZN(n8782) );
  INV_X1 U2605 ( .A(n6007), .ZN(n8783) );
  INV_X1 U2606 ( .A(n8783), .ZN(n8784) );
  BUF_X1 U2607 ( .A(n8789), .Z(n8785) );
  INV_X1 U2608 ( .A(n2475), .ZN(n8786) );
  INV_X1 U2609 ( .A(n8786), .ZN(n8787) );
  INV_X1 U2610 ( .A(n6008), .ZN(n8788) );
  INV_X1 U2611 ( .A(n8788), .ZN(n8789) );
  BUF_X1 U2612 ( .A(n8794), .Z(n8790) );
  INV_X1 U2613 ( .A(n2476), .ZN(n8791) );
  INV_X1 U2614 ( .A(n8791), .ZN(n8792) );
  INV_X1 U2615 ( .A(n6009), .ZN(n8793) );
  INV_X1 U2616 ( .A(n8793), .ZN(n8794) );
  BUF_X1 U2617 ( .A(n8798), .Z(n8795) );
  INV_X1 U2618 ( .A(matrix_mul_2D_4__6__0_), .ZN(n8796) );
  INV_X1 U2619 ( .A(n6010), .ZN(n8797) );
  INV_X1 U2620 ( .A(n8797), .ZN(n8798) );
  BUF_X1 U2621 ( .A(n27564), .Z(n8799) );
  BUF_X1 U2622 ( .A(n27565), .Z(n8800) );
  BUF_X1 U2623 ( .A(n27566), .Z(n8801) );
  BUF_X1 U2624 ( .A(n27567), .Z(n8802) );
  BUF_X1 U2625 ( .A(n27568), .Z(n8803) );
  BUF_X1 U2626 ( .A(n27569), .Z(n8804) );
  BUF_X1 U2627 ( .A(n8808), .Z(n8805) );
  INV_X1 U2628 ( .A(matrix_mul_2D_4__5__14_), .ZN(n8806) );
  INV_X1 U2629 ( .A(n59810), .ZN(n8807) );
  INV_X1 U2630 ( .A(n8807), .ZN(n8808) );
  BUF_X1 U2631 ( .A(n8812), .Z(n8809) );
  INV_X1 U2632 ( .A(matrix_mul_2D_4__5__13_), .ZN(n8810) );
  INV_X1 U2633 ( .A(n59820), .ZN(n8811) );
  INV_X1 U2634 ( .A(n8811), .ZN(n8812) );
  BUF_X1 U2635 ( .A(n8816), .Z(n8813) );
  INV_X1 U2636 ( .A(matrix_mul_2D_4__5__12_), .ZN(n8814) );
  INV_X1 U2637 ( .A(n59830), .ZN(n8815) );
  INV_X1 U2638 ( .A(n8815), .ZN(n8816) );
  BUF_X1 U2639 ( .A(n8820), .Z(n8817) );
  INV_X1 U2640 ( .A(matrix_mul_2D_4__5__11_), .ZN(n8818) );
  INV_X1 U2641 ( .A(n59840), .ZN(n8819) );
  INV_X1 U2642 ( .A(n8819), .ZN(n8820) );
  BUF_X1 U2643 ( .A(n8824), .Z(n8821) );
  INV_X1 U2644 ( .A(matrix_mul_2D_4__5__10_), .ZN(n8822) );
  INV_X1 U2645 ( .A(n59850), .ZN(n8823) );
  INV_X1 U2646 ( .A(n8823), .ZN(n8824) );
  BUF_X1 U2647 ( .A(n8828), .Z(n8825) );
  INV_X1 U2648 ( .A(matrix_mul_2D_4__5__9_), .ZN(n8826) );
  INV_X1 U2649 ( .A(n59860), .ZN(n8827) );
  INV_X1 U2650 ( .A(n8827), .ZN(n8828) );
  BUF_X1 U2651 ( .A(n8832), .Z(n8829) );
  INV_X1 U2652 ( .A(matrix_mul_2D_4__5__8_), .ZN(n8830) );
  INV_X1 U2653 ( .A(n59870), .ZN(n8831) );
  INV_X1 U2654 ( .A(n8831), .ZN(n8832) );
  BUF_X1 U2655 ( .A(n8836), .Z(n8833) );
  INV_X1 U2656 ( .A(matrix_mul_2D_4__5__7_), .ZN(n8834) );
  INV_X1 U2657 ( .A(n59880), .ZN(n8835) );
  INV_X1 U2658 ( .A(n8835), .ZN(n8836) );
  BUF_X1 U2659 ( .A(n8840), .Z(n8837) );
  INV_X1 U2660 ( .A(matrix_mul_2D_4__5__6_), .ZN(n8838) );
  INV_X1 U2661 ( .A(n59890), .ZN(n8839) );
  INV_X1 U2662 ( .A(n8839), .ZN(n8840) );
  BUF_X1 U2663 ( .A(n8844), .Z(n8841) );
  INV_X1 U2664 ( .A(matrix_mul_2D_4__5__5_), .ZN(n8842) );
  INV_X1 U2665 ( .A(n59900), .ZN(n8843) );
  INV_X1 U2666 ( .A(n8843), .ZN(n8844) );
  BUF_X1 U2667 ( .A(n8848), .Z(n8845) );
  INV_X1 U2668 ( .A(matrix_mul_2D_4__5__4_), .ZN(n8846) );
  INV_X1 U2669 ( .A(n59910), .ZN(n8847) );
  INV_X1 U2670 ( .A(n8847), .ZN(n8848) );
  BUF_X1 U2671 ( .A(n8852), .Z(n8849) );
  INV_X1 U2672 ( .A(matrix_mul_2D_4__5__3_), .ZN(n8850) );
  INV_X1 U2673 ( .A(n59920), .ZN(n8851) );
  INV_X1 U2674 ( .A(n8851), .ZN(n8852) );
  BUF_X1 U2675 ( .A(n8856), .Z(n8853) );
  INV_X1 U2676 ( .A(matrix_mul_2D_4__5__2_), .ZN(n8854) );
  INV_X1 U2677 ( .A(n59930), .ZN(n8855) );
  INV_X1 U2678 ( .A(n8855), .ZN(n8856) );
  BUF_X1 U2679 ( .A(n8860), .Z(n8857) );
  INV_X1 U2680 ( .A(matrix_mul_2D_4__5__1_), .ZN(n8858) );
  INV_X1 U2681 ( .A(n59940), .ZN(n8859) );
  INV_X1 U2682 ( .A(n8859), .ZN(n8860) );
  BUF_X1 U2683 ( .A(n8865), .Z(n8861) );
  INV_X1 U2684 ( .A(n2462), .ZN(n8862) );
  INV_X1 U2685 ( .A(n8862), .ZN(n8863) );
  INV_X1 U2686 ( .A(n59950), .ZN(n8864) );
  INV_X1 U2687 ( .A(n8864), .ZN(n8865) );
  BUF_X1 U2688 ( .A(n27558), .Z(n8866) );
  BUF_X1 U2689 ( .A(n27559), .Z(n8867) );
  BUF_X1 U2690 ( .A(n27560), .Z(n8868) );
  BUF_X1 U2691 ( .A(n27561), .Z(n8869) );
  BUF_X1 U2692 ( .A(n27562), .Z(n8870) );
  BUF_X1 U2693 ( .A(n27563), .Z(n8871) );
  BUF_X1 U2694 ( .A(n8875), .Z(n8872) );
  INV_X1 U2695 ( .A(matrix_mul_2D_4__4__14_), .ZN(n8873) );
  INV_X1 U2696 ( .A(n5966), .ZN(n8874) );
  INV_X1 U2697 ( .A(n8874), .ZN(n8875) );
  BUF_X1 U2698 ( .A(n8879), .Z(n8876) );
  INV_X1 U2699 ( .A(matrix_mul_2D_4__4__13_), .ZN(n8877) );
  INV_X1 U2700 ( .A(n5967), .ZN(n8878) );
  INV_X1 U2701 ( .A(n8878), .ZN(n8879) );
  BUF_X1 U2702 ( .A(n8883), .Z(n8880) );
  INV_X1 U2703 ( .A(matrix_mul_2D_4__4__12_), .ZN(n8881) );
  INV_X1 U2704 ( .A(n5968), .ZN(n8882) );
  INV_X1 U2705 ( .A(n8882), .ZN(n8883) );
  BUF_X1 U2706 ( .A(n8887), .Z(n8884) );
  INV_X1 U2707 ( .A(matrix_mul_2D_4__4__11_), .ZN(n8885) );
  INV_X1 U2708 ( .A(n5969), .ZN(n8886) );
  INV_X1 U2709 ( .A(n8886), .ZN(n8887) );
  BUF_X1 U2710 ( .A(n8891), .Z(n8888) );
  INV_X1 U2711 ( .A(matrix_mul_2D_4__4__10_), .ZN(n8889) );
  INV_X1 U2712 ( .A(n5970), .ZN(n8890) );
  INV_X1 U2713 ( .A(n8890), .ZN(n8891) );
  BUF_X1 U2714 ( .A(n8895), .Z(n8892) );
  INV_X1 U2715 ( .A(matrix_mul_2D_4__4__9_), .ZN(n8893) );
  INV_X1 U2716 ( .A(n5971), .ZN(n8894) );
  INV_X1 U2717 ( .A(n8894), .ZN(n8895) );
  BUF_X1 U2718 ( .A(n8899), .Z(n8896) );
  INV_X1 U2719 ( .A(matrix_mul_2D_4__4__8_), .ZN(n8897) );
  INV_X1 U2720 ( .A(n5972), .ZN(n8898) );
  INV_X1 U2721 ( .A(n8898), .ZN(n8899) );
  BUF_X1 U2722 ( .A(n8903), .Z(n8900) );
  INV_X1 U2723 ( .A(matrix_mul_2D_4__4__7_), .ZN(n8901) );
  INV_X1 U2724 ( .A(n5973), .ZN(n8902) );
  INV_X1 U2725 ( .A(n8902), .ZN(n8903) );
  BUF_X1 U2726 ( .A(n8907), .Z(n8904) );
  INV_X1 U2727 ( .A(matrix_mul_2D_4__4__6_), .ZN(n8905) );
  INV_X1 U2728 ( .A(n5974), .ZN(n8906) );
  INV_X1 U2729 ( .A(n8906), .ZN(n8907) );
  BUF_X1 U2730 ( .A(n8911), .Z(n8908) );
  INV_X1 U2731 ( .A(matrix_mul_2D_4__4__5_), .ZN(n8909) );
  INV_X1 U2732 ( .A(n5975), .ZN(n8910) );
  INV_X1 U2733 ( .A(n8910), .ZN(n8911) );
  BUF_X1 U2734 ( .A(n8915), .Z(n8912) );
  INV_X1 U2735 ( .A(matrix_mul_2D_4__4__4_), .ZN(n8913) );
  INV_X1 U2736 ( .A(n5976), .ZN(n8914) );
  INV_X1 U2737 ( .A(n8914), .ZN(n8915) );
  BUF_X1 U2738 ( .A(n8919), .Z(n8916) );
  INV_X1 U2739 ( .A(matrix_mul_2D_4__4__3_), .ZN(n8917) );
  INV_X1 U2740 ( .A(n5977), .ZN(n8918) );
  INV_X1 U2741 ( .A(n8918), .ZN(n8919) );
  BUF_X1 U2742 ( .A(n8923), .Z(n8920) );
  INV_X1 U2743 ( .A(matrix_mul_2D_4__4__2_), .ZN(n8921) );
  INV_X1 U2744 ( .A(n5978), .ZN(n8922) );
  INV_X1 U2745 ( .A(n8922), .ZN(n8923) );
  BUF_X1 U2746 ( .A(n8927), .Z(n8924) );
  INV_X1 U2747 ( .A(matrix_mul_2D_4__4__1_), .ZN(n8925) );
  INV_X1 U2748 ( .A(n5979), .ZN(n8926) );
  INV_X1 U2749 ( .A(n8926), .ZN(n8927) );
  BUF_X1 U2750 ( .A(n8932), .Z(n8928) );
  INV_X1 U2751 ( .A(n2447), .ZN(n8929) );
  INV_X1 U2752 ( .A(n8929), .ZN(n8930) );
  INV_X1 U2753 ( .A(n5980), .ZN(n8931) );
  INV_X1 U2754 ( .A(n8931), .ZN(n8932) );
  BUF_X1 U2755 ( .A(n27552), .Z(n8933) );
  BUF_X1 U2756 ( .A(n27553), .Z(n8934) );
  BUF_X1 U2757 ( .A(n27554), .Z(n8935) );
  BUF_X1 U2758 ( .A(n27555), .Z(n8936) );
  BUF_X1 U2759 ( .A(n27556), .Z(n8937) );
  BUF_X1 U2760 ( .A(n27557), .Z(n8938) );
  BUF_X1 U2761 ( .A(n8943), .Z(n8939) );
  INV_X1 U2762 ( .A(n2412), .ZN(n8940) );
  INV_X1 U2763 ( .A(n8940), .ZN(n8941) );
  INV_X1 U2764 ( .A(n5951), .ZN(n8942) );
  INV_X1 U2765 ( .A(n8942), .ZN(n8943) );
  BUF_X1 U2766 ( .A(n8948), .Z(n8944) );
  INV_X1 U2767 ( .A(n2413), .ZN(n8945) );
  INV_X1 U2768 ( .A(n8945), .ZN(n8946) );
  INV_X1 U2769 ( .A(n5952), .ZN(n8947) );
  INV_X1 U2770 ( .A(n8947), .ZN(n8948) );
  BUF_X1 U2771 ( .A(n8953), .Z(n8949) );
  INV_X1 U2772 ( .A(n2414), .ZN(n8950) );
  INV_X1 U2773 ( .A(n8950), .ZN(n8951) );
  INV_X1 U2774 ( .A(n5953), .ZN(n8952) );
  INV_X1 U2775 ( .A(n8952), .ZN(n8953) );
  BUF_X1 U2776 ( .A(n8958), .Z(n8954) );
  INV_X1 U2777 ( .A(n2415), .ZN(n8955) );
  INV_X1 U2778 ( .A(n8955), .ZN(n8956) );
  INV_X1 U2779 ( .A(n5954), .ZN(n8957) );
  INV_X1 U2780 ( .A(n8957), .ZN(n8958) );
  BUF_X1 U2781 ( .A(n8963), .Z(n8959) );
  INV_X1 U2782 ( .A(n2416), .ZN(n8960) );
  INV_X1 U2783 ( .A(n8960), .ZN(n8961) );
  INV_X1 U2784 ( .A(n5955), .ZN(n8962) );
  INV_X1 U2785 ( .A(n8962), .ZN(n8963) );
  BUF_X1 U2786 ( .A(n8968), .Z(n8964) );
  INV_X1 U2787 ( .A(n2417), .ZN(n8965) );
  INV_X1 U2788 ( .A(n8965), .ZN(n8966) );
  INV_X1 U2789 ( .A(n5956), .ZN(n8967) );
  INV_X1 U2790 ( .A(n8967), .ZN(n8968) );
  BUF_X1 U2791 ( .A(n8973), .Z(n8969) );
  INV_X1 U2792 ( .A(n2418), .ZN(n8970) );
  INV_X1 U2793 ( .A(n8970), .ZN(n8971) );
  INV_X1 U2794 ( .A(n5957), .ZN(n8972) );
  INV_X1 U2795 ( .A(n8972), .ZN(n8973) );
  BUF_X1 U2796 ( .A(n8978), .Z(n8974) );
  INV_X1 U2797 ( .A(n2419), .ZN(n8975) );
  INV_X1 U2798 ( .A(n8975), .ZN(n8976) );
  INV_X1 U2799 ( .A(n5958), .ZN(n8977) );
  INV_X1 U2800 ( .A(n8977), .ZN(n8978) );
  BUF_X1 U2801 ( .A(n8983), .Z(n8979) );
  INV_X1 U2802 ( .A(n2420), .ZN(n8980) );
  INV_X1 U2803 ( .A(n8980), .ZN(n8981) );
  INV_X1 U2804 ( .A(n5959), .ZN(n8982) );
  INV_X1 U2805 ( .A(n8982), .ZN(n8983) );
  BUF_X1 U2806 ( .A(n8988), .Z(n8984) );
  INV_X1 U2807 ( .A(n2421), .ZN(n8985) );
  INV_X1 U2808 ( .A(n8985), .ZN(n8986) );
  INV_X1 U2809 ( .A(n5960), .ZN(n8987) );
  INV_X1 U2810 ( .A(n8987), .ZN(n8988) );
  BUF_X1 U2811 ( .A(n8993), .Z(n8989) );
  INV_X1 U2812 ( .A(n2422), .ZN(n8990) );
  INV_X1 U2813 ( .A(n8990), .ZN(n8991) );
  INV_X1 U2814 ( .A(n5961), .ZN(n8992) );
  INV_X1 U2815 ( .A(n8992), .ZN(n8993) );
  BUF_X1 U2816 ( .A(n8998), .Z(n8994) );
  INV_X1 U2817 ( .A(n2423), .ZN(n8995) );
  INV_X1 U2818 ( .A(n8995), .ZN(n8996) );
  INV_X1 U2819 ( .A(n5962), .ZN(n8997) );
  INV_X1 U2820 ( .A(n8997), .ZN(n8998) );
  BUF_X1 U2821 ( .A(n9003), .Z(n8999) );
  INV_X1 U2822 ( .A(n2424), .ZN(n9000) );
  INV_X1 U2823 ( .A(n9000), .ZN(n9001) );
  INV_X1 U2824 ( .A(n5963), .ZN(n9002) );
  INV_X1 U2825 ( .A(n9002), .ZN(n9003) );
  BUF_X1 U2826 ( .A(n9008), .Z(n9004) );
  INV_X1 U2827 ( .A(n2425), .ZN(n9005) );
  INV_X1 U2828 ( .A(n9005), .ZN(n9006) );
  INV_X1 U2829 ( .A(n5964), .ZN(n9007) );
  INV_X1 U2830 ( .A(n9007), .ZN(n9008) );
  BUF_X1 U2831 ( .A(n9012), .Z(n9009) );
  INV_X1 U2832 ( .A(matrix_mul_2D_4__3__0_), .ZN(n9010) );
  INV_X1 U2833 ( .A(n5965), .ZN(n9011) );
  INV_X1 U2834 ( .A(n9011), .ZN(n9012) );
  BUF_X1 U2835 ( .A(n27546), .Z(n9013) );
  BUF_X1 U2836 ( .A(n27547), .Z(n9014) );
  BUF_X1 U2837 ( .A(n27548), .Z(n9015) );
  BUF_X1 U2838 ( .A(n27549), .Z(n9016) );
  BUF_X1 U2839 ( .A(n27550), .Z(n9017) );
  BUF_X1 U2840 ( .A(n27551), .Z(n9018) );
  BUF_X1 U2841 ( .A(n9023), .Z(n9019) );
  INV_X1 U2842 ( .A(n2397), .ZN(n9020) );
  INV_X1 U2843 ( .A(n9020), .ZN(n9021) );
  INV_X1 U2844 ( .A(n59360), .ZN(n9022) );
  INV_X1 U2845 ( .A(n9022), .ZN(n9023) );
  BUF_X1 U2846 ( .A(n9028), .Z(n9024) );
  INV_X1 U2847 ( .A(n2398), .ZN(n9025) );
  INV_X1 U2848 ( .A(n9025), .ZN(n9026) );
  INV_X1 U2849 ( .A(n59370), .ZN(n9027) );
  INV_X1 U2850 ( .A(n9027), .ZN(n9028) );
  BUF_X1 U2851 ( .A(n9033), .Z(n9029) );
  INV_X1 U2852 ( .A(n2399), .ZN(n9030) );
  INV_X1 U2853 ( .A(n9030), .ZN(n9031) );
  INV_X1 U2854 ( .A(n59380), .ZN(n9032) );
  INV_X1 U2855 ( .A(n9032), .ZN(n9033) );
  BUF_X1 U2856 ( .A(n9038), .Z(n9034) );
  INV_X1 U2857 ( .A(n2400), .ZN(n9035) );
  INV_X1 U2858 ( .A(n9035), .ZN(n9036) );
  INV_X1 U2859 ( .A(n59390), .ZN(n9037) );
  INV_X1 U2860 ( .A(n9037), .ZN(n9038) );
  BUF_X1 U2861 ( .A(n9043), .Z(n9039) );
  INV_X1 U2862 ( .A(n2401), .ZN(n9040) );
  INV_X1 U2863 ( .A(n9040), .ZN(n9041) );
  INV_X1 U2864 ( .A(n59400), .ZN(n9042) );
  INV_X1 U2865 ( .A(n9042), .ZN(n9043) );
  BUF_X1 U2866 ( .A(n9048), .Z(n9044) );
  INV_X1 U2867 ( .A(n2402), .ZN(n9045) );
  INV_X1 U2868 ( .A(n9045), .ZN(n9046) );
  INV_X1 U2869 ( .A(n59410), .ZN(n9047) );
  INV_X1 U2870 ( .A(n9047), .ZN(n9048) );
  BUF_X1 U2871 ( .A(n9053), .Z(n9049) );
  INV_X1 U2872 ( .A(n2403), .ZN(n9050) );
  INV_X1 U2873 ( .A(n9050), .ZN(n9051) );
  INV_X1 U2874 ( .A(n59420), .ZN(n9052) );
  INV_X1 U2875 ( .A(n9052), .ZN(n9053) );
  BUF_X1 U2876 ( .A(n9058), .Z(n9054) );
  INV_X1 U2877 ( .A(n2404), .ZN(n9055) );
  INV_X1 U2878 ( .A(n9055), .ZN(n9056) );
  INV_X1 U2879 ( .A(n59430), .ZN(n9057) );
  INV_X1 U2880 ( .A(n9057), .ZN(n9058) );
  BUF_X1 U2881 ( .A(n9063), .Z(n9059) );
  INV_X1 U2882 ( .A(n2405), .ZN(n9060) );
  INV_X1 U2883 ( .A(n9060), .ZN(n9061) );
  INV_X1 U2884 ( .A(n59440), .ZN(n9062) );
  INV_X1 U2885 ( .A(n9062), .ZN(n9063) );
  BUF_X1 U2886 ( .A(n9068), .Z(n9064) );
  INV_X1 U2887 ( .A(n2406), .ZN(n9065) );
  INV_X1 U2888 ( .A(n9065), .ZN(n9066) );
  INV_X1 U2889 ( .A(n59450), .ZN(n9067) );
  INV_X1 U2890 ( .A(n9067), .ZN(n9068) );
  BUF_X1 U2891 ( .A(n9073), .Z(n9069) );
  INV_X1 U2892 ( .A(n2407), .ZN(n9070) );
  INV_X1 U2893 ( .A(n9070), .ZN(n9071) );
  INV_X1 U2894 ( .A(n5946), .ZN(n9072) );
  INV_X1 U2895 ( .A(n9072), .ZN(n9073) );
  BUF_X1 U2896 ( .A(n9078), .Z(n9074) );
  INV_X1 U2897 ( .A(n2408), .ZN(n9075) );
  INV_X1 U2898 ( .A(n9075), .ZN(n9076) );
  INV_X1 U2899 ( .A(n5947), .ZN(n9077) );
  INV_X1 U2900 ( .A(n9077), .ZN(n9078) );
  BUF_X1 U2901 ( .A(n9083), .Z(n9079) );
  INV_X1 U2902 ( .A(n2409), .ZN(n9080) );
  INV_X1 U2903 ( .A(n9080), .ZN(n9081) );
  INV_X1 U2904 ( .A(n5948), .ZN(n9082) );
  INV_X1 U2905 ( .A(n9082), .ZN(n9083) );
  BUF_X1 U2906 ( .A(n9088), .Z(n9084) );
  INV_X1 U2907 ( .A(n2410), .ZN(n9085) );
  INV_X1 U2908 ( .A(n9085), .ZN(n9086) );
  INV_X1 U2909 ( .A(n5949), .ZN(n9087) );
  INV_X1 U2910 ( .A(n9087), .ZN(n9088) );
  BUF_X1 U2911 ( .A(n9092), .Z(n9089) );
  INV_X1 U2912 ( .A(matrix_mul_2D_4__2__0_), .ZN(n9090) );
  INV_X1 U2913 ( .A(n5950), .ZN(n9091) );
  INV_X1 U2914 ( .A(n9091), .ZN(n9092) );
  BUF_X1 U2915 ( .A(n27540), .Z(n9093) );
  BUF_X1 U2916 ( .A(n27541), .Z(n9094) );
  BUF_X1 U2917 ( .A(n27542), .Z(n9095) );
  BUF_X1 U2918 ( .A(n27543), .Z(n9096) );
  BUF_X1 U2919 ( .A(n27544), .Z(n9097) );
  BUF_X1 U2920 ( .A(n27545), .Z(n9098) );
  BUF_X1 U2921 ( .A(n9103), .Z(n9099) );
  INV_X1 U2922 ( .A(n2382), .ZN(n9100) );
  INV_X1 U2923 ( .A(n9100), .ZN(n9101) );
  INV_X1 U2924 ( .A(n5921), .ZN(n9102) );
  INV_X1 U2925 ( .A(n9102), .ZN(n9103) );
  BUF_X1 U2926 ( .A(n9108), .Z(n9104) );
  INV_X1 U2927 ( .A(n2383), .ZN(n9105) );
  INV_X1 U2928 ( .A(n9105), .ZN(n9106) );
  INV_X1 U2929 ( .A(n5922), .ZN(n9107) );
  INV_X1 U2930 ( .A(n9107), .ZN(n9108) );
  BUF_X1 U2931 ( .A(n9113), .Z(n9109) );
  INV_X1 U2932 ( .A(n2384), .ZN(n9110) );
  INV_X1 U2933 ( .A(n9110), .ZN(n9111) );
  INV_X1 U2934 ( .A(n5923), .ZN(n9112) );
  INV_X1 U2935 ( .A(n9112), .ZN(n9113) );
  BUF_X1 U2936 ( .A(n9118), .Z(n9114) );
  INV_X1 U2937 ( .A(n2385), .ZN(n9115) );
  INV_X1 U2938 ( .A(n9115), .ZN(n9116) );
  INV_X1 U2939 ( .A(n5924), .ZN(n9117) );
  INV_X1 U2940 ( .A(n9117), .ZN(n9118) );
  BUF_X1 U2941 ( .A(n9123), .Z(n9119) );
  INV_X1 U2942 ( .A(n2386), .ZN(n9120) );
  INV_X1 U2943 ( .A(n9120), .ZN(n9121) );
  INV_X1 U2944 ( .A(n59250), .ZN(n9122) );
  INV_X1 U2945 ( .A(n9122), .ZN(n9123) );
  BUF_X1 U2946 ( .A(n9128), .Z(n9124) );
  INV_X1 U2947 ( .A(n2387), .ZN(n9125) );
  INV_X1 U2948 ( .A(n9125), .ZN(n9126) );
  INV_X1 U2949 ( .A(n59260), .ZN(n9127) );
  INV_X1 U2950 ( .A(n9127), .ZN(n9128) );
  BUF_X1 U2951 ( .A(n9133), .Z(n9129) );
  INV_X1 U2952 ( .A(n2388), .ZN(n9130) );
  INV_X1 U2953 ( .A(n9130), .ZN(n9131) );
  INV_X1 U2954 ( .A(n59270), .ZN(n9132) );
  INV_X1 U2955 ( .A(n9132), .ZN(n9133) );
  BUF_X1 U2956 ( .A(n9138), .Z(n9134) );
  INV_X1 U2957 ( .A(n2389), .ZN(n9135) );
  INV_X1 U2958 ( .A(n9135), .ZN(n9136) );
  INV_X1 U2959 ( .A(n59280), .ZN(n9137) );
  INV_X1 U2960 ( .A(n9137), .ZN(n9138) );
  BUF_X1 U2961 ( .A(n9143), .Z(n9139) );
  INV_X1 U2962 ( .A(n2390), .ZN(n9140) );
  INV_X1 U2963 ( .A(n9140), .ZN(n9141) );
  INV_X1 U2964 ( .A(n59290), .ZN(n9142) );
  INV_X1 U2965 ( .A(n9142), .ZN(n9143) );
  BUF_X1 U2966 ( .A(n9148), .Z(n9144) );
  INV_X1 U2967 ( .A(n2391), .ZN(n9145) );
  INV_X1 U2968 ( .A(n9145), .ZN(n9146) );
  INV_X1 U2969 ( .A(n59300), .ZN(n9147) );
  INV_X1 U2970 ( .A(n9147), .ZN(n9148) );
  BUF_X1 U2971 ( .A(n9153), .Z(n9149) );
  INV_X1 U2972 ( .A(n2392), .ZN(n9150) );
  INV_X1 U2973 ( .A(n9150), .ZN(n9151) );
  INV_X1 U2974 ( .A(n59310), .ZN(n9152) );
  INV_X1 U2975 ( .A(n9152), .ZN(n9153) );
  BUF_X1 U2976 ( .A(n9158), .Z(n9154) );
  INV_X1 U2977 ( .A(n2393), .ZN(n9155) );
  INV_X1 U2978 ( .A(n9155), .ZN(n9156) );
  INV_X1 U2979 ( .A(n59320), .ZN(n9157) );
  INV_X1 U2980 ( .A(n9157), .ZN(n9158) );
  BUF_X1 U2981 ( .A(n9163), .Z(n9159) );
  INV_X1 U2982 ( .A(n2394), .ZN(n9160) );
  INV_X1 U2983 ( .A(n9160), .ZN(n9161) );
  INV_X1 U2984 ( .A(n59330), .ZN(n9162) );
  INV_X1 U2985 ( .A(n9162), .ZN(n9163) );
  BUF_X1 U2986 ( .A(n9168), .Z(n9164) );
  INV_X1 U2987 ( .A(n2395), .ZN(n9165) );
  INV_X1 U2988 ( .A(n9165), .ZN(n9166) );
  INV_X1 U2989 ( .A(n59340), .ZN(n9167) );
  INV_X1 U2990 ( .A(n9167), .ZN(n9168) );
  BUF_X1 U2991 ( .A(n9172), .Z(n9169) );
  INV_X1 U2992 ( .A(matrix_mul_2D_4__1__0_), .ZN(n9170) );
  INV_X1 U2993 ( .A(n59350), .ZN(n9171) );
  INV_X1 U2994 ( .A(n9171), .ZN(n9172) );
  BUF_X1 U2995 ( .A(n27534), .Z(n9173) );
  BUF_X1 U2996 ( .A(n27535), .Z(n9174) );
  BUF_X1 U2997 ( .A(n27536), .Z(n9175) );
  BUF_X1 U2998 ( .A(n27537), .Z(n9176) );
  BUF_X1 U2999 ( .A(n27538), .Z(n9177) );
  BUF_X1 U3000 ( .A(n27539), .Z(n9178) );
  BUF_X1 U3001 ( .A(n9183), .Z(n9179) );
  INV_X1 U3002 ( .A(n2367), .ZN(n9180) );
  INV_X1 U3003 ( .A(n9180), .ZN(n9181) );
  INV_X1 U3004 ( .A(n59060), .ZN(n9182) );
  INV_X1 U3005 ( .A(n9182), .ZN(n9183) );
  BUF_X1 U3006 ( .A(n9188), .Z(n9184) );
  INV_X1 U3007 ( .A(n2368), .ZN(n9185) );
  INV_X1 U3008 ( .A(n9185), .ZN(n9186) );
  INV_X1 U3009 ( .A(n59070), .ZN(n9187) );
  INV_X1 U3010 ( .A(n9187), .ZN(n9188) );
  BUF_X1 U3011 ( .A(n9193), .Z(n9189) );
  INV_X1 U3012 ( .A(n2369), .ZN(n9190) );
  INV_X1 U3013 ( .A(n9190), .ZN(n9191) );
  INV_X1 U3014 ( .A(n5908), .ZN(n9192) );
  INV_X1 U3015 ( .A(n9192), .ZN(n9193) );
  BUF_X1 U3016 ( .A(n9198), .Z(n9194) );
  INV_X1 U3017 ( .A(n2370), .ZN(n9195) );
  INV_X1 U3018 ( .A(n9195), .ZN(n9196) );
  INV_X1 U3019 ( .A(n5909), .ZN(n9197) );
  INV_X1 U3020 ( .A(n9197), .ZN(n9198) );
  BUF_X1 U3021 ( .A(n9203), .Z(n9199) );
  INV_X1 U3022 ( .A(n2371), .ZN(n9200) );
  INV_X1 U3023 ( .A(n9200), .ZN(n9201) );
  INV_X1 U3024 ( .A(n5910), .ZN(n9202) );
  INV_X1 U3025 ( .A(n9202), .ZN(n9203) );
  BUF_X1 U3026 ( .A(n9208), .Z(n9204) );
  INV_X1 U3027 ( .A(n2372), .ZN(n9205) );
  INV_X1 U3028 ( .A(n9205), .ZN(n9206) );
  INV_X1 U3029 ( .A(n5911), .ZN(n9207) );
  INV_X1 U3030 ( .A(n9207), .ZN(n9208) );
  BUF_X1 U3031 ( .A(n9213), .Z(n9209) );
  INV_X1 U3032 ( .A(n2373), .ZN(n9210) );
  INV_X1 U3033 ( .A(n9210), .ZN(n9211) );
  INV_X1 U3034 ( .A(n5912), .ZN(n9212) );
  INV_X1 U3035 ( .A(n9212), .ZN(n9213) );
  BUF_X1 U3036 ( .A(n9218), .Z(n9214) );
  INV_X1 U3037 ( .A(n2374), .ZN(n9215) );
  INV_X1 U3038 ( .A(n9215), .ZN(n9216) );
  INV_X1 U3039 ( .A(n5913), .ZN(n9217) );
  INV_X1 U3040 ( .A(n9217), .ZN(n9218) );
  BUF_X1 U3041 ( .A(n9223), .Z(n9219) );
  INV_X1 U3042 ( .A(n2375), .ZN(n9220) );
  INV_X1 U3043 ( .A(n9220), .ZN(n9221) );
  INV_X1 U3044 ( .A(n5914), .ZN(n9222) );
  INV_X1 U3045 ( .A(n9222), .ZN(n9223) );
  BUF_X1 U3046 ( .A(n9228), .Z(n9224) );
  INV_X1 U3047 ( .A(n2376), .ZN(n9225) );
  INV_X1 U3048 ( .A(n9225), .ZN(n9226) );
  INV_X1 U3049 ( .A(n5915), .ZN(n9227) );
  INV_X1 U3050 ( .A(n9227), .ZN(n9228) );
  BUF_X1 U3051 ( .A(n9233), .Z(n9229) );
  INV_X1 U3052 ( .A(n2377), .ZN(n9230) );
  INV_X1 U3053 ( .A(n9230), .ZN(n9231) );
  INV_X1 U3054 ( .A(n5916), .ZN(n9232) );
  INV_X1 U3055 ( .A(n9232), .ZN(n9233) );
  BUF_X1 U3056 ( .A(n9238), .Z(n9234) );
  INV_X1 U3057 ( .A(n2378), .ZN(n9235) );
  INV_X1 U3058 ( .A(n9235), .ZN(n9236) );
  INV_X1 U3059 ( .A(n5917), .ZN(n9237) );
  INV_X1 U3060 ( .A(n9237), .ZN(n9238) );
  BUF_X1 U3061 ( .A(n9243), .Z(n9239) );
  INV_X1 U3062 ( .A(n2379), .ZN(n9240) );
  INV_X1 U3063 ( .A(n9240), .ZN(n9241) );
  INV_X1 U3064 ( .A(n5918), .ZN(n9242) );
  INV_X1 U3065 ( .A(n9242), .ZN(n9243) );
  BUF_X1 U3066 ( .A(n9248), .Z(n9244) );
  INV_X1 U3067 ( .A(n2380), .ZN(n9245) );
  INV_X1 U3068 ( .A(n9245), .ZN(n9246) );
  INV_X1 U3069 ( .A(n5919), .ZN(n9247) );
  INV_X1 U3070 ( .A(n9247), .ZN(n9248) );
  BUF_X1 U3071 ( .A(n9252), .Z(n9249) );
  INV_X1 U3072 ( .A(matrix_mul_2D_4__0__0_), .ZN(n9250) );
  INV_X1 U3073 ( .A(n5920), .ZN(n9251) );
  INV_X1 U3074 ( .A(n9251), .ZN(n9252) );
  BUF_X1 U3075 ( .A(n27528), .Z(n9253) );
  BUF_X1 U3076 ( .A(n27529), .Z(n9254) );
  BUF_X1 U3077 ( .A(n27530), .Z(n9255) );
  BUF_X1 U3078 ( .A(n27531), .Z(n9256) );
  BUF_X1 U3079 ( .A(n27532), .Z(n9257) );
  BUF_X1 U3080 ( .A(n27533), .Z(n9258) );
  BUF_X1 U3081 ( .A(n9263), .Z(n9259) );
  INV_X1 U3082 ( .A(n2352), .ZN(n9260) );
  INV_X1 U3083 ( .A(n9260), .ZN(n9261) );
  INV_X1 U3084 ( .A(n5891), .ZN(n9262) );
  INV_X1 U3085 ( .A(n9262), .ZN(n9263) );
  BUF_X1 U3086 ( .A(n9268), .Z(n9264) );
  INV_X1 U3087 ( .A(n2353), .ZN(n9265) );
  INV_X1 U3088 ( .A(n9265), .ZN(n9266) );
  INV_X1 U3089 ( .A(n58920), .ZN(n9267) );
  INV_X1 U3090 ( .A(n9267), .ZN(n9268) );
  BUF_X1 U3091 ( .A(n9273), .Z(n9269) );
  INV_X1 U3092 ( .A(n2354), .ZN(n9270) );
  INV_X1 U3093 ( .A(n9270), .ZN(n9271) );
  INV_X1 U3094 ( .A(n58930), .ZN(n9272) );
  INV_X1 U3095 ( .A(n9272), .ZN(n9273) );
  BUF_X1 U3096 ( .A(n9278), .Z(n9274) );
  INV_X1 U3097 ( .A(n2355), .ZN(n9275) );
  INV_X1 U3098 ( .A(n9275), .ZN(n9276) );
  INV_X1 U3099 ( .A(n58940), .ZN(n9277) );
  INV_X1 U3100 ( .A(n9277), .ZN(n9278) );
  BUF_X1 U3101 ( .A(n9283), .Z(n9279) );
  INV_X1 U3102 ( .A(n2356), .ZN(n9280) );
  INV_X1 U3103 ( .A(n9280), .ZN(n9281) );
  INV_X1 U3104 ( .A(n58950), .ZN(n9282) );
  INV_X1 U3105 ( .A(n9282), .ZN(n9283) );
  BUF_X1 U3106 ( .A(n9288), .Z(n9284) );
  INV_X1 U3107 ( .A(n2357), .ZN(n9285) );
  INV_X1 U3108 ( .A(n9285), .ZN(n9286) );
  INV_X1 U3109 ( .A(n58960), .ZN(n9287) );
  INV_X1 U3110 ( .A(n9287), .ZN(n9288) );
  BUF_X1 U3111 ( .A(n9293), .Z(n9289) );
  INV_X1 U3112 ( .A(n2358), .ZN(n9290) );
  INV_X1 U3113 ( .A(n9290), .ZN(n9291) );
  INV_X1 U3114 ( .A(n58970), .ZN(n9292) );
  INV_X1 U3115 ( .A(n9292), .ZN(n9293) );
  BUF_X1 U3116 ( .A(n9298), .Z(n9294) );
  INV_X1 U3117 ( .A(n2359), .ZN(n9295) );
  INV_X1 U3118 ( .A(n9295), .ZN(n9296) );
  INV_X1 U3119 ( .A(n58980), .ZN(n9297) );
  INV_X1 U3120 ( .A(n9297), .ZN(n9298) );
  BUF_X1 U3121 ( .A(n9303), .Z(n9299) );
  INV_X1 U3122 ( .A(n2360), .ZN(n9300) );
  INV_X1 U3123 ( .A(n9300), .ZN(n9301) );
  INV_X1 U3124 ( .A(n58990), .ZN(n9302) );
  INV_X1 U3125 ( .A(n9302), .ZN(n9303) );
  BUF_X1 U3126 ( .A(n9308), .Z(n9304) );
  INV_X1 U3127 ( .A(n2361), .ZN(n9305) );
  INV_X1 U3128 ( .A(n9305), .ZN(n9306) );
  INV_X1 U3129 ( .A(n59000), .ZN(n9307) );
  INV_X1 U3130 ( .A(n9307), .ZN(n9308) );
  BUF_X1 U3131 ( .A(n9313), .Z(n9309) );
  INV_X1 U3132 ( .A(n2362), .ZN(n9310) );
  INV_X1 U3133 ( .A(n9310), .ZN(n9311) );
  INV_X1 U3134 ( .A(n59010), .ZN(n9312) );
  INV_X1 U3135 ( .A(n9312), .ZN(n9313) );
  BUF_X1 U3136 ( .A(n9318), .Z(n9314) );
  INV_X1 U3137 ( .A(n2363), .ZN(n9315) );
  INV_X1 U3138 ( .A(n9315), .ZN(n9316) );
  INV_X1 U3139 ( .A(n59020), .ZN(n9317) );
  INV_X1 U3140 ( .A(n9317), .ZN(n9318) );
  BUF_X1 U3141 ( .A(n9323), .Z(n9319) );
  INV_X1 U3142 ( .A(n2364), .ZN(n9320) );
  INV_X1 U3143 ( .A(n9320), .ZN(n9321) );
  INV_X1 U3144 ( .A(n59030), .ZN(n9322) );
  INV_X1 U3145 ( .A(n9322), .ZN(n9323) );
  BUF_X1 U3146 ( .A(n9328), .Z(n9324) );
  INV_X1 U3147 ( .A(n2365), .ZN(n9325) );
  INV_X1 U3148 ( .A(n9325), .ZN(n9326) );
  INV_X1 U3149 ( .A(n59040), .ZN(n9327) );
  INV_X1 U3150 ( .A(n9327), .ZN(n9328) );
  BUF_X1 U3151 ( .A(n9332), .Z(n9329) );
  INV_X1 U3152 ( .A(matrix_mul_2D_3__7__0_), .ZN(n9330) );
  INV_X1 U3153 ( .A(n59050), .ZN(n9331) );
  INV_X1 U3154 ( .A(n9331), .ZN(n9332) );
  BUF_X1 U3155 ( .A(n27522), .Z(n9333) );
  BUF_X1 U3156 ( .A(n27523), .Z(n9334) );
  BUF_X1 U3157 ( .A(n27524), .Z(n9335) );
  BUF_X1 U3158 ( .A(n27525), .Z(n9336) );
  BUF_X1 U3159 ( .A(n27526), .Z(n9337) );
  BUF_X1 U3160 ( .A(n27527), .Z(n9338) );
  BUF_X1 U3161 ( .A(n9343), .Z(n9339) );
  INV_X1 U3162 ( .A(n2337), .ZN(n9340) );
  INV_X1 U3163 ( .A(n9340), .ZN(n9341) );
  INV_X1 U3164 ( .A(n5876), .ZN(n9342) );
  INV_X1 U3165 ( .A(n9342), .ZN(n9343) );
  BUF_X1 U3166 ( .A(n9348), .Z(n9344) );
  INV_X1 U3167 ( .A(n2338), .ZN(n9345) );
  INV_X1 U3168 ( .A(n9345), .ZN(n9346) );
  INV_X1 U3169 ( .A(n5877), .ZN(n9347) );
  INV_X1 U3170 ( .A(n9347), .ZN(n9348) );
  BUF_X1 U3171 ( .A(n9353), .Z(n9349) );
  INV_X1 U3172 ( .A(n2339), .ZN(n9350) );
  INV_X1 U3173 ( .A(n9350), .ZN(n9351) );
  INV_X1 U3174 ( .A(n5878), .ZN(n9352) );
  INV_X1 U3175 ( .A(n9352), .ZN(n9353) );
  BUF_X1 U3176 ( .A(n9358), .Z(n9354) );
  INV_X1 U3177 ( .A(n2340), .ZN(n9355) );
  INV_X1 U3178 ( .A(n9355), .ZN(n9356) );
  INV_X1 U3179 ( .A(n5879), .ZN(n9357) );
  INV_X1 U3180 ( .A(n9357), .ZN(n9358) );
  BUF_X1 U3181 ( .A(n9363), .Z(n9359) );
  INV_X1 U3182 ( .A(n2341), .ZN(n9360) );
  INV_X1 U3183 ( .A(n9360), .ZN(n9361) );
  INV_X1 U3184 ( .A(n5880), .ZN(n9362) );
  INV_X1 U3185 ( .A(n9362), .ZN(n9363) );
  BUF_X1 U3186 ( .A(n9368), .Z(n9364) );
  INV_X1 U3187 ( .A(n2342), .ZN(n9365) );
  INV_X1 U3188 ( .A(n9365), .ZN(n9366) );
  INV_X1 U3189 ( .A(n5881), .ZN(n9367) );
  INV_X1 U3190 ( .A(n9367), .ZN(n9368) );
  BUF_X1 U3191 ( .A(n9373), .Z(n9369) );
  INV_X1 U3192 ( .A(n2343), .ZN(n9370) );
  INV_X1 U3193 ( .A(n9370), .ZN(n9371) );
  INV_X1 U3194 ( .A(n5882), .ZN(n9372) );
  INV_X1 U3195 ( .A(n9372), .ZN(n9373) );
  BUF_X1 U3196 ( .A(n9378), .Z(n9374) );
  INV_X1 U3197 ( .A(n2344), .ZN(n9375) );
  INV_X1 U3198 ( .A(n9375), .ZN(n9376) );
  INV_X1 U3199 ( .A(n5883), .ZN(n9377) );
  INV_X1 U3200 ( .A(n9377), .ZN(n9378) );
  BUF_X1 U3201 ( .A(n9383), .Z(n9379) );
  INV_X1 U3202 ( .A(n2345), .ZN(n9380) );
  INV_X1 U3203 ( .A(n9380), .ZN(n9381) );
  INV_X1 U3204 ( .A(n5884), .ZN(n9382) );
  INV_X1 U3205 ( .A(n9382), .ZN(n9383) );
  BUF_X1 U3206 ( .A(n9388), .Z(n9384) );
  INV_X1 U3207 ( .A(n2346), .ZN(n9385) );
  INV_X1 U3208 ( .A(n9385), .ZN(n9386) );
  INV_X1 U3209 ( .A(n5885), .ZN(n9387) );
  INV_X1 U3210 ( .A(n9387), .ZN(n9388) );
  BUF_X1 U3211 ( .A(n9393), .Z(n9389) );
  INV_X1 U3212 ( .A(n2347), .ZN(n9390) );
  INV_X1 U3213 ( .A(n9390), .ZN(n9391) );
  INV_X1 U3214 ( .A(n5886), .ZN(n9392) );
  INV_X1 U3215 ( .A(n9392), .ZN(n9393) );
  BUF_X1 U3216 ( .A(n9398), .Z(n9394) );
  INV_X1 U3217 ( .A(n2348), .ZN(n9395) );
  INV_X1 U3218 ( .A(n9395), .ZN(n9396) );
  INV_X1 U3219 ( .A(n5887), .ZN(n9397) );
  INV_X1 U3220 ( .A(n9397), .ZN(n9398) );
  BUF_X1 U3221 ( .A(n9403), .Z(n9399) );
  INV_X1 U3222 ( .A(n2349), .ZN(n9400) );
  INV_X1 U3223 ( .A(n9400), .ZN(n9401) );
  INV_X1 U3224 ( .A(n58880), .ZN(n9402) );
  INV_X1 U3225 ( .A(n9402), .ZN(n9403) );
  BUF_X1 U3226 ( .A(n9408), .Z(n9404) );
  INV_X1 U3227 ( .A(n2350), .ZN(n9405) );
  INV_X1 U3228 ( .A(n9405), .ZN(n9406) );
  INV_X1 U3229 ( .A(n5889), .ZN(n9407) );
  INV_X1 U3230 ( .A(n9407), .ZN(n9408) );
  BUF_X1 U3231 ( .A(n9412), .Z(n9409) );
  INV_X1 U3232 ( .A(matrix_mul_2D_3__6__0_), .ZN(n9410) );
  INV_X1 U3233 ( .A(n5890), .ZN(n9411) );
  INV_X1 U3234 ( .A(n9411), .ZN(n9412) );
  BUF_X1 U3235 ( .A(n27516), .Z(n9413) );
  BUF_X1 U3236 ( .A(n27517), .Z(n9414) );
  BUF_X1 U3237 ( .A(n27518), .Z(n9415) );
  BUF_X1 U3238 ( .A(n27519), .Z(n9416) );
  BUF_X1 U3239 ( .A(n27520), .Z(n9417) );
  BUF_X1 U3240 ( .A(n27521), .Z(n9418) );
  BUF_X1 U3241 ( .A(n9423), .Z(n9419) );
  INV_X1 U3242 ( .A(n2322), .ZN(n9420) );
  INV_X1 U3243 ( .A(n9420), .ZN(n9421) );
  INV_X1 U3244 ( .A(n58610), .ZN(n9422) );
  INV_X1 U3245 ( .A(n9422), .ZN(n9423) );
  BUF_X1 U3246 ( .A(n9428), .Z(n9424) );
  INV_X1 U3247 ( .A(n2323), .ZN(n9425) );
  INV_X1 U3248 ( .A(n9425), .ZN(n9426) );
  INV_X1 U3249 ( .A(n58620), .ZN(n9427) );
  INV_X1 U3250 ( .A(n9427), .ZN(n9428) );
  BUF_X1 U3251 ( .A(n9433), .Z(n9429) );
  INV_X1 U3252 ( .A(n2324), .ZN(n9430) );
  INV_X1 U3253 ( .A(n9430), .ZN(n9431) );
  INV_X1 U3254 ( .A(n58630), .ZN(n9432) );
  INV_X1 U3255 ( .A(n9432), .ZN(n9433) );
  BUF_X1 U3256 ( .A(n9438), .Z(n9434) );
  INV_X1 U3257 ( .A(n2325), .ZN(n9435) );
  INV_X1 U3258 ( .A(n9435), .ZN(n9436) );
  INV_X1 U3259 ( .A(n5864), .ZN(n9437) );
  INV_X1 U3260 ( .A(n9437), .ZN(n9438) );
  BUF_X1 U3261 ( .A(n9443), .Z(n9439) );
  INV_X1 U3262 ( .A(n2326), .ZN(n9440) );
  INV_X1 U3263 ( .A(n9440), .ZN(n9441) );
  INV_X1 U3264 ( .A(n5865), .ZN(n9442) );
  INV_X1 U3265 ( .A(n9442), .ZN(n9443) );
  BUF_X1 U3266 ( .A(n9448), .Z(n9444) );
  INV_X1 U3267 ( .A(n2327), .ZN(n9445) );
  INV_X1 U3268 ( .A(n9445), .ZN(n9446) );
  INV_X1 U3269 ( .A(n5866), .ZN(n9447) );
  INV_X1 U3270 ( .A(n9447), .ZN(n9448) );
  BUF_X1 U3271 ( .A(n9453), .Z(n9449) );
  INV_X1 U3272 ( .A(n2328), .ZN(n9450) );
  INV_X1 U3273 ( .A(n9450), .ZN(n9451) );
  INV_X1 U3274 ( .A(n5867), .ZN(n9452) );
  INV_X1 U3275 ( .A(n9452), .ZN(n9453) );
  BUF_X1 U3276 ( .A(n9458), .Z(n9454) );
  INV_X1 U3277 ( .A(n2329), .ZN(n9455) );
  INV_X1 U3278 ( .A(n9455), .ZN(n9456) );
  INV_X1 U3279 ( .A(n5868), .ZN(n9457) );
  INV_X1 U3280 ( .A(n9457), .ZN(n9458) );
  BUF_X1 U3281 ( .A(n9463), .Z(n9459) );
  INV_X1 U3282 ( .A(n2330), .ZN(n9460) );
  INV_X1 U3283 ( .A(n9460), .ZN(n9461) );
  INV_X1 U3284 ( .A(n5869), .ZN(n9462) );
  INV_X1 U3285 ( .A(n9462), .ZN(n9463) );
  BUF_X1 U3286 ( .A(n9468), .Z(n9464) );
  INV_X1 U3287 ( .A(n2331), .ZN(n9465) );
  INV_X1 U3288 ( .A(n9465), .ZN(n9466) );
  INV_X1 U3289 ( .A(n5870), .ZN(n9467) );
  INV_X1 U3290 ( .A(n9467), .ZN(n9468) );
  BUF_X1 U3291 ( .A(n9473), .Z(n9469) );
  INV_X1 U3292 ( .A(n2332), .ZN(n9470) );
  INV_X1 U3293 ( .A(n9470), .ZN(n9471) );
  INV_X1 U3294 ( .A(n5871), .ZN(n9472) );
  INV_X1 U3295 ( .A(n9472), .ZN(n9473) );
  BUF_X1 U3296 ( .A(n9478), .Z(n9474) );
  INV_X1 U3297 ( .A(n2333), .ZN(n9475) );
  INV_X1 U3298 ( .A(n9475), .ZN(n9476) );
  INV_X1 U3299 ( .A(n5872), .ZN(n9477) );
  INV_X1 U3300 ( .A(n9477), .ZN(n9478) );
  BUF_X1 U3301 ( .A(n9483), .Z(n9479) );
  INV_X1 U3302 ( .A(n2334), .ZN(n9480) );
  INV_X1 U3303 ( .A(n9480), .ZN(n9481) );
  INV_X1 U3304 ( .A(n5873), .ZN(n9482) );
  INV_X1 U3305 ( .A(n9482), .ZN(n9483) );
  BUF_X1 U3306 ( .A(n9488), .Z(n9484) );
  INV_X1 U3307 ( .A(n2335), .ZN(n9485) );
  INV_X1 U3308 ( .A(n9485), .ZN(n9486) );
  INV_X1 U3309 ( .A(n5874), .ZN(n9487) );
  INV_X1 U3310 ( .A(n9487), .ZN(n9488) );
  BUF_X1 U3311 ( .A(n9492), .Z(n9489) );
  INV_X1 U3312 ( .A(matrix_mul_2D_3__5__0_), .ZN(n9490) );
  INV_X1 U3313 ( .A(n5875), .ZN(n9491) );
  INV_X1 U3314 ( .A(n9491), .ZN(n9492) );
  BUF_X1 U3315 ( .A(n27510), .Z(n9493) );
  BUF_X1 U3316 ( .A(n27511), .Z(n9494) );
  BUF_X1 U3317 ( .A(n27512), .Z(n9495) );
  BUF_X1 U3318 ( .A(n27513), .Z(n9496) );
  BUF_X1 U3319 ( .A(n27514), .Z(n9497) );
  BUF_X1 U3320 ( .A(n27515), .Z(n9498) );
  BUF_X1 U3321 ( .A(n9502), .Z(n9499) );
  INV_X1 U3322 ( .A(matrix_mul_2D_3__4__14_), .ZN(n9500) );
  INV_X1 U3323 ( .A(n58460), .ZN(n9501) );
  INV_X1 U3324 ( .A(n9501), .ZN(n9502) );
  BUF_X1 U3325 ( .A(n9506), .Z(n9503) );
  INV_X1 U3326 ( .A(matrix_mul_2D_3__4__13_), .ZN(n9504) );
  INV_X1 U3327 ( .A(n58470), .ZN(n9505) );
  INV_X1 U3328 ( .A(n9505), .ZN(n9506) );
  BUF_X1 U3329 ( .A(n9510), .Z(n9507) );
  INV_X1 U3330 ( .A(matrix_mul_2D_3__4__12_), .ZN(n9508) );
  INV_X1 U3331 ( .A(n58480), .ZN(n9509) );
  INV_X1 U3332 ( .A(n9509), .ZN(n9510) );
  BUF_X1 U3333 ( .A(n9514), .Z(n9511) );
  INV_X1 U3334 ( .A(matrix_mul_2D_3__4__11_), .ZN(n9512) );
  INV_X1 U3335 ( .A(n58490), .ZN(n9513) );
  INV_X1 U3336 ( .A(n9513), .ZN(n9514) );
  BUF_X1 U3337 ( .A(n9518), .Z(n9515) );
  INV_X1 U3338 ( .A(matrix_mul_2D_3__4__10_), .ZN(n9516) );
  INV_X1 U3339 ( .A(n58500), .ZN(n9517) );
  INV_X1 U3340 ( .A(n9517), .ZN(n9518) );
  BUF_X1 U3341 ( .A(n9522), .Z(n9519) );
  INV_X1 U3342 ( .A(matrix_mul_2D_3__4__9_), .ZN(n9520) );
  INV_X1 U3343 ( .A(n58510), .ZN(n9521) );
  INV_X1 U3344 ( .A(n9521), .ZN(n9522) );
  BUF_X1 U3345 ( .A(n9526), .Z(n9523) );
  INV_X1 U3346 ( .A(matrix_mul_2D_3__4__8_), .ZN(n9524) );
  INV_X1 U3347 ( .A(n58520), .ZN(n9525) );
  INV_X1 U3348 ( .A(n9525), .ZN(n9526) );
  BUF_X1 U3349 ( .A(n9530), .Z(n9527) );
  INV_X1 U3350 ( .A(matrix_mul_2D_3__4__7_), .ZN(n9528) );
  INV_X1 U3351 ( .A(n58530), .ZN(n9529) );
  INV_X1 U3352 ( .A(n9529), .ZN(n9530) );
  BUF_X1 U3353 ( .A(n9534), .Z(n9531) );
  INV_X1 U3354 ( .A(matrix_mul_2D_3__4__6_), .ZN(n9532) );
  INV_X1 U3355 ( .A(n58540), .ZN(n9533) );
  INV_X1 U3356 ( .A(n9533), .ZN(n9534) );
  BUF_X1 U3357 ( .A(n9538), .Z(n9535) );
  INV_X1 U3358 ( .A(matrix_mul_2D_3__4__5_), .ZN(n9536) );
  INV_X1 U3359 ( .A(n58550), .ZN(n9537) );
  INV_X1 U3360 ( .A(n9537), .ZN(n9538) );
  BUF_X1 U3361 ( .A(n9542), .Z(n9539) );
  INV_X1 U3362 ( .A(matrix_mul_2D_3__4__4_), .ZN(n9540) );
  INV_X1 U3363 ( .A(n58560), .ZN(n9541) );
  INV_X1 U3364 ( .A(n9541), .ZN(n9542) );
  BUF_X1 U3365 ( .A(n9546), .Z(n9543) );
  INV_X1 U3366 ( .A(matrix_mul_2D_3__4__3_), .ZN(n9544) );
  INV_X1 U3367 ( .A(n58570), .ZN(n9545) );
  INV_X1 U3368 ( .A(n9545), .ZN(n9546) );
  BUF_X1 U3369 ( .A(n9550), .Z(n9547) );
  INV_X1 U3370 ( .A(matrix_mul_2D_3__4__2_), .ZN(n9548) );
  INV_X1 U3371 ( .A(n58580), .ZN(n9549) );
  INV_X1 U3372 ( .A(n9549), .ZN(n9550) );
  BUF_X1 U3373 ( .A(n9554), .Z(n9551) );
  INV_X1 U3374 ( .A(matrix_mul_2D_3__4__1_), .ZN(n9552) );
  INV_X1 U3375 ( .A(n58590), .ZN(n9553) );
  INV_X1 U3376 ( .A(n9553), .ZN(n9554) );
  BUF_X1 U3377 ( .A(n9559), .Z(n9555) );
  INV_X1 U3378 ( .A(n2321), .ZN(n9556) );
  INV_X1 U3379 ( .A(n9556), .ZN(n9557) );
  INV_X1 U3380 ( .A(n58600), .ZN(n9558) );
  INV_X1 U3381 ( .A(n9558), .ZN(n9559) );
  BUF_X1 U3382 ( .A(n27504), .Z(n9560) );
  BUF_X1 U3383 ( .A(n27505), .Z(n9561) );
  BUF_X1 U3384 ( .A(n27506), .Z(n9562) );
  BUF_X1 U3385 ( .A(n27507), .Z(n9563) );
  BUF_X1 U3386 ( .A(n27508), .Z(n9564) );
  BUF_X1 U3387 ( .A(n27509), .Z(n9565) );
  BUF_X1 U3388 ( .A(n9569), .Z(n9566) );
  INV_X1 U3389 ( .A(matrix_mul_2D_3__3__14_), .ZN(n9567) );
  INV_X1 U3390 ( .A(n5831), .ZN(n9568) );
  INV_X1 U3391 ( .A(n9568), .ZN(n9569) );
  BUF_X1 U3392 ( .A(n9573), .Z(n9570) );
  INV_X1 U3393 ( .A(matrix_mul_2D_3__3__13_), .ZN(n9571) );
  INV_X1 U3394 ( .A(n5832), .ZN(n9572) );
  INV_X1 U3395 ( .A(n9572), .ZN(n9573) );
  BUF_X1 U3396 ( .A(n9577), .Z(n9574) );
  INV_X1 U3397 ( .A(matrix_mul_2D_3__3__12_), .ZN(n9575) );
  INV_X1 U3398 ( .A(n5833), .ZN(n9576) );
  INV_X1 U3399 ( .A(n9576), .ZN(n9577) );
  BUF_X1 U3400 ( .A(n9581), .Z(n9578) );
  INV_X1 U3401 ( .A(matrix_mul_2D_3__3__11_), .ZN(n9579) );
  INV_X1 U3402 ( .A(n5834), .ZN(n9580) );
  INV_X1 U3403 ( .A(n9580), .ZN(n9581) );
  BUF_X1 U3404 ( .A(n9585), .Z(n9582) );
  INV_X1 U3405 ( .A(matrix_mul_2D_3__3__10_), .ZN(n9583) );
  INV_X1 U3406 ( .A(n5835), .ZN(n9584) );
  INV_X1 U3407 ( .A(n9584), .ZN(n9585) );
  BUF_X1 U3408 ( .A(n9589), .Z(n9586) );
  INV_X1 U3409 ( .A(matrix_mul_2D_3__3__9_), .ZN(n9587) );
  INV_X1 U3410 ( .A(n5836), .ZN(n9588) );
  INV_X1 U3411 ( .A(n9588), .ZN(n9589) );
  BUF_X1 U3412 ( .A(n9593), .Z(n9590) );
  INV_X1 U3413 ( .A(matrix_mul_2D_3__3__8_), .ZN(n9591) );
  INV_X1 U3414 ( .A(n5837), .ZN(n9592) );
  INV_X1 U3415 ( .A(n9592), .ZN(n9593) );
  BUF_X1 U3416 ( .A(n9597), .Z(n9594) );
  INV_X1 U3417 ( .A(matrix_mul_2D_3__3__7_), .ZN(n9595) );
  INV_X1 U3418 ( .A(n5838), .ZN(n9596) );
  INV_X1 U3419 ( .A(n9596), .ZN(n9597) );
  BUF_X1 U3420 ( .A(n9601), .Z(n9598) );
  INV_X1 U3421 ( .A(matrix_mul_2D_3__3__6_), .ZN(n9599) );
  INV_X1 U3422 ( .A(n5839), .ZN(n9600) );
  INV_X1 U3423 ( .A(n9600), .ZN(n9601) );
  BUF_X1 U3424 ( .A(n9605), .Z(n9602) );
  INV_X1 U3425 ( .A(matrix_mul_2D_3__3__5_), .ZN(n9603) );
  INV_X1 U3426 ( .A(n5840), .ZN(n9604) );
  INV_X1 U3427 ( .A(n9604), .ZN(n9605) );
  BUF_X1 U3428 ( .A(n9609), .Z(n9606) );
  INV_X1 U3429 ( .A(matrix_mul_2D_3__3__4_), .ZN(n9607) );
  INV_X1 U3430 ( .A(n5841), .ZN(n9608) );
  INV_X1 U3431 ( .A(n9608), .ZN(n9609) );
  BUF_X1 U3432 ( .A(n9613), .Z(n9610) );
  INV_X1 U3433 ( .A(matrix_mul_2D_3__3__3_), .ZN(n9611) );
  INV_X1 U3434 ( .A(n5842), .ZN(n9612) );
  INV_X1 U3435 ( .A(n9612), .ZN(n9613) );
  BUF_X1 U3436 ( .A(n9617), .Z(n9614) );
  INV_X1 U3437 ( .A(matrix_mul_2D_3__3__2_), .ZN(n9615) );
  INV_X1 U3438 ( .A(n58430), .ZN(n9616) );
  INV_X1 U3439 ( .A(n9616), .ZN(n9617) );
  BUF_X1 U3440 ( .A(n9621), .Z(n9618) );
  INV_X1 U3441 ( .A(matrix_mul_2D_3__3__1_), .ZN(n9619) );
  INV_X1 U3442 ( .A(n58440), .ZN(n9620) );
  INV_X1 U3443 ( .A(n9620), .ZN(n9621) );
  BUF_X1 U3444 ( .A(n9626), .Z(n9622) );
  INV_X1 U3445 ( .A(n2306), .ZN(n9623) );
  INV_X1 U3446 ( .A(n9623), .ZN(n9624) );
  INV_X1 U3447 ( .A(n58450), .ZN(n9625) );
  INV_X1 U3448 ( .A(n9625), .ZN(n9626) );
  BUF_X1 U3449 ( .A(n27498), .Z(n9627) );
  BUF_X1 U3450 ( .A(n27499), .Z(n9628) );
  BUF_X1 U3451 ( .A(n27500), .Z(n9629) );
  BUF_X1 U3452 ( .A(n27501), .Z(n9630) );
  BUF_X1 U3453 ( .A(n27502), .Z(n9631) );
  BUF_X1 U3454 ( .A(n27503), .Z(n9632) );
  BUF_X1 U3455 ( .A(n9637), .Z(n9633) );
  INV_X1 U3456 ( .A(n2271), .ZN(n9634) );
  INV_X1 U3457 ( .A(n9634), .ZN(n9635) );
  INV_X1 U3458 ( .A(n58160), .ZN(n9636) );
  INV_X1 U3459 ( .A(n9636), .ZN(n9637) );
  BUF_X1 U3460 ( .A(n9642), .Z(n9638) );
  INV_X1 U3461 ( .A(n2272), .ZN(n9639) );
  INV_X1 U3462 ( .A(n9639), .ZN(n9640) );
  INV_X1 U3463 ( .A(n58170), .ZN(n9641) );
  INV_X1 U3464 ( .A(n9641), .ZN(n9642) );
  BUF_X1 U3465 ( .A(n9647), .Z(n9643) );
  INV_X1 U3466 ( .A(n2273), .ZN(n9644) );
  INV_X1 U3467 ( .A(n9644), .ZN(n9645) );
  INV_X1 U3468 ( .A(n58180), .ZN(n9646) );
  INV_X1 U3469 ( .A(n9646), .ZN(n9647) );
  BUF_X1 U3470 ( .A(n9652), .Z(n9648) );
  INV_X1 U3471 ( .A(n2274), .ZN(n9649) );
  INV_X1 U3472 ( .A(n9649), .ZN(n9650) );
  INV_X1 U3473 ( .A(n58190), .ZN(n9651) );
  INV_X1 U3474 ( .A(n9651), .ZN(n9652) );
  BUF_X1 U3475 ( .A(n9657), .Z(n9653) );
  INV_X1 U3476 ( .A(n2275), .ZN(n9654) );
  INV_X1 U3477 ( .A(n9654), .ZN(n9655) );
  INV_X1 U3478 ( .A(n58200), .ZN(n9656) );
  INV_X1 U3479 ( .A(n9656), .ZN(n9657) );
  BUF_X1 U3480 ( .A(n9662), .Z(n9658) );
  INV_X1 U3481 ( .A(n2276), .ZN(n9659) );
  INV_X1 U3482 ( .A(n9659), .ZN(n9660) );
  INV_X1 U3483 ( .A(n58210), .ZN(n9661) );
  INV_X1 U3484 ( .A(n9661), .ZN(n9662) );
  BUF_X1 U3485 ( .A(n9667), .Z(n9663) );
  INV_X1 U3486 ( .A(n2277), .ZN(n9664) );
  INV_X1 U3487 ( .A(n9664), .ZN(n9665) );
  INV_X1 U3488 ( .A(n58220), .ZN(n9666) );
  INV_X1 U3489 ( .A(n9666), .ZN(n9667) );
  BUF_X1 U3490 ( .A(n9672), .Z(n9668) );
  INV_X1 U3491 ( .A(n2278), .ZN(n9669) );
  INV_X1 U3492 ( .A(n9669), .ZN(n9670) );
  INV_X1 U3493 ( .A(n58230), .ZN(n9671) );
  INV_X1 U3494 ( .A(n9671), .ZN(n9672) );
  BUF_X1 U3495 ( .A(n9677), .Z(n9673) );
  INV_X1 U3496 ( .A(n2279), .ZN(n9674) );
  INV_X1 U3497 ( .A(n9674), .ZN(n9675) );
  INV_X1 U3498 ( .A(n58240), .ZN(n9676) );
  INV_X1 U3499 ( .A(n9676), .ZN(n9677) );
  BUF_X1 U3500 ( .A(n9682), .Z(n9678) );
  INV_X1 U3501 ( .A(n2280), .ZN(n9679) );
  INV_X1 U3502 ( .A(n9679), .ZN(n9680) );
  INV_X1 U3503 ( .A(n58250), .ZN(n9681) );
  INV_X1 U3504 ( .A(n9681), .ZN(n9682) );
  BUF_X1 U3505 ( .A(n9687), .Z(n9683) );
  INV_X1 U3506 ( .A(n2281), .ZN(n9684) );
  INV_X1 U3507 ( .A(n9684), .ZN(n9685) );
  INV_X1 U3508 ( .A(n5826), .ZN(n9686) );
  INV_X1 U3509 ( .A(n9686), .ZN(n9687) );
  BUF_X1 U3510 ( .A(n9692), .Z(n9688) );
  INV_X1 U3511 ( .A(n2282), .ZN(n9689) );
  INV_X1 U3512 ( .A(n9689), .ZN(n9690) );
  INV_X1 U3513 ( .A(n5827), .ZN(n9691) );
  INV_X1 U3514 ( .A(n9691), .ZN(n9692) );
  BUF_X1 U3515 ( .A(n9697), .Z(n9693) );
  INV_X1 U3516 ( .A(n2283), .ZN(n9694) );
  INV_X1 U3517 ( .A(n9694), .ZN(n9695) );
  INV_X1 U3518 ( .A(n5828), .ZN(n9696) );
  INV_X1 U3519 ( .A(n9696), .ZN(n9697) );
  BUF_X1 U3520 ( .A(n9702), .Z(n9698) );
  INV_X1 U3521 ( .A(n2284), .ZN(n9699) );
  INV_X1 U3522 ( .A(n9699), .ZN(n9700) );
  INV_X1 U3523 ( .A(n5829), .ZN(n9701) );
  INV_X1 U3524 ( .A(n9701), .ZN(n9702) );
  BUF_X1 U3525 ( .A(n9706), .Z(n9703) );
  INV_X1 U3526 ( .A(matrix_mul_2D_3__2__0_), .ZN(n9704) );
  INV_X1 U3527 ( .A(n5830), .ZN(n9705) );
  INV_X1 U3528 ( .A(n9705), .ZN(n9706) );
  BUF_X1 U3529 ( .A(n27492), .Z(n9707) );
  BUF_X1 U3530 ( .A(n27493), .Z(n9708) );
  BUF_X1 U3531 ( .A(n27494), .Z(n9709) );
  BUF_X1 U3532 ( .A(n27495), .Z(n9710) );
  BUF_X1 U3533 ( .A(n27496), .Z(n9711) );
  BUF_X1 U3534 ( .A(n27497), .Z(n9712) );
  BUF_X1 U3535 ( .A(n9717), .Z(n9713) );
  INV_X1 U3536 ( .A(n2256), .ZN(n9714) );
  INV_X1 U3537 ( .A(n9714), .ZN(n9715) );
  INV_X1 U3538 ( .A(n5801), .ZN(n9716) );
  INV_X1 U3539 ( .A(n9716), .ZN(n9717) );
  BUF_X1 U3540 ( .A(n9722), .Z(n9718) );
  INV_X1 U3541 ( .A(n2257), .ZN(n9719) );
  INV_X1 U3542 ( .A(n9719), .ZN(n9720) );
  INV_X1 U3543 ( .A(n5802), .ZN(n9721) );
  INV_X1 U3544 ( .A(n9721), .ZN(n9722) );
  BUF_X1 U3545 ( .A(n9727), .Z(n9723) );
  INV_X1 U3546 ( .A(n2258), .ZN(n9724) );
  INV_X1 U3547 ( .A(n9724), .ZN(n9725) );
  INV_X1 U3548 ( .A(n5803), .ZN(n9726) );
  INV_X1 U3549 ( .A(n9726), .ZN(n9727) );
  BUF_X1 U3550 ( .A(n9732), .Z(n9728) );
  INV_X1 U3551 ( .A(n2259), .ZN(n9729) );
  INV_X1 U3552 ( .A(n9729), .ZN(n9730) );
  INV_X1 U3553 ( .A(n5804), .ZN(n9731) );
  INV_X1 U3554 ( .A(n9731), .ZN(n9732) );
  BUF_X1 U3555 ( .A(n9737), .Z(n9733) );
  INV_X1 U3556 ( .A(n2260), .ZN(n9734) );
  INV_X1 U3557 ( .A(n9734), .ZN(n9735) );
  INV_X1 U3558 ( .A(n5805), .ZN(n9736) );
  INV_X1 U3559 ( .A(n9736), .ZN(n9737) );
  BUF_X1 U3560 ( .A(n9742), .Z(n9738) );
  INV_X1 U3561 ( .A(n2261), .ZN(n9739) );
  INV_X1 U3562 ( .A(n9739), .ZN(n9740) );
  INV_X1 U3563 ( .A(n5806), .ZN(n9741) );
  INV_X1 U3564 ( .A(n9741), .ZN(n9742) );
  BUF_X1 U3565 ( .A(n9747), .Z(n9743) );
  INV_X1 U3566 ( .A(n2262), .ZN(n9744) );
  INV_X1 U3567 ( .A(n9744), .ZN(n9745) );
  INV_X1 U3568 ( .A(n5807), .ZN(n9746) );
  INV_X1 U3569 ( .A(n9746), .ZN(n9747) );
  BUF_X1 U3570 ( .A(n9752), .Z(n9748) );
  INV_X1 U3571 ( .A(n2263), .ZN(n9749) );
  INV_X1 U3572 ( .A(n9749), .ZN(n9750) );
  INV_X1 U3573 ( .A(n5808), .ZN(n9751) );
  INV_X1 U3574 ( .A(n9751), .ZN(n9752) );
  BUF_X1 U3575 ( .A(n9757), .Z(n9753) );
  INV_X1 U3576 ( .A(n2264), .ZN(n9754) );
  INV_X1 U3577 ( .A(n9754), .ZN(n9755) );
  INV_X1 U3578 ( .A(n5809), .ZN(n9756) );
  INV_X1 U3579 ( .A(n9756), .ZN(n9757) );
  BUF_X1 U3580 ( .A(n9762), .Z(n9758) );
  INV_X1 U3581 ( .A(n2265), .ZN(n9759) );
  INV_X1 U3582 ( .A(n9759), .ZN(n9760) );
  INV_X1 U3583 ( .A(n58100), .ZN(n9761) );
  INV_X1 U3584 ( .A(n9761), .ZN(n9762) );
  BUF_X1 U3585 ( .A(n9767), .Z(n9763) );
  INV_X1 U3586 ( .A(n2266), .ZN(n9764) );
  INV_X1 U3587 ( .A(n9764), .ZN(n9765) );
  INV_X1 U3588 ( .A(n58110), .ZN(n9766) );
  INV_X1 U3589 ( .A(n9766), .ZN(n9767) );
  BUF_X1 U3590 ( .A(n9772), .Z(n9768) );
  INV_X1 U3591 ( .A(n2267), .ZN(n9769) );
  INV_X1 U3592 ( .A(n9769), .ZN(n9770) );
  INV_X1 U3593 ( .A(n58120), .ZN(n9771) );
  INV_X1 U3594 ( .A(n9771), .ZN(n9772) );
  BUF_X1 U3595 ( .A(n9777), .Z(n9773) );
  INV_X1 U3596 ( .A(n2268), .ZN(n9774) );
  INV_X1 U3597 ( .A(n9774), .ZN(n9775) );
  INV_X1 U3598 ( .A(n58130), .ZN(n9776) );
  INV_X1 U3599 ( .A(n9776), .ZN(n9777) );
  BUF_X1 U3600 ( .A(n9782), .Z(n9778) );
  INV_X1 U3601 ( .A(n2269), .ZN(n9779) );
  INV_X1 U3602 ( .A(n9779), .ZN(n9780) );
  INV_X1 U3603 ( .A(n58140), .ZN(n9781) );
  INV_X1 U3604 ( .A(n9781), .ZN(n9782) );
  BUF_X1 U3605 ( .A(n9786), .Z(n9783) );
  INV_X1 U3606 ( .A(matrix_mul_2D_3__1__0_), .ZN(n9784) );
  INV_X1 U3607 ( .A(n58150), .ZN(n9785) );
  INV_X1 U3608 ( .A(n9785), .ZN(n9786) );
  BUF_X1 U3609 ( .A(n27486), .Z(n9787) );
  BUF_X1 U3610 ( .A(n27487), .Z(n9788) );
  BUF_X1 U3611 ( .A(n27488), .Z(n9789) );
  BUF_X1 U3612 ( .A(n27489), .Z(n9790) );
  BUF_X1 U3613 ( .A(n27490), .Z(n9791) );
  BUF_X1 U3614 ( .A(n27491), .Z(n9792) );
  BUF_X1 U3615 ( .A(n9797), .Z(n9793) );
  INV_X1 U3616 ( .A(n2241), .ZN(n9794) );
  INV_X1 U3617 ( .A(n9794), .ZN(n9795) );
  INV_X1 U3618 ( .A(n5786), .ZN(n9796) );
  INV_X1 U3619 ( .A(n9796), .ZN(n9797) );
  BUF_X1 U3620 ( .A(n9802), .Z(n9798) );
  INV_X1 U3621 ( .A(n2242), .ZN(n9799) );
  INV_X1 U3622 ( .A(n9799), .ZN(n9800) );
  INV_X1 U3623 ( .A(n5787), .ZN(n9801) );
  INV_X1 U3624 ( .A(n9801), .ZN(n9802) );
  BUF_X1 U3625 ( .A(n9807), .Z(n9803) );
  INV_X1 U3626 ( .A(n2243), .ZN(n9804) );
  INV_X1 U3627 ( .A(n9804), .ZN(n9805) );
  INV_X1 U3628 ( .A(n5788), .ZN(n9806) );
  INV_X1 U3629 ( .A(n9806), .ZN(n9807) );
  BUF_X1 U3630 ( .A(n9812), .Z(n9808) );
  INV_X1 U3631 ( .A(n2244), .ZN(n9809) );
  INV_X1 U3632 ( .A(n9809), .ZN(n9810) );
  INV_X1 U3633 ( .A(n5789), .ZN(n9811) );
  INV_X1 U3634 ( .A(n9811), .ZN(n9812) );
  BUF_X1 U3635 ( .A(n9817), .Z(n9813) );
  INV_X1 U3636 ( .A(n2245), .ZN(n9814) );
  INV_X1 U3637 ( .A(n9814), .ZN(n9815) );
  INV_X1 U3638 ( .A(n5790), .ZN(n9816) );
  INV_X1 U3639 ( .A(n9816), .ZN(n9817) );
  BUF_X1 U3640 ( .A(n9822), .Z(n9818) );
  INV_X1 U3641 ( .A(n2246), .ZN(n9819) );
  INV_X1 U3642 ( .A(n9819), .ZN(n9820) );
  INV_X1 U3643 ( .A(n5791), .ZN(n9821) );
  INV_X1 U3644 ( .A(n9821), .ZN(n9822) );
  BUF_X1 U3645 ( .A(n9827), .Z(n9823) );
  INV_X1 U3646 ( .A(n2247), .ZN(n9824) );
  INV_X1 U3647 ( .A(n9824), .ZN(n9825) );
  INV_X1 U3648 ( .A(n5792), .ZN(n9826) );
  INV_X1 U3649 ( .A(n9826), .ZN(n9827) );
  BUF_X1 U3650 ( .A(n9832), .Z(n9828) );
  INV_X1 U3651 ( .A(n2248), .ZN(n9829) );
  INV_X1 U3652 ( .A(n9829), .ZN(n9830) );
  INV_X1 U3653 ( .A(n5793), .ZN(n9831) );
  INV_X1 U3654 ( .A(n9831), .ZN(n9832) );
  BUF_X1 U3655 ( .A(n9837), .Z(n9833) );
  INV_X1 U3656 ( .A(n2249), .ZN(n9834) );
  INV_X1 U3657 ( .A(n9834), .ZN(n9835) );
  INV_X1 U3658 ( .A(n5794), .ZN(n9836) );
  INV_X1 U3659 ( .A(n9836), .ZN(n9837) );
  BUF_X1 U3660 ( .A(n9842), .Z(n9838) );
  INV_X1 U3661 ( .A(n2250), .ZN(n9839) );
  INV_X1 U3662 ( .A(n9839), .ZN(n9840) );
  INV_X1 U3663 ( .A(n5795), .ZN(n9841) );
  INV_X1 U3664 ( .A(n9841), .ZN(n9842) );
  BUF_X1 U3665 ( .A(n9847), .Z(n9843) );
  INV_X1 U3666 ( .A(n2251), .ZN(n9844) );
  INV_X1 U3667 ( .A(n9844), .ZN(n9845) );
  INV_X1 U3668 ( .A(n5796), .ZN(n9846) );
  INV_X1 U3669 ( .A(n9846), .ZN(n9847) );
  BUF_X1 U3670 ( .A(n9852), .Z(n9848) );
  INV_X1 U3671 ( .A(n2252), .ZN(n9849) );
  INV_X1 U3672 ( .A(n9849), .ZN(n9850) );
  INV_X1 U3673 ( .A(n5797), .ZN(n9851) );
  INV_X1 U3674 ( .A(n9851), .ZN(n9852) );
  BUF_X1 U3675 ( .A(n9857), .Z(n9853) );
  INV_X1 U3676 ( .A(n2253), .ZN(n9854) );
  INV_X1 U3677 ( .A(n9854), .ZN(n9855) );
  INV_X1 U3678 ( .A(n5798), .ZN(n9856) );
  INV_X1 U3679 ( .A(n9856), .ZN(n9857) );
  BUF_X1 U3680 ( .A(n9862), .Z(n9858) );
  INV_X1 U3681 ( .A(n2254), .ZN(n9859) );
  INV_X1 U3682 ( .A(n9859), .ZN(n9860) );
  INV_X1 U3683 ( .A(n5799), .ZN(n9861) );
  INV_X1 U3684 ( .A(n9861), .ZN(n9862) );
  BUF_X1 U3685 ( .A(n9866), .Z(n9863) );
  INV_X1 U3686 ( .A(matrix_mul_2D_3__0__0_), .ZN(n9864) );
  INV_X1 U3687 ( .A(n5800), .ZN(n9865) );
  INV_X1 U3688 ( .A(n9865), .ZN(n9866) );
  BUF_X1 U3689 ( .A(n274801), .Z(n9867) );
  BUF_X1 U3690 ( .A(n27481), .Z(n9868) );
  BUF_X1 U3691 ( .A(n27482), .Z(n9869) );
  BUF_X1 U3692 ( .A(n27483), .Z(n9870) );
  BUF_X1 U3693 ( .A(n27484), .Z(n9871) );
  BUF_X1 U3694 ( .A(n27485), .Z(n9872) );
  BUF_X1 U3695 ( .A(n9876), .Z(n9873) );
  INV_X1 U3696 ( .A(matrix_mul_2D_2__7__14_), .ZN(n9874) );
  INV_X1 U3697 ( .A(n57710), .ZN(n9875) );
  INV_X1 U3698 ( .A(n9875), .ZN(n9876) );
  BUF_X1 U3699 ( .A(n9880), .Z(n9877) );
  INV_X1 U3700 ( .A(matrix_mul_2D_2__7__13_), .ZN(n9878) );
  INV_X1 U3701 ( .A(n57720), .ZN(n9879) );
  INV_X1 U3702 ( .A(n9879), .ZN(n9880) );
  BUF_X1 U3703 ( .A(n9884), .Z(n9881) );
  INV_X1 U3704 ( .A(matrix_mul_2D_2__7__12_), .ZN(n9882) );
  INV_X1 U3705 ( .A(n57730), .ZN(n9883) );
  INV_X1 U3706 ( .A(n9883), .ZN(n9884) );
  BUF_X1 U3707 ( .A(n9888), .Z(n9885) );
  INV_X1 U3708 ( .A(matrix_mul_2D_2__7__11_), .ZN(n9886) );
  INV_X1 U3709 ( .A(n57740), .ZN(n9887) );
  INV_X1 U3710 ( .A(n9887), .ZN(n9888) );
  BUF_X1 U3711 ( .A(n9892), .Z(n9889) );
  INV_X1 U3712 ( .A(matrix_mul_2D_2__7__10_), .ZN(n9890) );
  INV_X1 U3713 ( .A(n5775), .ZN(n9891) );
  INV_X1 U3714 ( .A(n9891), .ZN(n9892) );
  BUF_X1 U3715 ( .A(n9896), .Z(n9893) );
  INV_X1 U3716 ( .A(matrix_mul_2D_2__7__9_), .ZN(n9894) );
  INV_X1 U3717 ( .A(n5776), .ZN(n9895) );
  INV_X1 U3718 ( .A(n9895), .ZN(n9896) );
  BUF_X1 U3719 ( .A(n9900), .Z(n9897) );
  INV_X1 U3720 ( .A(matrix_mul_2D_2__7__8_), .ZN(n9898) );
  INV_X1 U3721 ( .A(n5777), .ZN(n9899) );
  INV_X1 U3722 ( .A(n9899), .ZN(n9900) );
  BUF_X1 U3723 ( .A(n9904), .Z(n9901) );
  INV_X1 U3724 ( .A(matrix_mul_2D_2__7__7_), .ZN(n9902) );
  INV_X1 U3725 ( .A(n5778), .ZN(n9903) );
  INV_X1 U3726 ( .A(n9903), .ZN(n9904) );
  BUF_X1 U3727 ( .A(n9908), .Z(n9905) );
  INV_X1 U3728 ( .A(matrix_mul_2D_2__7__6_), .ZN(n9906) );
  INV_X1 U3729 ( .A(n5779), .ZN(n9907) );
  INV_X1 U3730 ( .A(n9907), .ZN(n9908) );
  BUF_X1 U3731 ( .A(n9912), .Z(n9909) );
  INV_X1 U3732 ( .A(matrix_mul_2D_2__7__5_), .ZN(n9910) );
  INV_X1 U3733 ( .A(n5780), .ZN(n9911) );
  INV_X1 U3734 ( .A(n9911), .ZN(n9912) );
  BUF_X1 U3735 ( .A(n9916), .Z(n9913) );
  INV_X1 U3736 ( .A(matrix_mul_2D_2__7__4_), .ZN(n9914) );
  INV_X1 U3737 ( .A(n5781), .ZN(n9915) );
  INV_X1 U3738 ( .A(n9915), .ZN(n9916) );
  BUF_X1 U3739 ( .A(n9920), .Z(n9917) );
  INV_X1 U3740 ( .A(matrix_mul_2D_2__7__3_), .ZN(n9918) );
  INV_X1 U3741 ( .A(n5782), .ZN(n9919) );
  INV_X1 U3742 ( .A(n9919), .ZN(n9920) );
  BUF_X1 U3743 ( .A(n9924), .Z(n9921) );
  INV_X1 U3744 ( .A(matrix_mul_2D_2__7__2_), .ZN(n9922) );
  INV_X1 U3745 ( .A(n5783), .ZN(n9923) );
  INV_X1 U3746 ( .A(n9923), .ZN(n9924) );
  BUF_X1 U3747 ( .A(n9928), .Z(n9925) );
  INV_X1 U3748 ( .A(matrix_mul_2D_2__7__1_), .ZN(n9926) );
  INV_X1 U3749 ( .A(n5784), .ZN(n9927) );
  INV_X1 U3750 ( .A(n9927), .ZN(n9928) );
  BUF_X1 U3751 ( .A(n9933), .Z(n9929) );
  INV_X1 U3752 ( .A(n2240), .ZN(n9930) );
  INV_X1 U3753 ( .A(n9930), .ZN(n9931) );
  INV_X1 U3754 ( .A(n5785), .ZN(n9932) );
  INV_X1 U3755 ( .A(n9932), .ZN(n9933) );
  BUF_X1 U3756 ( .A(n27474), .Z(n9934) );
  BUF_X1 U3757 ( .A(n27475), .Z(n9935) );
  BUF_X1 U3758 ( .A(n27476), .Z(n9936) );
  BUF_X1 U3759 ( .A(n27477), .Z(n9937) );
  BUF_X1 U3760 ( .A(n27478), .Z(n9938) );
  BUF_X1 U3761 ( .A(n27479), .Z(n9939) );
  BUF_X1 U3762 ( .A(n9943), .Z(n9940) );
  INV_X1 U3763 ( .A(matrix_mul_2D_2__6__14_), .ZN(n9941) );
  INV_X1 U3764 ( .A(n57560), .ZN(n9942) );
  INV_X1 U3765 ( .A(n9942), .ZN(n9943) );
  BUF_X1 U3766 ( .A(n9947), .Z(n9944) );
  INV_X1 U3767 ( .A(matrix_mul_2D_2__6__13_), .ZN(n9945) );
  INV_X1 U3768 ( .A(n57570), .ZN(n9946) );
  INV_X1 U3769 ( .A(n9946), .ZN(n9947) );
  BUF_X1 U3770 ( .A(n9951), .Z(n9948) );
  INV_X1 U3771 ( .A(matrix_mul_2D_2__6__12_), .ZN(n9949) );
  INV_X1 U3772 ( .A(n57580), .ZN(n9950) );
  INV_X1 U3773 ( .A(n9950), .ZN(n9951) );
  BUF_X1 U3774 ( .A(n9955), .Z(n9952) );
  INV_X1 U3775 ( .A(matrix_mul_2D_2__6__11_), .ZN(n9953) );
  INV_X1 U3776 ( .A(n57590), .ZN(n9954) );
  INV_X1 U3777 ( .A(n9954), .ZN(n9955) );
  BUF_X1 U3778 ( .A(n9959), .Z(n9956) );
  INV_X1 U3779 ( .A(matrix_mul_2D_2__6__10_), .ZN(n9957) );
  INV_X1 U3780 ( .A(n57600), .ZN(n9958) );
  INV_X1 U3781 ( .A(n9958), .ZN(n9959) );
  BUF_X1 U3782 ( .A(n9963), .Z(n9960) );
  INV_X1 U3783 ( .A(matrix_mul_2D_2__6__9_), .ZN(n9961) );
  INV_X1 U3784 ( .A(n57610), .ZN(n9962) );
  INV_X1 U3785 ( .A(n9962), .ZN(n9963) );
  BUF_X1 U3786 ( .A(n9967), .Z(n9964) );
  INV_X1 U3787 ( .A(matrix_mul_2D_2__6__8_), .ZN(n9965) );
  INV_X1 U3788 ( .A(n57620), .ZN(n9966) );
  INV_X1 U3789 ( .A(n9966), .ZN(n9967) );
  BUF_X1 U3790 ( .A(n9971), .Z(n9968) );
  INV_X1 U3791 ( .A(matrix_mul_2D_2__6__7_), .ZN(n9969) );
  INV_X1 U3792 ( .A(n57630), .ZN(n9970) );
  INV_X1 U3793 ( .A(n9970), .ZN(n9971) );
  BUF_X1 U3794 ( .A(n9975), .Z(n9972) );
  INV_X1 U3795 ( .A(matrix_mul_2D_2__6__6_), .ZN(n9973) );
  INV_X1 U3796 ( .A(n57640), .ZN(n9974) );
  INV_X1 U3797 ( .A(n9974), .ZN(n9975) );
  BUF_X1 U3798 ( .A(n9979), .Z(n9976) );
  INV_X1 U3799 ( .A(matrix_mul_2D_2__6__5_), .ZN(n9977) );
  INV_X1 U3800 ( .A(n57650), .ZN(n9978) );
  INV_X1 U3801 ( .A(n9978), .ZN(n9979) );
  BUF_X1 U3802 ( .A(n9983), .Z(n9980) );
  INV_X1 U3803 ( .A(matrix_mul_2D_2__6__4_), .ZN(n9981) );
  INV_X1 U3804 ( .A(n57660), .ZN(n9982) );
  INV_X1 U3805 ( .A(n9982), .ZN(n9983) );
  BUF_X1 U3806 ( .A(n9987), .Z(n9984) );
  INV_X1 U3807 ( .A(matrix_mul_2D_2__6__3_), .ZN(n9985) );
  INV_X1 U3808 ( .A(n57670), .ZN(n9986) );
  INV_X1 U3809 ( .A(n9986), .ZN(n9987) );
  BUF_X1 U3810 ( .A(n9991), .Z(n9988) );
  INV_X1 U3811 ( .A(matrix_mul_2D_2__6__2_), .ZN(n9989) );
  INV_X1 U3812 ( .A(n57680), .ZN(n9990) );
  INV_X1 U3813 ( .A(n9990), .ZN(n9991) );
  BUF_X1 U3814 ( .A(n9995), .Z(n9992) );
  INV_X1 U3815 ( .A(matrix_mul_2D_2__6__1_), .ZN(n9993) );
  INV_X1 U3816 ( .A(n57690), .ZN(n9994) );
  INV_X1 U3817 ( .A(n9994), .ZN(n9995) );
  BUF_X1 U3818 ( .A(n10000), .Z(n9996) );
  INV_X1 U3819 ( .A(n2225), .ZN(n9997) );
  INV_X1 U3820 ( .A(n9997), .ZN(n9998) );
  INV_X1 U3821 ( .A(n57700), .ZN(n9999) );
  INV_X1 U3822 ( .A(n9999), .ZN(n10000) );
  BUF_X1 U3823 ( .A(n27468), .Z(n10001) );
  BUF_X1 U3824 ( .A(n27469), .Z(n10002) );
  BUF_X1 U3825 ( .A(n274701), .Z(n10003) );
  BUF_X1 U3826 ( .A(n27471), .Z(n10004) );
  BUF_X1 U3827 ( .A(n27472), .Z(n10005) );
  BUF_X1 U3828 ( .A(n27473), .Z(n10006) );
  BUF_X1 U3829 ( .A(n10011), .Z(n10007) );
  INV_X1 U3830 ( .A(n2190), .ZN(n10008) );
  INV_X1 U3831 ( .A(n10008), .ZN(n10009) );
  INV_X1 U3832 ( .A(n5741), .ZN(n10010) );
  INV_X1 U3833 ( .A(n10010), .ZN(n10011) );
  BUF_X1 U3834 ( .A(n10016), .Z(n10012) );
  INV_X1 U3835 ( .A(n2191), .ZN(n10013) );
  INV_X1 U3836 ( .A(n10013), .ZN(n10014) );
  INV_X1 U3837 ( .A(n5742), .ZN(n10015) );
  INV_X1 U3838 ( .A(n10015), .ZN(n10016) );
  BUF_X1 U3839 ( .A(n10021), .Z(n10017) );
  INV_X1 U3840 ( .A(n2192), .ZN(n10018) );
  INV_X1 U3841 ( .A(n10018), .ZN(n10019) );
  INV_X1 U3842 ( .A(n5743), .ZN(n10020) );
  INV_X1 U3843 ( .A(n10020), .ZN(n10021) );
  BUF_X1 U3844 ( .A(n10026), .Z(n10022) );
  INV_X1 U3845 ( .A(n2193), .ZN(n10023) );
  INV_X1 U3846 ( .A(n10023), .ZN(n10024) );
  INV_X1 U3847 ( .A(n5744), .ZN(n10025) );
  INV_X1 U3848 ( .A(n10025), .ZN(n10026) );
  BUF_X1 U3849 ( .A(n10031), .Z(n10027) );
  INV_X1 U3850 ( .A(n2194), .ZN(n10028) );
  INV_X1 U3851 ( .A(n10028), .ZN(n10029) );
  INV_X1 U3852 ( .A(n5745), .ZN(n10030) );
  INV_X1 U3853 ( .A(n10030), .ZN(n10031) );
  BUF_X1 U3854 ( .A(n10036), .Z(n10032) );
  INV_X1 U3855 ( .A(n2195), .ZN(n10033) );
  INV_X1 U3856 ( .A(n10033), .ZN(n10034) );
  INV_X1 U3857 ( .A(n5746), .ZN(n10035) );
  INV_X1 U3858 ( .A(n10035), .ZN(n10036) );
  BUF_X1 U3859 ( .A(n10041), .Z(n10037) );
  INV_X1 U3860 ( .A(n2196), .ZN(n10038) );
  INV_X1 U3861 ( .A(n10038), .ZN(n10039) );
  INV_X1 U3862 ( .A(n5747), .ZN(n10040) );
  INV_X1 U3863 ( .A(n10040), .ZN(n10041) );
  BUF_X1 U3864 ( .A(n10046), .Z(n10042) );
  INV_X1 U3865 ( .A(n2197), .ZN(n10043) );
  INV_X1 U3866 ( .A(n10043), .ZN(n10044) );
  INV_X1 U3867 ( .A(n5748), .ZN(n10045) );
  INV_X1 U3868 ( .A(n10045), .ZN(n10046) );
  BUF_X1 U3869 ( .A(n10051), .Z(n10047) );
  INV_X1 U3870 ( .A(n2198), .ZN(n10048) );
  INV_X1 U3871 ( .A(n10048), .ZN(n10049) );
  INV_X1 U3872 ( .A(n5749), .ZN(n10050) );
  INV_X1 U3873 ( .A(n10050), .ZN(n10051) );
  BUF_X1 U3874 ( .A(n10056), .Z(n10052) );
  INV_X1 U3875 ( .A(n2199), .ZN(n10053) );
  INV_X1 U3876 ( .A(n10053), .ZN(n10054) );
  INV_X1 U3877 ( .A(n5750), .ZN(n10055) );
  INV_X1 U3878 ( .A(n10055), .ZN(n10056) );
  BUF_X1 U3879 ( .A(n10061), .Z(n10057) );
  INV_X1 U3880 ( .A(n2200), .ZN(n10058) );
  INV_X1 U3881 ( .A(n10058), .ZN(n10059) );
  INV_X1 U3882 ( .A(n5751), .ZN(n10060) );
  INV_X1 U3883 ( .A(n10060), .ZN(n10061) );
  BUF_X1 U3884 ( .A(n10066), .Z(n10062) );
  INV_X1 U3885 ( .A(n2201), .ZN(n10063) );
  INV_X1 U3886 ( .A(n10063), .ZN(n10064) );
  INV_X1 U3887 ( .A(n5752), .ZN(n10065) );
  INV_X1 U3888 ( .A(n10065), .ZN(n10066) );
  BUF_X1 U3889 ( .A(n10071), .Z(n10067) );
  INV_X1 U3890 ( .A(n2202), .ZN(n10068) );
  INV_X1 U3891 ( .A(n10068), .ZN(n10069) );
  INV_X1 U3892 ( .A(n5753), .ZN(n10070) );
  INV_X1 U3893 ( .A(n10070), .ZN(n10071) );
  BUF_X1 U3894 ( .A(n10076), .Z(n10072) );
  INV_X1 U3895 ( .A(n2203), .ZN(n10073) );
  INV_X1 U3896 ( .A(n10073), .ZN(n10074) );
  INV_X1 U3897 ( .A(n57540), .ZN(n10075) );
  INV_X1 U3898 ( .A(n10075), .ZN(n10076) );
  BUF_X1 U3899 ( .A(n10080), .Z(n10077) );
  INV_X1 U3900 ( .A(matrix_mul_2D_2__5__0_), .ZN(n10078) );
  INV_X1 U3901 ( .A(n57550), .ZN(n10079) );
  INV_X1 U3902 ( .A(n10079), .ZN(n10080) );
  BUF_X1 U3903 ( .A(n27462), .Z(n10081) );
  BUF_X1 U3904 ( .A(n27463), .Z(n10082) );
  BUF_X1 U3905 ( .A(n27464), .Z(n10083) );
  BUF_X1 U3906 ( .A(n27465), .Z(n10084) );
  BUF_X1 U3907 ( .A(n27466), .Z(n10085) );
  BUF_X1 U3908 ( .A(n27467), .Z(n10086) );
  BUF_X1 U3909 ( .A(n10091), .Z(n10087) );
  INV_X1 U3910 ( .A(n2175), .ZN(n10088) );
  INV_X1 U3911 ( .A(n10088), .ZN(n10089) );
  INV_X1 U3912 ( .A(n57260), .ZN(n10090) );
  INV_X1 U3913 ( .A(n10090), .ZN(n10091) );
  BUF_X1 U3914 ( .A(n10096), .Z(n10092) );
  INV_X1 U3915 ( .A(n2176), .ZN(n10093) );
  INV_X1 U3916 ( .A(n10093), .ZN(n10094) );
  INV_X1 U3917 ( .A(n57270), .ZN(n10095) );
  INV_X1 U3918 ( .A(n10095), .ZN(n10096) );
  BUF_X1 U3919 ( .A(n10101), .Z(n10097) );
  INV_X1 U3920 ( .A(n2177), .ZN(n10098) );
  INV_X1 U3921 ( .A(n10098), .ZN(n10099) );
  INV_X1 U3922 ( .A(n57280), .ZN(n10100) );
  INV_X1 U3923 ( .A(n10100), .ZN(n10101) );
  BUF_X1 U3924 ( .A(n10106), .Z(n10102) );
  INV_X1 U3925 ( .A(n2178), .ZN(n10103) );
  INV_X1 U3926 ( .A(n10103), .ZN(n10104) );
  INV_X1 U3927 ( .A(n57290), .ZN(n10105) );
  INV_X1 U3928 ( .A(n10105), .ZN(n10106) );
  BUF_X1 U3929 ( .A(n10111), .Z(n10107) );
  INV_X1 U3930 ( .A(n2179), .ZN(n10108) );
  INV_X1 U3931 ( .A(n10108), .ZN(n10109) );
  INV_X1 U3932 ( .A(n57300), .ZN(n10110) );
  INV_X1 U3933 ( .A(n10110), .ZN(n10111) );
  BUF_X1 U3934 ( .A(n10116), .Z(n10112) );
  INV_X1 U3935 ( .A(n2180), .ZN(n10113) );
  INV_X1 U3936 ( .A(n10113), .ZN(n10114) );
  INV_X1 U3937 ( .A(n57310), .ZN(n10115) );
  INV_X1 U3938 ( .A(n10115), .ZN(n10116) );
  BUF_X1 U3939 ( .A(n10121), .Z(n10117) );
  INV_X1 U3940 ( .A(n2181), .ZN(n10118) );
  INV_X1 U3941 ( .A(n10118), .ZN(n10119) );
  INV_X1 U3942 ( .A(n57320), .ZN(n10120) );
  INV_X1 U3943 ( .A(n10120), .ZN(n10121) );
  BUF_X1 U3944 ( .A(n10126), .Z(n10122) );
  INV_X1 U3945 ( .A(n2182), .ZN(n10123) );
  INV_X1 U3946 ( .A(n10123), .ZN(n10124) );
  INV_X1 U3947 ( .A(n57330), .ZN(n10125) );
  INV_X1 U3948 ( .A(n10125), .ZN(n10126) );
  BUF_X1 U3949 ( .A(n10131), .Z(n10127) );
  INV_X1 U3950 ( .A(n2183), .ZN(n10128) );
  INV_X1 U3951 ( .A(n10128), .ZN(n10129) );
  INV_X1 U3952 ( .A(n57340), .ZN(n10130) );
  INV_X1 U3953 ( .A(n10130), .ZN(n10131) );
  BUF_X1 U3954 ( .A(n10136), .Z(n10132) );
  INV_X1 U3955 ( .A(n2184), .ZN(n10133) );
  INV_X1 U3956 ( .A(n10133), .ZN(n10134) );
  INV_X1 U3957 ( .A(n57350), .ZN(n10135) );
  INV_X1 U3958 ( .A(n10135), .ZN(n10136) );
  BUF_X1 U3959 ( .A(n10141), .Z(n10137) );
  INV_X1 U3960 ( .A(n2185), .ZN(n10138) );
  INV_X1 U3961 ( .A(n10138), .ZN(n10139) );
  INV_X1 U3962 ( .A(n57360), .ZN(n10140) );
  INV_X1 U3963 ( .A(n10140), .ZN(n10141) );
  BUF_X1 U3964 ( .A(n10146), .Z(n10142) );
  INV_X1 U3965 ( .A(n2186), .ZN(n10143) );
  INV_X1 U3966 ( .A(n10143), .ZN(n10144) );
  INV_X1 U3967 ( .A(n5737), .ZN(n10145) );
  INV_X1 U3968 ( .A(n10145), .ZN(n10146) );
  BUF_X1 U3969 ( .A(n10151), .Z(n10147) );
  INV_X1 U3970 ( .A(n2187), .ZN(n10148) );
  INV_X1 U3971 ( .A(n10148), .ZN(n10149) );
  INV_X1 U3972 ( .A(n5738), .ZN(n10150) );
  INV_X1 U3973 ( .A(n10150), .ZN(n10151) );
  BUF_X1 U3974 ( .A(n10156), .Z(n10152) );
  INV_X1 U3975 ( .A(n2188), .ZN(n10153) );
  INV_X1 U3976 ( .A(n10153), .ZN(n10154) );
  INV_X1 U3977 ( .A(n5739), .ZN(n10155) );
  INV_X1 U3978 ( .A(n10155), .ZN(n10156) );
  BUF_X1 U3979 ( .A(n10160), .Z(n10157) );
  INV_X1 U3980 ( .A(matrix_mul_2D_2__4__0_), .ZN(n10158) );
  INV_X1 U3981 ( .A(n5740), .ZN(n10159) );
  INV_X1 U3982 ( .A(n10159), .ZN(n10160) );
  BUF_X1 U3983 ( .A(n27456), .Z(n10161) );
  BUF_X1 U3984 ( .A(n27457), .Z(n10162) );
  BUF_X1 U3985 ( .A(n27458), .Z(n10163) );
  BUF_X1 U3986 ( .A(n27459), .Z(n10164) );
  BUF_X1 U3987 ( .A(n274601), .Z(n10165) );
  BUF_X1 U3988 ( .A(n27461), .Z(n10166) );
  BUF_X1 U3989 ( .A(n10171), .Z(n10167) );
  INV_X1 U3990 ( .A(n2160), .ZN(n10168) );
  INV_X1 U3991 ( .A(n10168), .ZN(n10169) );
  INV_X1 U3992 ( .A(n5711), .ZN(n10170) );
  INV_X1 U3993 ( .A(n10170), .ZN(n10171) );
  BUF_X1 U3994 ( .A(n10176), .Z(n10172) );
  INV_X1 U3995 ( .A(n2161), .ZN(n10173) );
  INV_X1 U3996 ( .A(n10173), .ZN(n10174) );
  INV_X1 U3997 ( .A(n5712), .ZN(n10175) );
  INV_X1 U3998 ( .A(n10175), .ZN(n10176) );
  BUF_X1 U3999 ( .A(n10181), .Z(n10177) );
  INV_X1 U4000 ( .A(n2162), .ZN(n10178) );
  INV_X1 U4001 ( .A(n10178), .ZN(n10179) );
  INV_X1 U4002 ( .A(n5713), .ZN(n10180) );
  INV_X1 U4003 ( .A(n10180), .ZN(n10181) );
  BUF_X1 U4004 ( .A(n10186), .Z(n10182) );
  INV_X1 U4005 ( .A(n2163), .ZN(n10183) );
  INV_X1 U4006 ( .A(n10183), .ZN(n10184) );
  INV_X1 U4007 ( .A(n5714), .ZN(n10185) );
  INV_X1 U4008 ( .A(n10185), .ZN(n10186) );
  BUF_X1 U4009 ( .A(n10191), .Z(n10187) );
  INV_X1 U4010 ( .A(n2164), .ZN(n10188) );
  INV_X1 U4011 ( .A(n10188), .ZN(n10189) );
  INV_X1 U4012 ( .A(n5715), .ZN(n10190) );
  INV_X1 U4013 ( .A(n10190), .ZN(n10191) );
  BUF_X1 U4014 ( .A(n10196), .Z(n10192) );
  INV_X1 U4015 ( .A(n2165), .ZN(n10193) );
  INV_X1 U4016 ( .A(n10193), .ZN(n10194) );
  INV_X1 U4017 ( .A(n5716), .ZN(n10195) );
  INV_X1 U4018 ( .A(n10195), .ZN(n10196) );
  BUF_X1 U4019 ( .A(n10201), .Z(n10197) );
  INV_X1 U4020 ( .A(n2166), .ZN(n10198) );
  INV_X1 U4021 ( .A(n10198), .ZN(n10199) );
  INV_X1 U4022 ( .A(n5717), .ZN(n10200) );
  INV_X1 U4023 ( .A(n10200), .ZN(n10201) );
  BUF_X1 U4024 ( .A(n10206), .Z(n10202) );
  INV_X1 U4025 ( .A(n2167), .ZN(n10203) );
  INV_X1 U4026 ( .A(n10203), .ZN(n10204) );
  INV_X1 U4027 ( .A(n5718), .ZN(n10205) );
  INV_X1 U4028 ( .A(n10205), .ZN(n10206) );
  BUF_X1 U4029 ( .A(n10211), .Z(n10207) );
  INV_X1 U4030 ( .A(n2168), .ZN(n10208) );
  INV_X1 U4031 ( .A(n10208), .ZN(n10209) );
  INV_X1 U4032 ( .A(n5719), .ZN(n10210) );
  INV_X1 U4033 ( .A(n10210), .ZN(n10211) );
  BUF_X1 U4034 ( .A(n10216), .Z(n10212) );
  INV_X1 U4035 ( .A(n2169), .ZN(n10213) );
  INV_X1 U4036 ( .A(n10213), .ZN(n10214) );
  INV_X1 U4037 ( .A(n5720), .ZN(n10215) );
  INV_X1 U4038 ( .A(n10215), .ZN(n10216) );
  BUF_X1 U4039 ( .A(n10221), .Z(n10217) );
  INV_X1 U4040 ( .A(n2170), .ZN(n10218) );
  INV_X1 U4041 ( .A(n10218), .ZN(n10219) );
  INV_X1 U4042 ( .A(n57210), .ZN(n10220) );
  INV_X1 U4043 ( .A(n10220), .ZN(n10221) );
  BUF_X1 U4044 ( .A(n10226), .Z(n10222) );
  INV_X1 U4045 ( .A(n2171), .ZN(n10223) );
  INV_X1 U4046 ( .A(n10223), .ZN(n10224) );
  INV_X1 U4047 ( .A(n57220), .ZN(n10225) );
  INV_X1 U4048 ( .A(n10225), .ZN(n10226) );
  BUF_X1 U4049 ( .A(n10231), .Z(n10227) );
  INV_X1 U4050 ( .A(n2172), .ZN(n10228) );
  INV_X1 U4051 ( .A(n10228), .ZN(n10229) );
  INV_X1 U4052 ( .A(n57230), .ZN(n10230) );
  INV_X1 U4053 ( .A(n10230), .ZN(n10231) );
  BUF_X1 U4054 ( .A(n10236), .Z(n10232) );
  INV_X1 U4055 ( .A(n2173), .ZN(n10233) );
  INV_X1 U4056 ( .A(n10233), .ZN(n10234) );
  INV_X1 U4057 ( .A(n57240), .ZN(n10235) );
  INV_X1 U4058 ( .A(n10235), .ZN(n10236) );
  BUF_X1 U4059 ( .A(n10240), .Z(n10237) );
  INV_X1 U4060 ( .A(matrix_mul_2D_2__3__0_), .ZN(n10238) );
  INV_X1 U4061 ( .A(n57250), .ZN(n10239) );
  INV_X1 U4062 ( .A(n10239), .ZN(n10240) );
  BUF_X1 U4063 ( .A(n274501), .Z(n10241) );
  BUF_X1 U4064 ( .A(n27451), .Z(n10242) );
  BUF_X1 U4065 ( .A(n27452), .Z(n10243) );
  BUF_X1 U4066 ( .A(n27453), .Z(n10244) );
  BUF_X1 U4067 ( .A(n27454), .Z(n10245) );
  BUF_X1 U4068 ( .A(n27455), .Z(n10246) );
  BUF_X1 U4069 ( .A(n10251), .Z(n10247) );
  INV_X1 U4070 ( .A(n2145), .ZN(n10248) );
  INV_X1 U4071 ( .A(n10248), .ZN(n10249) );
  INV_X1 U4072 ( .A(n5696), .ZN(n10250) );
  INV_X1 U4073 ( .A(n10250), .ZN(n10251) );
  BUF_X1 U4074 ( .A(n10256), .Z(n10252) );
  INV_X1 U4075 ( .A(n2146), .ZN(n10253) );
  INV_X1 U4076 ( .A(n10253), .ZN(n10254) );
  INV_X1 U4077 ( .A(n5697), .ZN(n10255) );
  INV_X1 U4078 ( .A(n10255), .ZN(n10256) );
  BUF_X1 U4079 ( .A(n10261), .Z(n10257) );
  INV_X1 U4080 ( .A(n2147), .ZN(n10258) );
  INV_X1 U4081 ( .A(n10258), .ZN(n10259) );
  INV_X1 U4082 ( .A(n5698), .ZN(n10260) );
  INV_X1 U4083 ( .A(n10260), .ZN(n10261) );
  BUF_X1 U4084 ( .A(n10266), .Z(n10262) );
  INV_X1 U4085 ( .A(n2148), .ZN(n10263) );
  INV_X1 U4086 ( .A(n10263), .ZN(n10264) );
  INV_X1 U4087 ( .A(n5699), .ZN(n10265) );
  INV_X1 U4088 ( .A(n10265), .ZN(n10266) );
  BUF_X1 U4089 ( .A(n10271), .Z(n10267) );
  INV_X1 U4090 ( .A(n2149), .ZN(n10268) );
  INV_X1 U4091 ( .A(n10268), .ZN(n10269) );
  INV_X1 U4092 ( .A(n5700), .ZN(n10270) );
  INV_X1 U4093 ( .A(n10270), .ZN(n10271) );
  BUF_X1 U4094 ( .A(n10276), .Z(n10272) );
  INV_X1 U4095 ( .A(n2150), .ZN(n10273) );
  INV_X1 U4096 ( .A(n10273), .ZN(n10274) );
  INV_X1 U4097 ( .A(n5701), .ZN(n10275) );
  INV_X1 U4098 ( .A(n10275), .ZN(n10276) );
  BUF_X1 U4099 ( .A(n10281), .Z(n10277) );
  INV_X1 U4100 ( .A(n2151), .ZN(n10278) );
  INV_X1 U4101 ( .A(n10278), .ZN(n10279) );
  INV_X1 U4102 ( .A(n5702), .ZN(n10280) );
  INV_X1 U4103 ( .A(n10280), .ZN(n10281) );
  BUF_X1 U4104 ( .A(n10286), .Z(n10282) );
  INV_X1 U4105 ( .A(n2152), .ZN(n10283) );
  INV_X1 U4106 ( .A(n10283), .ZN(n10284) );
  INV_X1 U4107 ( .A(n5703), .ZN(n10285) );
  INV_X1 U4108 ( .A(n10285), .ZN(n10286) );
  BUF_X1 U4109 ( .A(n10291), .Z(n10287) );
  INV_X1 U4110 ( .A(n2153), .ZN(n10288) );
  INV_X1 U4111 ( .A(n10288), .ZN(n10289) );
  INV_X1 U4112 ( .A(n5704), .ZN(n10290) );
  INV_X1 U4113 ( .A(n10290), .ZN(n10291) );
  BUF_X1 U4114 ( .A(n10296), .Z(n10292) );
  INV_X1 U4115 ( .A(n2154), .ZN(n10293) );
  INV_X1 U4116 ( .A(n10293), .ZN(n10294) );
  INV_X1 U4117 ( .A(n5705), .ZN(n10295) );
  INV_X1 U4118 ( .A(n10295), .ZN(n10296) );
  BUF_X1 U4119 ( .A(n10301), .Z(n10297) );
  INV_X1 U4120 ( .A(n2155), .ZN(n10298) );
  INV_X1 U4121 ( .A(n10298), .ZN(n10299) );
  INV_X1 U4122 ( .A(n5706), .ZN(n10300) );
  INV_X1 U4123 ( .A(n10300), .ZN(n10301) );
  BUF_X1 U4124 ( .A(n10306), .Z(n10302) );
  INV_X1 U4125 ( .A(n2156), .ZN(n10303) );
  INV_X1 U4126 ( .A(n10303), .ZN(n10304) );
  INV_X1 U4127 ( .A(n5707), .ZN(n10305) );
  INV_X1 U4128 ( .A(n10305), .ZN(n10306) );
  BUF_X1 U4129 ( .A(n10311), .Z(n10307) );
  INV_X1 U4130 ( .A(n2157), .ZN(n10308) );
  INV_X1 U4131 ( .A(n10308), .ZN(n10309) );
  INV_X1 U4132 ( .A(n5708), .ZN(n10310) );
  INV_X1 U4133 ( .A(n10310), .ZN(n10311) );
  BUF_X1 U4134 ( .A(n10316), .Z(n10312) );
  INV_X1 U4135 ( .A(n2158), .ZN(n10313) );
  INV_X1 U4136 ( .A(n10313), .ZN(n10314) );
  INV_X1 U4137 ( .A(n5709), .ZN(n10315) );
  INV_X1 U4138 ( .A(n10315), .ZN(n10316) );
  BUF_X1 U4139 ( .A(n10320), .Z(n10317) );
  INV_X1 U4140 ( .A(matrix_mul_2D_2__2__0_), .ZN(n10318) );
  INV_X1 U4141 ( .A(n5710), .ZN(n10319) );
  INV_X1 U4142 ( .A(n10319), .ZN(n10320) );
  BUF_X1 U4143 ( .A(n27444), .Z(n10321) );
  BUF_X1 U4144 ( .A(n27445), .Z(n10322) );
  BUF_X1 U4145 ( .A(n27446), .Z(n10323) );
  BUF_X1 U4146 ( .A(n27447), .Z(n10324) );
  BUF_X1 U4147 ( .A(n27448), .Z(n10325) );
  BUF_X1 U4148 ( .A(n27449), .Z(n10326) );
  BUF_X1 U4149 ( .A(n10331), .Z(n10327) );
  INV_X1 U4150 ( .A(n2130), .ZN(n10328) );
  INV_X1 U4151 ( .A(n10328), .ZN(n10329) );
  INV_X1 U4152 ( .A(n56810), .ZN(n10330) );
  INV_X1 U4153 ( .A(n10330), .ZN(n10331) );
  BUF_X1 U4154 ( .A(n10336), .Z(n10332) );
  INV_X1 U4155 ( .A(n2131), .ZN(n10333) );
  INV_X1 U4156 ( .A(n10333), .ZN(n10334) );
  INV_X1 U4157 ( .A(n56820), .ZN(n10335) );
  INV_X1 U4158 ( .A(n10335), .ZN(n10336) );
  BUF_X1 U4159 ( .A(n10341), .Z(n10337) );
  INV_X1 U4160 ( .A(n2132), .ZN(n10338) );
  INV_X1 U4161 ( .A(n10338), .ZN(n10339) );
  INV_X1 U4162 ( .A(n56830), .ZN(n10340) );
  INV_X1 U4163 ( .A(n10340), .ZN(n10341) );
  BUF_X1 U4164 ( .A(n10346), .Z(n10342) );
  INV_X1 U4165 ( .A(n2133), .ZN(n10343) );
  INV_X1 U4166 ( .A(n10343), .ZN(n10344) );
  INV_X1 U4167 ( .A(n56840), .ZN(n10345) );
  INV_X1 U4168 ( .A(n10345), .ZN(n10346) );
  BUF_X1 U4169 ( .A(n10351), .Z(n10347) );
  INV_X1 U4170 ( .A(n2134), .ZN(n10348) );
  INV_X1 U4171 ( .A(n10348), .ZN(n10349) );
  INV_X1 U4172 ( .A(n56850), .ZN(n10350) );
  INV_X1 U4173 ( .A(n10350), .ZN(n10351) );
  BUF_X1 U4174 ( .A(n10356), .Z(n10352) );
  INV_X1 U4175 ( .A(n2135), .ZN(n10353) );
  INV_X1 U4176 ( .A(n10353), .ZN(n10354) );
  INV_X1 U4177 ( .A(n56860), .ZN(n10355) );
  INV_X1 U4178 ( .A(n10355), .ZN(n10356) );
  BUF_X1 U4179 ( .A(n10361), .Z(n10357) );
  INV_X1 U4180 ( .A(n2136), .ZN(n10358) );
  INV_X1 U4181 ( .A(n10358), .ZN(n10359) );
  INV_X1 U4182 ( .A(n56870), .ZN(n10360) );
  INV_X1 U4183 ( .A(n10360), .ZN(n10361) );
  BUF_X1 U4184 ( .A(n10366), .Z(n10362) );
  INV_X1 U4185 ( .A(n2137), .ZN(n10363) );
  INV_X1 U4186 ( .A(n10363), .ZN(n10364) );
  INV_X1 U4187 ( .A(n56880), .ZN(n10365) );
  INV_X1 U4188 ( .A(n10365), .ZN(n10366) );
  BUF_X1 U4189 ( .A(n10371), .Z(n10367) );
  INV_X1 U4190 ( .A(n2138), .ZN(n10368) );
  INV_X1 U4191 ( .A(n10368), .ZN(n10369) );
  INV_X1 U4192 ( .A(n56890), .ZN(n10370) );
  INV_X1 U4193 ( .A(n10370), .ZN(n10371) );
  BUF_X1 U4194 ( .A(n10376), .Z(n10372) );
  INV_X1 U4195 ( .A(n2139), .ZN(n10373) );
  INV_X1 U4196 ( .A(n10373), .ZN(n10374) );
  INV_X1 U4197 ( .A(n56900), .ZN(n10375) );
  INV_X1 U4198 ( .A(n10375), .ZN(n10376) );
  BUF_X1 U4199 ( .A(n10381), .Z(n10377) );
  INV_X1 U4200 ( .A(n2140), .ZN(n10378) );
  INV_X1 U4201 ( .A(n10378), .ZN(n10379) );
  INV_X1 U4202 ( .A(n56910), .ZN(n10380) );
  INV_X1 U4203 ( .A(n10380), .ZN(n10381) );
  BUF_X1 U4204 ( .A(n10386), .Z(n10382) );
  INV_X1 U4205 ( .A(n2141), .ZN(n10383) );
  INV_X1 U4206 ( .A(n10383), .ZN(n10384) );
  INV_X1 U4207 ( .A(n56920), .ZN(n10385) );
  INV_X1 U4208 ( .A(n10385), .ZN(n10386) );
  BUF_X1 U4209 ( .A(n10391), .Z(n10387) );
  INV_X1 U4210 ( .A(n2142), .ZN(n10388) );
  INV_X1 U4211 ( .A(n10388), .ZN(n10389) );
  INV_X1 U4212 ( .A(n56930), .ZN(n10390) );
  INV_X1 U4213 ( .A(n10390), .ZN(n10391) );
  BUF_X1 U4214 ( .A(n10396), .Z(n10392) );
  INV_X1 U4215 ( .A(n2143), .ZN(n10393) );
  INV_X1 U4216 ( .A(n10393), .ZN(n10394) );
  INV_X1 U4217 ( .A(n56940), .ZN(n10395) );
  INV_X1 U4218 ( .A(n10395), .ZN(n10396) );
  BUF_X1 U4219 ( .A(n10400), .Z(n10397) );
  INV_X1 U4220 ( .A(matrix_mul_2D_2__1__0_), .ZN(n10398) );
  INV_X1 U4221 ( .A(n56950), .ZN(n10399) );
  INV_X1 U4222 ( .A(n10399), .ZN(n10400) );
  BUF_X1 U4223 ( .A(n27438), .Z(n10401) );
  BUF_X1 U4224 ( .A(n27439), .Z(n10402) );
  BUF_X1 U4225 ( .A(n274401), .Z(n10403) );
  BUF_X1 U4226 ( .A(n27441), .Z(n10404) );
  BUF_X1 U4227 ( .A(n27442), .Z(n10405) );
  BUF_X1 U4228 ( .A(n27443), .Z(n10406) );
  BUF_X1 U4229 ( .A(n10411), .Z(n10407) );
  INV_X1 U4230 ( .A(n2115), .ZN(n10408) );
  INV_X1 U4231 ( .A(n10408), .ZN(n10409) );
  INV_X1 U4232 ( .A(n5666), .ZN(n10410) );
  INV_X1 U4233 ( .A(n10410), .ZN(n10411) );
  BUF_X1 U4234 ( .A(n10416), .Z(n10412) );
  INV_X1 U4235 ( .A(n2116), .ZN(n10413) );
  INV_X1 U4236 ( .A(n10413), .ZN(n10414) );
  INV_X1 U4237 ( .A(n5667), .ZN(n10415) );
  INV_X1 U4238 ( .A(n10415), .ZN(n10416) );
  BUF_X1 U4239 ( .A(n10421), .Z(n10417) );
  INV_X1 U4240 ( .A(n2117), .ZN(n10418) );
  INV_X1 U4241 ( .A(n10418), .ZN(n10419) );
  INV_X1 U4242 ( .A(n5668), .ZN(n10420) );
  INV_X1 U4243 ( .A(n10420), .ZN(n10421) );
  BUF_X1 U4244 ( .A(n10426), .Z(n10422) );
  INV_X1 U4245 ( .A(n2118), .ZN(n10423) );
  INV_X1 U4246 ( .A(n10423), .ZN(n10424) );
  INV_X1 U4247 ( .A(n5669), .ZN(n10425) );
  INV_X1 U4248 ( .A(n10425), .ZN(n10426) );
  BUF_X1 U4249 ( .A(n10431), .Z(n10427) );
  INV_X1 U4250 ( .A(n2119), .ZN(n10428) );
  INV_X1 U4251 ( .A(n10428), .ZN(n10429) );
  INV_X1 U4252 ( .A(n5670), .ZN(n10430) );
  INV_X1 U4253 ( .A(n10430), .ZN(n10431) );
  BUF_X1 U4254 ( .A(n10436), .Z(n10432) );
  INV_X1 U4255 ( .A(n2120), .ZN(n10433) );
  INV_X1 U4256 ( .A(n10433), .ZN(n10434) );
  INV_X1 U4257 ( .A(n5671), .ZN(n10435) );
  INV_X1 U4258 ( .A(n10435), .ZN(n10436) );
  BUF_X1 U4259 ( .A(n10441), .Z(n10437) );
  INV_X1 U4260 ( .A(n2121), .ZN(n10438) );
  INV_X1 U4261 ( .A(n10438), .ZN(n10439) );
  INV_X1 U4262 ( .A(n5672), .ZN(n10440) );
  INV_X1 U4263 ( .A(n10440), .ZN(n10441) );
  BUF_X1 U4264 ( .A(n10446), .Z(n10442) );
  INV_X1 U4265 ( .A(n2122), .ZN(n10443) );
  INV_X1 U4266 ( .A(n10443), .ZN(n10444) );
  INV_X1 U4267 ( .A(n5673), .ZN(n10445) );
  INV_X1 U4268 ( .A(n10445), .ZN(n10446) );
  BUF_X1 U4269 ( .A(n10451), .Z(n10447) );
  INV_X1 U4270 ( .A(n2123), .ZN(n10448) );
  INV_X1 U4271 ( .A(n10448), .ZN(n10449) );
  INV_X1 U4272 ( .A(n5674), .ZN(n10450) );
  INV_X1 U4273 ( .A(n10450), .ZN(n10451) );
  BUF_X1 U4274 ( .A(n10456), .Z(n10452) );
  INV_X1 U4275 ( .A(n2124), .ZN(n10453) );
  INV_X1 U4276 ( .A(n10453), .ZN(n10454) );
  INV_X1 U4277 ( .A(n56750), .ZN(n10455) );
  INV_X1 U4278 ( .A(n10455), .ZN(n10456) );
  BUF_X1 U4279 ( .A(n10461), .Z(n10457) );
  INV_X1 U4280 ( .A(n2125), .ZN(n10458) );
  INV_X1 U4281 ( .A(n10458), .ZN(n10459) );
  INV_X1 U4282 ( .A(n56760), .ZN(n10460) );
  INV_X1 U4283 ( .A(n10460), .ZN(n10461) );
  BUF_X1 U4284 ( .A(n10466), .Z(n10462) );
  INV_X1 U4285 ( .A(n2126), .ZN(n10463) );
  INV_X1 U4286 ( .A(n10463), .ZN(n10464) );
  INV_X1 U4287 ( .A(n56770), .ZN(n10465) );
  INV_X1 U4288 ( .A(n10465), .ZN(n10466) );
  BUF_X1 U4289 ( .A(n10471), .Z(n10467) );
  INV_X1 U4290 ( .A(n2127), .ZN(n10468) );
  INV_X1 U4291 ( .A(n10468), .ZN(n10469) );
  INV_X1 U4292 ( .A(n56780), .ZN(n10470) );
  INV_X1 U4293 ( .A(n10470), .ZN(n10471) );
  BUF_X1 U4294 ( .A(n10476), .Z(n10472) );
  INV_X1 U4295 ( .A(n2128), .ZN(n10473) );
  INV_X1 U4296 ( .A(n10473), .ZN(n10474) );
  INV_X1 U4297 ( .A(n56790), .ZN(n10475) );
  INV_X1 U4298 ( .A(n10475), .ZN(n10476) );
  BUF_X1 U4299 ( .A(n10480), .Z(n10477) );
  INV_X1 U4300 ( .A(matrix_mul_2D_2__0__0_), .ZN(n10478) );
  INV_X1 U4301 ( .A(n56800), .ZN(n10479) );
  INV_X1 U4302 ( .A(n10479), .ZN(n10480) );
  BUF_X1 U4303 ( .A(n27432), .Z(n10481) );
  BUF_X1 U4304 ( .A(n27433), .Z(n10482) );
  BUF_X1 U4305 ( .A(n27434), .Z(n10483) );
  BUF_X1 U4306 ( .A(n27435), .Z(n10484) );
  BUF_X1 U4307 ( .A(n27436), .Z(n10485) );
  BUF_X1 U4308 ( .A(n27437), .Z(n10486) );
  BUF_X1 U4309 ( .A(n10491), .Z(n10487) );
  INV_X1 U4310 ( .A(n2100), .ZN(n10488) );
  INV_X1 U4311 ( .A(n10488), .ZN(n10489) );
  INV_X1 U4312 ( .A(n56510), .ZN(n10490) );
  INV_X1 U4313 ( .A(n10490), .ZN(n10491) );
  BUF_X1 U4314 ( .A(n10496), .Z(n10492) );
  INV_X1 U4315 ( .A(n2101), .ZN(n10493) );
  INV_X1 U4316 ( .A(n10493), .ZN(n10494) );
  INV_X1 U4317 ( .A(n56520), .ZN(n10495) );
  INV_X1 U4318 ( .A(n10495), .ZN(n10496) );
  BUF_X1 U4319 ( .A(n10501), .Z(n10497) );
  INV_X1 U4320 ( .A(n2102), .ZN(n10498) );
  INV_X1 U4321 ( .A(n10498), .ZN(n10499) );
  INV_X1 U4322 ( .A(n56530), .ZN(n10500) );
  INV_X1 U4323 ( .A(n10500), .ZN(n10501) );
  BUF_X1 U4324 ( .A(n10506), .Z(n10502) );
  INV_X1 U4325 ( .A(n2103), .ZN(n10503) );
  INV_X1 U4326 ( .A(n10503), .ZN(n10504) );
  INV_X1 U4327 ( .A(n56540), .ZN(n10505) );
  INV_X1 U4328 ( .A(n10505), .ZN(n10506) );
  BUF_X1 U4329 ( .A(n10511), .Z(n10507) );
  INV_X1 U4330 ( .A(n2104), .ZN(n10508) );
  INV_X1 U4331 ( .A(n10508), .ZN(n10509) );
  INV_X1 U4332 ( .A(n56550), .ZN(n10510) );
  INV_X1 U4333 ( .A(n10510), .ZN(n10511) );
  BUF_X1 U4334 ( .A(n10516), .Z(n10512) );
  INV_X1 U4335 ( .A(n2105), .ZN(n10513) );
  INV_X1 U4336 ( .A(n10513), .ZN(n10514) );
  INV_X1 U4337 ( .A(n56560), .ZN(n10515) );
  INV_X1 U4338 ( .A(n10515), .ZN(n10516) );
  BUF_X1 U4339 ( .A(n10521), .Z(n10517) );
  INV_X1 U4340 ( .A(n2106), .ZN(n10518) );
  INV_X1 U4341 ( .A(n10518), .ZN(n10519) );
  INV_X1 U4342 ( .A(n56570), .ZN(n10520) );
  INV_X1 U4343 ( .A(n10520), .ZN(n10521) );
  BUF_X1 U4344 ( .A(n10526), .Z(n10522) );
  INV_X1 U4345 ( .A(n2107), .ZN(n10523) );
  INV_X1 U4346 ( .A(n10523), .ZN(n10524) );
  INV_X1 U4347 ( .A(n5658), .ZN(n10525) );
  INV_X1 U4348 ( .A(n10525), .ZN(n10526) );
  BUF_X1 U4349 ( .A(n10531), .Z(n10527) );
  INV_X1 U4350 ( .A(n2108), .ZN(n10528) );
  INV_X1 U4351 ( .A(n10528), .ZN(n10529) );
  INV_X1 U4352 ( .A(n5659), .ZN(n10530) );
  INV_X1 U4353 ( .A(n10530), .ZN(n10531) );
  BUF_X1 U4354 ( .A(n10536), .Z(n10532) );
  INV_X1 U4355 ( .A(n2109), .ZN(n10533) );
  INV_X1 U4356 ( .A(n10533), .ZN(n10534) );
  INV_X1 U4357 ( .A(n5660), .ZN(n10535) );
  INV_X1 U4358 ( .A(n10535), .ZN(n10536) );
  BUF_X1 U4359 ( .A(n10541), .Z(n10537) );
  INV_X1 U4360 ( .A(n2110), .ZN(n10538) );
  INV_X1 U4361 ( .A(n10538), .ZN(n10539) );
  INV_X1 U4362 ( .A(n5661), .ZN(n10540) );
  INV_X1 U4363 ( .A(n10540), .ZN(n10541) );
  BUF_X1 U4364 ( .A(n10546), .Z(n10542) );
  INV_X1 U4365 ( .A(n2111), .ZN(n10543) );
  INV_X1 U4366 ( .A(n10543), .ZN(n10544) );
  INV_X1 U4367 ( .A(n5662), .ZN(n10545) );
  INV_X1 U4368 ( .A(n10545), .ZN(n10546) );
  BUF_X1 U4369 ( .A(n10551), .Z(n10547) );
  INV_X1 U4370 ( .A(n2112), .ZN(n10548) );
  INV_X1 U4371 ( .A(n10548), .ZN(n10549) );
  INV_X1 U4372 ( .A(n5663), .ZN(n10550) );
  INV_X1 U4373 ( .A(n10550), .ZN(n10551) );
  BUF_X1 U4374 ( .A(n10556), .Z(n10552) );
  INV_X1 U4375 ( .A(n2113), .ZN(n10553) );
  INV_X1 U4376 ( .A(n10553), .ZN(n10554) );
  INV_X1 U4377 ( .A(n5664), .ZN(n10555) );
  INV_X1 U4378 ( .A(n10555), .ZN(n10556) );
  BUF_X1 U4379 ( .A(n10560), .Z(n10557) );
  INV_X1 U4380 ( .A(matrix_mul_2D_1__7__0_), .ZN(n10558) );
  INV_X1 U4381 ( .A(n5665), .ZN(n10559) );
  INV_X1 U4382 ( .A(n10559), .ZN(n10560) );
  BUF_X1 U4383 ( .A(n27426), .Z(n10561) );
  BUF_X1 U4384 ( .A(n27427), .Z(n10562) );
  BUF_X1 U4385 ( .A(n27428), .Z(n10563) );
  BUF_X1 U4386 ( .A(n27429), .Z(n10564) );
  BUF_X1 U4387 ( .A(n274301), .Z(n10565) );
  BUF_X1 U4388 ( .A(n27431), .Z(n10566) );
  BUF_X1 U4389 ( .A(n10571), .Z(n10567) );
  INV_X1 U4390 ( .A(n2085), .ZN(n10568) );
  INV_X1 U4391 ( .A(n10568), .ZN(n10569) );
  INV_X1 U4392 ( .A(n5636), .ZN(n10570) );
  INV_X1 U4393 ( .A(n10570), .ZN(n10571) );
  BUF_X1 U4394 ( .A(n10576), .Z(n10572) );
  INV_X1 U4395 ( .A(n2086), .ZN(n10573) );
  INV_X1 U4396 ( .A(n10573), .ZN(n10574) );
  INV_X1 U4397 ( .A(n5637), .ZN(n10575) );
  INV_X1 U4398 ( .A(n10575), .ZN(n10576) );
  BUF_X1 U4399 ( .A(n10581), .Z(n10577) );
  INV_X1 U4400 ( .A(n2087), .ZN(n10578) );
  INV_X1 U4401 ( .A(n10578), .ZN(n10579) );
  INV_X1 U4402 ( .A(n5638), .ZN(n10580) );
  INV_X1 U4403 ( .A(n10580), .ZN(n10581) );
  BUF_X1 U4404 ( .A(n10586), .Z(n10582) );
  INV_X1 U4405 ( .A(n2088), .ZN(n10583) );
  INV_X1 U4406 ( .A(n10583), .ZN(n10584) );
  INV_X1 U4407 ( .A(n5639), .ZN(n10585) );
  INV_X1 U4408 ( .A(n10585), .ZN(n10586) );
  BUF_X1 U4409 ( .A(n10591), .Z(n10587) );
  INV_X1 U4410 ( .A(n2089), .ZN(n10588) );
  INV_X1 U4411 ( .A(n10588), .ZN(n10589) );
  INV_X1 U4412 ( .A(n5640), .ZN(n10590) );
  INV_X1 U4413 ( .A(n10590), .ZN(n10591) );
  BUF_X1 U4414 ( .A(n10596), .Z(n10592) );
  INV_X1 U4415 ( .A(n2090), .ZN(n10593) );
  INV_X1 U4416 ( .A(n10593), .ZN(n10594) );
  INV_X1 U4417 ( .A(n5641), .ZN(n10595) );
  INV_X1 U4418 ( .A(n10595), .ZN(n10596) );
  BUF_X1 U4419 ( .A(n10601), .Z(n10597) );
  INV_X1 U4420 ( .A(n2091), .ZN(n10598) );
  INV_X1 U4421 ( .A(n10598), .ZN(n10599) );
  INV_X1 U4422 ( .A(n56420), .ZN(n10600) );
  INV_X1 U4423 ( .A(n10600), .ZN(n10601) );
  BUF_X1 U4424 ( .A(n10606), .Z(n10602) );
  INV_X1 U4425 ( .A(n2092), .ZN(n10603) );
  INV_X1 U4426 ( .A(n10603), .ZN(n10604) );
  INV_X1 U4427 ( .A(n56430), .ZN(n10605) );
  INV_X1 U4428 ( .A(n10605), .ZN(n10606) );
  BUF_X1 U4429 ( .A(n10611), .Z(n10607) );
  INV_X1 U4430 ( .A(n2093), .ZN(n10608) );
  INV_X1 U4431 ( .A(n10608), .ZN(n10609) );
  INV_X1 U4432 ( .A(n56440), .ZN(n10610) );
  INV_X1 U4433 ( .A(n10610), .ZN(n10611) );
  BUF_X1 U4434 ( .A(n10616), .Z(n10612) );
  INV_X1 U4435 ( .A(n2094), .ZN(n10613) );
  INV_X1 U4436 ( .A(n10613), .ZN(n10614) );
  INV_X1 U4437 ( .A(n56450), .ZN(n10615) );
  INV_X1 U4438 ( .A(n10615), .ZN(n10616) );
  BUF_X1 U4439 ( .A(n10621), .Z(n10617) );
  INV_X1 U4440 ( .A(n2095), .ZN(n10618) );
  INV_X1 U4441 ( .A(n10618), .ZN(n10619) );
  INV_X1 U4442 ( .A(n56460), .ZN(n10620) );
  INV_X1 U4443 ( .A(n10620), .ZN(n10621) );
  BUF_X1 U4444 ( .A(n10626), .Z(n10622) );
  INV_X1 U4445 ( .A(n2096), .ZN(n10623) );
  INV_X1 U4446 ( .A(n10623), .ZN(n10624) );
  INV_X1 U4447 ( .A(n56470), .ZN(n10625) );
  INV_X1 U4448 ( .A(n10625), .ZN(n10626) );
  BUF_X1 U4449 ( .A(n10631), .Z(n10627) );
  INV_X1 U4450 ( .A(n2097), .ZN(n10628) );
  INV_X1 U4451 ( .A(n10628), .ZN(n10629) );
  INV_X1 U4452 ( .A(n56480), .ZN(n10630) );
  INV_X1 U4453 ( .A(n10630), .ZN(n10631) );
  BUF_X1 U4454 ( .A(n10636), .Z(n10632) );
  INV_X1 U4455 ( .A(n2098), .ZN(n10633) );
  INV_X1 U4456 ( .A(n10633), .ZN(n10634) );
  INV_X1 U4457 ( .A(n56490), .ZN(n10635) );
  INV_X1 U4458 ( .A(n10635), .ZN(n10636) );
  BUF_X1 U4459 ( .A(n10640), .Z(n10637) );
  INV_X1 U4460 ( .A(matrix_mul_2D_1__6__0_), .ZN(n10638) );
  INV_X1 U4461 ( .A(n56500), .ZN(n10639) );
  INV_X1 U4462 ( .A(n10639), .ZN(n10640) );
  BUF_X1 U4463 ( .A(n10643), .Z(n10641) );
  INV_X1 U4464 ( .A(n274201), .ZN(n10642) );
  INV_X1 U4465 ( .A(n10642), .ZN(n10643) );
  BUF_X1 U4466 ( .A(n10646), .Z(n10644) );
  INV_X1 U4467 ( .A(n27421), .ZN(n10645) );
  INV_X1 U4468 ( .A(n10645), .ZN(n10646) );
  BUF_X1 U4469 ( .A(n10649), .Z(n10647) );
  INV_X1 U4470 ( .A(n27422), .ZN(n10648) );
  INV_X1 U4471 ( .A(n10648), .ZN(n10649) );
  BUF_X1 U4472 ( .A(n10652), .Z(n10650) );
  INV_X1 U4473 ( .A(n27423), .ZN(n10651) );
  INV_X1 U4474 ( .A(n10651), .ZN(n10652) );
  BUF_X1 U4475 ( .A(n10655), .Z(n10653) );
  INV_X1 U4476 ( .A(n27424), .ZN(n10654) );
  INV_X1 U4477 ( .A(n10654), .ZN(n10655) );
  BUF_X1 U4478 ( .A(n10658), .Z(n10656) );
  INV_X1 U4479 ( .A(n27425), .ZN(n10657) );
  INV_X1 U4480 ( .A(n10657), .ZN(n10658) );
  BUF_X1 U4481 ( .A(n10662), .Z(n10659) );
  INV_X1 U4482 ( .A(matrix_mul_2D_1__5__14_), .ZN(n10660) );
  INV_X1 U4483 ( .A(n5621), .ZN(n10661) );
  INV_X1 U4484 ( .A(n10661), .ZN(n10662) );
  BUF_X1 U4485 ( .A(n10666), .Z(n10663) );
  INV_X1 U4486 ( .A(matrix_mul_2D_1__5__13_), .ZN(n10664) );
  INV_X1 U4487 ( .A(n5622), .ZN(n10665) );
  INV_X1 U4488 ( .A(n10665), .ZN(n10666) );
  BUF_X1 U4489 ( .A(n10670), .Z(n10667) );
  INV_X1 U4490 ( .A(matrix_mul_2D_1__5__12_), .ZN(n10668) );
  INV_X1 U4491 ( .A(n5623), .ZN(n10669) );
  INV_X1 U4492 ( .A(n10669), .ZN(n10670) );
  BUF_X1 U4493 ( .A(n10674), .Z(n10671) );
  INV_X1 U4494 ( .A(matrix_mul_2D_1__5__11_), .ZN(n10672) );
  INV_X1 U4495 ( .A(n5624), .ZN(n10673) );
  INV_X1 U4496 ( .A(n10673), .ZN(n10674) );
  BUF_X1 U4497 ( .A(n10678), .Z(n10675) );
  INV_X1 U4498 ( .A(matrix_mul_2D_1__5__10_), .ZN(n10676) );
  INV_X1 U4499 ( .A(n5625), .ZN(n10677) );
  INV_X1 U4500 ( .A(n10677), .ZN(n10678) );
  BUF_X1 U4501 ( .A(n10682), .Z(n10679) );
  INV_X1 U4502 ( .A(matrix_mul_2D_1__5__9_), .ZN(n10680) );
  INV_X1 U4503 ( .A(n5626), .ZN(n10681) );
  INV_X1 U4504 ( .A(n10681), .ZN(n10682) );
  BUF_X1 U4505 ( .A(n10686), .Z(n10683) );
  INV_X1 U4506 ( .A(matrix_mul_2D_1__5__8_), .ZN(n10684) );
  INV_X1 U4507 ( .A(n5627), .ZN(n10685) );
  INV_X1 U4508 ( .A(n10685), .ZN(n10686) );
  BUF_X1 U4509 ( .A(n10690), .Z(n10687) );
  INV_X1 U4510 ( .A(matrix_mul_2D_1__5__7_), .ZN(n10688) );
  INV_X1 U4511 ( .A(n5628), .ZN(n10689) );
  INV_X1 U4512 ( .A(n10689), .ZN(n10690) );
  BUF_X1 U4513 ( .A(n10694), .Z(n10691) );
  INV_X1 U4514 ( .A(matrix_mul_2D_1__5__6_), .ZN(n10692) );
  INV_X1 U4515 ( .A(n5629), .ZN(n10693) );
  INV_X1 U4516 ( .A(n10693), .ZN(n10694) );
  BUF_X1 U4517 ( .A(n10698), .Z(n10695) );
  INV_X1 U4518 ( .A(matrix_mul_2D_1__5__5_), .ZN(n10696) );
  INV_X1 U4519 ( .A(n5630), .ZN(n10697) );
  INV_X1 U4520 ( .A(n10697), .ZN(n10698) );
  BUF_X1 U4521 ( .A(n10702), .Z(n10699) );
  INV_X1 U4522 ( .A(matrix_mul_2D_1__5__4_), .ZN(n10700) );
  INV_X1 U4523 ( .A(n5631), .ZN(n10701) );
  INV_X1 U4524 ( .A(n10701), .ZN(n10702) );
  BUF_X1 U4525 ( .A(n10706), .Z(n10703) );
  INV_X1 U4526 ( .A(matrix_mul_2D_1__5__3_), .ZN(n10704) );
  INV_X1 U4527 ( .A(n5632), .ZN(n10705) );
  INV_X1 U4528 ( .A(n10705), .ZN(n10706) );
  BUF_X1 U4529 ( .A(n10710), .Z(n10707) );
  INV_X1 U4530 ( .A(matrix_mul_2D_1__5__2_), .ZN(n10708) );
  INV_X1 U4531 ( .A(n5633), .ZN(n10709) );
  INV_X1 U4532 ( .A(n10709), .ZN(n10710) );
  BUF_X1 U4533 ( .A(n10714), .Z(n10711) );
  INV_X1 U4534 ( .A(matrix_mul_2D_1__5__1_), .ZN(n10712) );
  INV_X1 U4535 ( .A(n5634), .ZN(n10713) );
  INV_X1 U4536 ( .A(n10713), .ZN(n10714) );
  BUF_X1 U4537 ( .A(n10719), .Z(n10715) );
  INV_X1 U4538 ( .A(n2084), .ZN(n10716) );
  INV_X1 U4539 ( .A(n10716), .ZN(n10717) );
  INV_X1 U4540 ( .A(n5635), .ZN(n10718) );
  INV_X1 U4541 ( .A(n10718), .ZN(n10719) );
  BUF_X1 U4542 ( .A(n10722), .Z(n10720) );
  INV_X1 U4543 ( .A(n27414), .ZN(n10721) );
  INV_X1 U4544 ( .A(n10721), .ZN(n10722) );
  BUF_X1 U4545 ( .A(n10725), .Z(n10723) );
  INV_X1 U4546 ( .A(n27415), .ZN(n10724) );
  INV_X1 U4547 ( .A(n10724), .ZN(n10725) );
  BUF_X1 U4548 ( .A(n10728), .Z(n10726) );
  INV_X1 U4549 ( .A(n27416), .ZN(n10727) );
  INV_X1 U4550 ( .A(n10727), .ZN(n10728) );
  BUF_X1 U4551 ( .A(n10731), .Z(n10729) );
  INV_X1 U4552 ( .A(n27417), .ZN(n10730) );
  INV_X1 U4553 ( .A(n10730), .ZN(n10731) );
  BUF_X1 U4554 ( .A(n10734), .Z(n10732) );
  INV_X1 U4555 ( .A(n27418), .ZN(n10733) );
  INV_X1 U4556 ( .A(n10733), .ZN(n10734) );
  BUF_X1 U4557 ( .A(n10737), .Z(n10735) );
  INV_X1 U4558 ( .A(n27419), .ZN(n10736) );
  INV_X1 U4559 ( .A(n10736), .ZN(n10737) );
  BUF_X1 U4560 ( .A(n10741), .Z(n10738) );
  INV_X1 U4561 ( .A(matrix_mul_2D_1__4__14_), .ZN(n10739) );
  INV_X1 U4562 ( .A(n56060), .ZN(n10740) );
  INV_X1 U4563 ( .A(n10740), .ZN(n10741) );
  BUF_X1 U4564 ( .A(n10745), .Z(n10742) );
  INV_X1 U4565 ( .A(matrix_mul_2D_1__4__13_), .ZN(n10743) );
  INV_X1 U4566 ( .A(n5607), .ZN(n10744) );
  INV_X1 U4567 ( .A(n10744), .ZN(n10745) );
  BUF_X1 U4568 ( .A(n10749), .Z(n10746) );
  INV_X1 U4569 ( .A(matrix_mul_2D_1__4__12_), .ZN(n10747) );
  INV_X1 U4570 ( .A(n5608), .ZN(n10748) );
  INV_X1 U4571 ( .A(n10748), .ZN(n10749) );
  BUF_X1 U4572 ( .A(n10753), .Z(n10750) );
  INV_X1 U4573 ( .A(matrix_mul_2D_1__4__11_), .ZN(n10751) );
  INV_X1 U4574 ( .A(n5609), .ZN(n10752) );
  INV_X1 U4575 ( .A(n10752), .ZN(n10753) );
  BUF_X1 U4576 ( .A(n10757), .Z(n10754) );
  INV_X1 U4577 ( .A(matrix_mul_2D_1__4__10_), .ZN(n10755) );
  INV_X1 U4578 ( .A(n5610), .ZN(n10756) );
  INV_X1 U4579 ( .A(n10756), .ZN(n10757) );
  BUF_X1 U4580 ( .A(n10761), .Z(n10758) );
  INV_X1 U4581 ( .A(matrix_mul_2D_1__4__9_), .ZN(n10759) );
  INV_X1 U4582 ( .A(n5611), .ZN(n10760) );
  INV_X1 U4583 ( .A(n10760), .ZN(n10761) );
  BUF_X1 U4584 ( .A(n10765), .Z(n10762) );
  INV_X1 U4585 ( .A(matrix_mul_2D_1__4__8_), .ZN(n10763) );
  INV_X1 U4586 ( .A(n5612), .ZN(n10764) );
  INV_X1 U4587 ( .A(n10764), .ZN(n10765) );
  BUF_X1 U4588 ( .A(n10769), .Z(n10766) );
  INV_X1 U4589 ( .A(matrix_mul_2D_1__4__7_), .ZN(n10767) );
  INV_X1 U4590 ( .A(n5613), .ZN(n10768) );
  INV_X1 U4591 ( .A(n10768), .ZN(n10769) );
  BUF_X1 U4592 ( .A(n10773), .Z(n10770) );
  INV_X1 U4593 ( .A(matrix_mul_2D_1__4__6_), .ZN(n10771) );
  INV_X1 U4594 ( .A(n5614), .ZN(n10772) );
  INV_X1 U4595 ( .A(n10772), .ZN(n10773) );
  BUF_X1 U4596 ( .A(n10777), .Z(n10774) );
  INV_X1 U4597 ( .A(matrix_mul_2D_1__4__5_), .ZN(n10775) );
  INV_X1 U4598 ( .A(n5615), .ZN(n10776) );
  INV_X1 U4599 ( .A(n10776), .ZN(n10777) );
  BUF_X1 U4600 ( .A(n10781), .Z(n10778) );
  INV_X1 U4601 ( .A(matrix_mul_2D_1__4__4_), .ZN(n10779) );
  INV_X1 U4602 ( .A(n5616), .ZN(n10780) );
  INV_X1 U4603 ( .A(n10780), .ZN(n10781) );
  BUF_X1 U4604 ( .A(n10785), .Z(n10782) );
  INV_X1 U4605 ( .A(matrix_mul_2D_1__4__3_), .ZN(n10783) );
  INV_X1 U4606 ( .A(n5617), .ZN(n10784) );
  INV_X1 U4607 ( .A(n10784), .ZN(n10785) );
  BUF_X1 U4608 ( .A(n10789), .Z(n10786) );
  INV_X1 U4609 ( .A(matrix_mul_2D_1__4__2_), .ZN(n10787) );
  INV_X1 U4610 ( .A(n5618), .ZN(n10788) );
  INV_X1 U4611 ( .A(n10788), .ZN(n10789) );
  BUF_X1 U4612 ( .A(n10793), .Z(n10790) );
  INV_X1 U4613 ( .A(matrix_mul_2D_1__4__1_), .ZN(n10791) );
  INV_X1 U4614 ( .A(n5619), .ZN(n10792) );
  INV_X1 U4615 ( .A(n10792), .ZN(n10793) );
  BUF_X1 U4616 ( .A(n10798), .Z(n10794) );
  INV_X1 U4617 ( .A(n2063), .ZN(n10795) );
  INV_X1 U4618 ( .A(n10795), .ZN(n10796) );
  INV_X1 U4619 ( .A(n5620), .ZN(n10797) );
  INV_X1 U4620 ( .A(n10797), .ZN(n10798) );
  BUF_X1 U4621 ( .A(n10801), .Z(n10799) );
  INV_X1 U4622 ( .A(n27408), .ZN(n10800) );
  INV_X1 U4623 ( .A(n10800), .ZN(n10801) );
  BUF_X1 U4624 ( .A(n10804), .Z(n10802) );
  INV_X1 U4625 ( .A(n27409), .ZN(n10803) );
  INV_X1 U4626 ( .A(n10803), .ZN(n10804) );
  BUF_X1 U4627 ( .A(n10807), .Z(n10805) );
  INV_X1 U4628 ( .A(n274101), .ZN(n10806) );
  INV_X1 U4629 ( .A(n10806), .ZN(n10807) );
  BUF_X1 U4630 ( .A(n10810), .Z(n10808) );
  INV_X1 U4631 ( .A(n27411), .ZN(n10809) );
  INV_X1 U4632 ( .A(n10809), .ZN(n10810) );
  BUF_X1 U4633 ( .A(n10813), .Z(n10811) );
  INV_X1 U4634 ( .A(n27412), .ZN(n10812) );
  INV_X1 U4635 ( .A(n10812), .ZN(n10813) );
  BUF_X1 U4636 ( .A(n10816), .Z(n10814) );
  INV_X1 U4637 ( .A(n27413), .ZN(n10815) );
  INV_X1 U4638 ( .A(n10815), .ZN(n10816) );
  BUF_X1 U4639 ( .A(n10820), .Z(n10817) );
  INV_X1 U4640 ( .A(matrix_mul_2D_1__3__14_), .ZN(n10818) );
  INV_X1 U4641 ( .A(n55910), .ZN(n10819) );
  INV_X1 U4642 ( .A(n10819), .ZN(n10820) );
  BUF_X1 U4643 ( .A(n10824), .Z(n10821) );
  INV_X1 U4644 ( .A(matrix_mul_2D_1__3__13_), .ZN(n10822) );
  INV_X1 U4645 ( .A(n55920), .ZN(n10823) );
  INV_X1 U4646 ( .A(n10823), .ZN(n10824) );
  BUF_X1 U4647 ( .A(n10828), .Z(n10825) );
  INV_X1 U4648 ( .A(matrix_mul_2D_1__3__12_), .ZN(n10826) );
  INV_X1 U4649 ( .A(n55930), .ZN(n10827) );
  INV_X1 U4650 ( .A(n10827), .ZN(n10828) );
  BUF_X1 U4651 ( .A(n10832), .Z(n10829) );
  INV_X1 U4652 ( .A(matrix_mul_2D_1__3__11_), .ZN(n10830) );
  INV_X1 U4653 ( .A(n55940), .ZN(n10831) );
  INV_X1 U4654 ( .A(n10831), .ZN(n10832) );
  BUF_X1 U4655 ( .A(n10836), .Z(n10833) );
  INV_X1 U4656 ( .A(matrix_mul_2D_1__3__10_), .ZN(n10834) );
  INV_X1 U4657 ( .A(n55950), .ZN(n10835) );
  INV_X1 U4658 ( .A(n10835), .ZN(n10836) );
  BUF_X1 U4659 ( .A(n10840), .Z(n10837) );
  INV_X1 U4660 ( .A(matrix_mul_2D_1__3__9_), .ZN(n10838) );
  INV_X1 U4661 ( .A(n55960), .ZN(n10839) );
  INV_X1 U4662 ( .A(n10839), .ZN(n10840) );
  BUF_X1 U4663 ( .A(n10844), .Z(n10841) );
  INV_X1 U4664 ( .A(matrix_mul_2D_1__3__8_), .ZN(n10842) );
  INV_X1 U4665 ( .A(n55970), .ZN(n10843) );
  INV_X1 U4666 ( .A(n10843), .ZN(n10844) );
  BUF_X1 U4667 ( .A(n10848), .Z(n10845) );
  INV_X1 U4668 ( .A(matrix_mul_2D_1__3__7_), .ZN(n10846) );
  INV_X1 U4669 ( .A(n55980), .ZN(n10847) );
  INV_X1 U4670 ( .A(n10847), .ZN(n10848) );
  BUF_X1 U4671 ( .A(n10852), .Z(n10849) );
  INV_X1 U4672 ( .A(matrix_mul_2D_1__3__6_), .ZN(n10850) );
  INV_X1 U4673 ( .A(n55990), .ZN(n10851) );
  INV_X1 U4674 ( .A(n10851), .ZN(n10852) );
  BUF_X1 U4675 ( .A(n10856), .Z(n10853) );
  INV_X1 U4676 ( .A(matrix_mul_2D_1__3__5_), .ZN(n10854) );
  INV_X1 U4677 ( .A(n56000), .ZN(n10855) );
  INV_X1 U4678 ( .A(n10855), .ZN(n10856) );
  BUF_X1 U4679 ( .A(n10860), .Z(n10857) );
  INV_X1 U4680 ( .A(matrix_mul_2D_1__3__4_), .ZN(n10858) );
  INV_X1 U4681 ( .A(n56010), .ZN(n10859) );
  INV_X1 U4682 ( .A(n10859), .ZN(n10860) );
  BUF_X1 U4683 ( .A(n10864), .Z(n10861) );
  INV_X1 U4684 ( .A(matrix_mul_2D_1__3__3_), .ZN(n10862) );
  INV_X1 U4685 ( .A(n56020), .ZN(n10863) );
  INV_X1 U4686 ( .A(n10863), .ZN(n10864) );
  BUF_X1 U4687 ( .A(n10868), .Z(n10865) );
  INV_X1 U4688 ( .A(matrix_mul_2D_1__3__2_), .ZN(n10866) );
  INV_X1 U4689 ( .A(n56030), .ZN(n10867) );
  INV_X1 U4690 ( .A(n10867), .ZN(n10868) );
  BUF_X1 U4691 ( .A(n10872), .Z(n10869) );
  INV_X1 U4692 ( .A(matrix_mul_2D_1__3__1_), .ZN(n10870) );
  INV_X1 U4693 ( .A(n56040), .ZN(n10871) );
  INV_X1 U4694 ( .A(n10871), .ZN(n10872) );
  BUF_X1 U4695 ( .A(n10877), .Z(n10873) );
  INV_X1 U4696 ( .A(n2042), .ZN(n10874) );
  INV_X1 U4697 ( .A(n10874), .ZN(n10875) );
  INV_X1 U4698 ( .A(n56050), .ZN(n10876) );
  INV_X1 U4699 ( .A(n10876), .ZN(n10877) );
  BUF_X1 U4700 ( .A(n10880), .Z(n10878) );
  INV_X1 U4701 ( .A(n27402), .ZN(n10879) );
  INV_X1 U4702 ( .A(n10879), .ZN(n10880) );
  BUF_X1 U4703 ( .A(n10883), .Z(n10881) );
  INV_X1 U4704 ( .A(n27403), .ZN(n10882) );
  INV_X1 U4705 ( .A(n10882), .ZN(n10883) );
  BUF_X1 U4706 ( .A(n10886), .Z(n10884) );
  INV_X1 U4707 ( .A(n27404), .ZN(n10885) );
  INV_X1 U4708 ( .A(n10885), .ZN(n10886) );
  BUF_X1 U4709 ( .A(n10889), .Z(n10887) );
  INV_X1 U4710 ( .A(n27405), .ZN(n10888) );
  INV_X1 U4711 ( .A(n10888), .ZN(n10889) );
  BUF_X1 U4712 ( .A(n10892), .Z(n10890) );
  INV_X1 U4713 ( .A(n27406), .ZN(n10891) );
  INV_X1 U4714 ( .A(n10891), .ZN(n10892) );
  BUF_X1 U4715 ( .A(n10895), .Z(n10893) );
  INV_X1 U4716 ( .A(n27407), .ZN(n10894) );
  INV_X1 U4717 ( .A(n10894), .ZN(n10895) );
  BUF_X1 U4718 ( .A(n10899), .Z(n10896) );
  INV_X1 U4719 ( .A(matrix_mul_2D_1__2__14_), .ZN(n10897) );
  INV_X1 U4720 ( .A(n5576), .ZN(n10898) );
  INV_X1 U4721 ( .A(n10898), .ZN(n10899) );
  BUF_X1 U4722 ( .A(n10903), .Z(n10900) );
  INV_X1 U4723 ( .A(matrix_mul_2D_1__2__13_), .ZN(n10901) );
  INV_X1 U4724 ( .A(n5577), .ZN(n10902) );
  INV_X1 U4725 ( .A(n10902), .ZN(n10903) );
  BUF_X1 U4726 ( .A(n10907), .Z(n10904) );
  INV_X1 U4727 ( .A(matrix_mul_2D_1__2__12_), .ZN(n10905) );
  INV_X1 U4728 ( .A(n5578), .ZN(n10906) );
  INV_X1 U4729 ( .A(n10906), .ZN(n10907) );
  BUF_X1 U4730 ( .A(n10911), .Z(n10908) );
  INV_X1 U4731 ( .A(matrix_mul_2D_1__2__11_), .ZN(n10909) );
  INV_X1 U4732 ( .A(n5579), .ZN(n10910) );
  INV_X1 U4733 ( .A(n10910), .ZN(n10911) );
  BUF_X1 U4734 ( .A(n10915), .Z(n10912) );
  INV_X1 U4735 ( .A(matrix_mul_2D_1__2__10_), .ZN(n10913) );
  INV_X1 U4736 ( .A(n5580), .ZN(n10914) );
  INV_X1 U4737 ( .A(n10914), .ZN(n10915) );
  BUF_X1 U4738 ( .A(n10919), .Z(n10916) );
  INV_X1 U4739 ( .A(matrix_mul_2D_1__2__9_), .ZN(n10917) );
  INV_X1 U4740 ( .A(n5581), .ZN(n10918) );
  INV_X1 U4741 ( .A(n10918), .ZN(n10919) );
  BUF_X1 U4742 ( .A(n10923), .Z(n10920) );
  INV_X1 U4743 ( .A(matrix_mul_2D_1__2__8_), .ZN(n10921) );
  INV_X1 U4744 ( .A(n5582), .ZN(n10922) );
  INV_X1 U4745 ( .A(n10922), .ZN(n10923) );
  BUF_X1 U4746 ( .A(n10927), .Z(n10924) );
  INV_X1 U4747 ( .A(matrix_mul_2D_1__2__7_), .ZN(n10925) );
  INV_X1 U4748 ( .A(n5583), .ZN(n10926) );
  INV_X1 U4749 ( .A(n10926), .ZN(n10927) );
  BUF_X1 U4750 ( .A(n10931), .Z(n10928) );
  INV_X1 U4751 ( .A(matrix_mul_2D_1__2__6_), .ZN(n10929) );
  INV_X1 U4752 ( .A(n5584), .ZN(n10930) );
  INV_X1 U4753 ( .A(n10930), .ZN(n10931) );
  BUF_X1 U4754 ( .A(n10935), .Z(n10932) );
  INV_X1 U4755 ( .A(matrix_mul_2D_1__2__5_), .ZN(n10933) );
  INV_X1 U4756 ( .A(n5585), .ZN(n10934) );
  INV_X1 U4757 ( .A(n10934), .ZN(n10935) );
  BUF_X1 U4758 ( .A(n10939), .Z(n10936) );
  INV_X1 U4759 ( .A(matrix_mul_2D_1__2__4_), .ZN(n10937) );
  INV_X1 U4760 ( .A(n55860), .ZN(n10938) );
  INV_X1 U4761 ( .A(n10938), .ZN(n10939) );
  BUF_X1 U4762 ( .A(n10943), .Z(n10940) );
  INV_X1 U4763 ( .A(matrix_mul_2D_1__2__3_), .ZN(n10941) );
  INV_X1 U4764 ( .A(n55870), .ZN(n10942) );
  INV_X1 U4765 ( .A(n10942), .ZN(n10943) );
  BUF_X1 U4766 ( .A(n10947), .Z(n10944) );
  INV_X1 U4767 ( .A(matrix_mul_2D_1__2__2_), .ZN(n10945) );
  INV_X1 U4768 ( .A(n55880), .ZN(n10946) );
  INV_X1 U4769 ( .A(n10946), .ZN(n10947) );
  BUF_X1 U4770 ( .A(n10951), .Z(n10948) );
  INV_X1 U4771 ( .A(matrix_mul_2D_1__2__1_), .ZN(n10949) );
  INV_X1 U4772 ( .A(n55890), .ZN(n10950) );
  INV_X1 U4773 ( .A(n10950), .ZN(n10951) );
  BUF_X1 U4774 ( .A(n10956), .Z(n10952) );
  INV_X1 U4775 ( .A(n2021), .ZN(n10953) );
  INV_X1 U4776 ( .A(n10953), .ZN(n10954) );
  INV_X1 U4777 ( .A(n55900), .ZN(n10955) );
  INV_X1 U4778 ( .A(n10955), .ZN(n10956) );
  BUF_X1 U4779 ( .A(n27396), .Z(n10957) );
  BUF_X1 U4780 ( .A(n27397), .Z(n10958) );
  BUF_X1 U4781 ( .A(n27398), .Z(n10959) );
  BUF_X1 U4782 ( .A(n27399), .Z(n10960) );
  BUF_X1 U4783 ( .A(n274001), .Z(n10961) );
  BUF_X1 U4784 ( .A(n27401), .Z(n10962) );
  BUF_X1 U4785 ( .A(n10967), .Z(n10963) );
  INV_X1 U4786 ( .A(n1986), .ZN(n10964) );
  INV_X1 U4787 ( .A(n10964), .ZN(n10965) );
  INV_X1 U4788 ( .A(n55610), .ZN(n10966) );
  INV_X1 U4789 ( .A(n10966), .ZN(n10967) );
  BUF_X1 U4790 ( .A(n10972), .Z(n10968) );
  INV_X1 U4791 ( .A(n1987), .ZN(n10969) );
  INV_X1 U4792 ( .A(n10969), .ZN(n10970) );
  INV_X1 U4793 ( .A(n55620), .ZN(n10971) );
  INV_X1 U4794 ( .A(n10971), .ZN(n10972) );
  BUF_X1 U4795 ( .A(n10977), .Z(n10973) );
  INV_X1 U4796 ( .A(n1988), .ZN(n10974) );
  INV_X1 U4797 ( .A(n10974), .ZN(n10975) );
  INV_X1 U4798 ( .A(n55630), .ZN(n10976) );
  INV_X1 U4799 ( .A(n10976), .ZN(n10977) );
  BUF_X1 U4800 ( .A(n10982), .Z(n10978) );
  INV_X1 U4801 ( .A(n1989), .ZN(n10979) );
  INV_X1 U4802 ( .A(n10979), .ZN(n10980) );
  INV_X1 U4803 ( .A(n55640), .ZN(n10981) );
  INV_X1 U4804 ( .A(n10981), .ZN(n10982) );
  BUF_X1 U4805 ( .A(n10987), .Z(n10983) );
  INV_X1 U4806 ( .A(n1990), .ZN(n10984) );
  INV_X1 U4807 ( .A(n10984), .ZN(n10985) );
  INV_X1 U4808 ( .A(n55650), .ZN(n10986) );
  INV_X1 U4809 ( .A(n10986), .ZN(n10987) );
  BUF_X1 U4810 ( .A(n10992), .Z(n10988) );
  INV_X1 U4811 ( .A(n1991), .ZN(n10989) );
  INV_X1 U4812 ( .A(n10989), .ZN(n10990) );
  INV_X1 U4813 ( .A(n55660), .ZN(n10991) );
  INV_X1 U4814 ( .A(n10991), .ZN(n10992) );
  BUF_X1 U4815 ( .A(n10997), .Z(n10993) );
  INV_X1 U4816 ( .A(n1992), .ZN(n10994) );
  INV_X1 U4817 ( .A(n10994), .ZN(n10995) );
  INV_X1 U4818 ( .A(n55670), .ZN(n10996) );
  INV_X1 U4819 ( .A(n10996), .ZN(n10997) );
  BUF_X1 U4820 ( .A(n11002), .Z(n10998) );
  INV_X1 U4821 ( .A(n1993), .ZN(n10999) );
  INV_X1 U4822 ( .A(n10999), .ZN(n11000) );
  INV_X1 U4823 ( .A(n55680), .ZN(n11001) );
  INV_X1 U4824 ( .A(n11001), .ZN(n11002) );
  BUF_X1 U4825 ( .A(n11007), .Z(n11003) );
  INV_X1 U4826 ( .A(n1994), .ZN(n11004) );
  INV_X1 U4827 ( .A(n11004), .ZN(n11005) );
  INV_X1 U4828 ( .A(n5569), .ZN(n11006) );
  INV_X1 U4829 ( .A(n11006), .ZN(n11007) );
  BUF_X1 U4830 ( .A(n11012), .Z(n11008) );
  INV_X1 U4831 ( .A(n1995), .ZN(n11009) );
  INV_X1 U4832 ( .A(n11009), .ZN(n11010) );
  INV_X1 U4833 ( .A(n5570), .ZN(n11011) );
  INV_X1 U4834 ( .A(n11011), .ZN(n11012) );
  BUF_X1 U4835 ( .A(n11017), .Z(n11013) );
  INV_X1 U4836 ( .A(n1996), .ZN(n11014) );
  INV_X1 U4837 ( .A(n11014), .ZN(n11015) );
  INV_X1 U4838 ( .A(n5571), .ZN(n11016) );
  INV_X1 U4839 ( .A(n11016), .ZN(n11017) );
  BUF_X1 U4840 ( .A(n11022), .Z(n11018) );
  INV_X1 U4841 ( .A(n1997), .ZN(n11019) );
  INV_X1 U4842 ( .A(n11019), .ZN(n11020) );
  INV_X1 U4843 ( .A(n5572), .ZN(n11021) );
  INV_X1 U4844 ( .A(n11021), .ZN(n11022) );
  BUF_X1 U4845 ( .A(n11027), .Z(n11023) );
  INV_X1 U4846 ( .A(n1998), .ZN(n11024) );
  INV_X1 U4847 ( .A(n11024), .ZN(n11025) );
  INV_X1 U4848 ( .A(n5573), .ZN(n11026) );
  INV_X1 U4849 ( .A(n11026), .ZN(n11027) );
  BUF_X1 U4850 ( .A(n11032), .Z(n11028) );
  INV_X1 U4851 ( .A(n1999), .ZN(n11029) );
  INV_X1 U4852 ( .A(n11029), .ZN(n11030) );
  INV_X1 U4853 ( .A(n5574), .ZN(n11031) );
  INV_X1 U4854 ( .A(n11031), .ZN(n11032) );
  BUF_X1 U4855 ( .A(n11036), .Z(n11033) );
  INV_X1 U4856 ( .A(matrix_mul_2D_1__1__0_), .ZN(n11034) );
  INV_X1 U4857 ( .A(n5575), .ZN(n11035) );
  INV_X1 U4858 ( .A(n11035), .ZN(n11036) );
  BUF_X1 U4859 ( .A(n273901), .Z(n11037) );
  BUF_X1 U4860 ( .A(n27391), .Z(n11038) );
  BUF_X1 U4861 ( .A(n27392), .Z(n11039) );
  BUF_X1 U4862 ( .A(n27393), .Z(n11040) );
  BUF_X1 U4863 ( .A(n27394), .Z(n11041) );
  BUF_X1 U4864 ( .A(n27395), .Z(n11042) );
  BUF_X1 U4865 ( .A(n11047), .Z(n11043) );
  INV_X1 U4866 ( .A(n1971), .ZN(n11044) );
  INV_X1 U4867 ( .A(n11044), .ZN(n11045) );
  INV_X1 U4868 ( .A(n5546), .ZN(n11046) );
  INV_X1 U4869 ( .A(n11046), .ZN(n11047) );
  BUF_X1 U4870 ( .A(n11052), .Z(n11048) );
  INV_X1 U4871 ( .A(n1972), .ZN(n11049) );
  INV_X1 U4872 ( .A(n11049), .ZN(n11050) );
  INV_X1 U4873 ( .A(n5547), .ZN(n11051) );
  INV_X1 U4874 ( .A(n11051), .ZN(n11052) );
  BUF_X1 U4875 ( .A(n11057), .Z(n11053) );
  INV_X1 U4876 ( .A(n1973), .ZN(n11054) );
  INV_X1 U4877 ( .A(n11054), .ZN(n11055) );
  INV_X1 U4878 ( .A(n5548), .ZN(n11056) );
  INV_X1 U4879 ( .A(n11056), .ZN(n11057) );
  BUF_X1 U4880 ( .A(n11062), .Z(n11058) );
  INV_X1 U4881 ( .A(n1974), .ZN(n11059) );
  INV_X1 U4882 ( .A(n11059), .ZN(n11060) );
  INV_X1 U4883 ( .A(n5549), .ZN(n11061) );
  INV_X1 U4884 ( .A(n11061), .ZN(n11062) );
  BUF_X1 U4885 ( .A(n11067), .Z(n11063) );
  INV_X1 U4886 ( .A(n1975), .ZN(n11064) );
  INV_X1 U4887 ( .A(n11064), .ZN(n11065) );
  INV_X1 U4888 ( .A(n5550), .ZN(n11066) );
  INV_X1 U4889 ( .A(n11066), .ZN(n11067) );
  BUF_X1 U4890 ( .A(n11072), .Z(n11068) );
  INV_X1 U4891 ( .A(n1976), .ZN(n11069) );
  INV_X1 U4892 ( .A(n11069), .ZN(n11070) );
  INV_X1 U4893 ( .A(n5551), .ZN(n11071) );
  INV_X1 U4894 ( .A(n11071), .ZN(n11072) );
  BUF_X1 U4895 ( .A(n11077), .Z(n11073) );
  INV_X1 U4896 ( .A(n1977), .ZN(n11074) );
  INV_X1 U4897 ( .A(n11074), .ZN(n11075) );
  INV_X1 U4898 ( .A(n5552), .ZN(n11076) );
  INV_X1 U4899 ( .A(n11076), .ZN(n11077) );
  BUF_X1 U4900 ( .A(n11082), .Z(n11078) );
  INV_X1 U4901 ( .A(n1978), .ZN(n11079) );
  INV_X1 U4902 ( .A(n11079), .ZN(n11080) );
  INV_X1 U4903 ( .A(n55530), .ZN(n11081) );
  INV_X1 U4904 ( .A(n11081), .ZN(n11082) );
  BUF_X1 U4905 ( .A(n11087), .Z(n11083) );
  INV_X1 U4906 ( .A(n1979), .ZN(n11084) );
  INV_X1 U4907 ( .A(n11084), .ZN(n11085) );
  INV_X1 U4908 ( .A(n55540), .ZN(n11086) );
  INV_X1 U4909 ( .A(n11086), .ZN(n11087) );
  BUF_X1 U4910 ( .A(n11092), .Z(n11088) );
  INV_X1 U4911 ( .A(n1980), .ZN(n11089) );
  INV_X1 U4912 ( .A(n11089), .ZN(n11090) );
  INV_X1 U4913 ( .A(n55550), .ZN(n11091) );
  INV_X1 U4914 ( .A(n11091), .ZN(n11092) );
  BUF_X1 U4915 ( .A(n11097), .Z(n11093) );
  INV_X1 U4916 ( .A(n1981), .ZN(n11094) );
  INV_X1 U4917 ( .A(n11094), .ZN(n11095) );
  INV_X1 U4918 ( .A(n55560), .ZN(n11096) );
  INV_X1 U4919 ( .A(n11096), .ZN(n11097) );
  BUF_X1 U4920 ( .A(n11102), .Z(n11098) );
  INV_X1 U4921 ( .A(n1982), .ZN(n11099) );
  INV_X1 U4922 ( .A(n11099), .ZN(n11100) );
  INV_X1 U4923 ( .A(n55570), .ZN(n11101) );
  INV_X1 U4924 ( .A(n11101), .ZN(n11102) );
  BUF_X1 U4925 ( .A(n11107), .Z(n11103) );
  INV_X1 U4926 ( .A(n1983), .ZN(n11104) );
  INV_X1 U4927 ( .A(n11104), .ZN(n11105) );
  INV_X1 U4928 ( .A(n55580), .ZN(n11106) );
  INV_X1 U4929 ( .A(n11106), .ZN(n11107) );
  BUF_X1 U4930 ( .A(n11112), .Z(n11108) );
  INV_X1 U4931 ( .A(n1984), .ZN(n11109) );
  INV_X1 U4932 ( .A(n11109), .ZN(n11110) );
  INV_X1 U4933 ( .A(n55590), .ZN(n11111) );
  INV_X1 U4934 ( .A(n11111), .ZN(n11112) );
  BUF_X1 U4935 ( .A(n11116), .Z(n11113) );
  INV_X1 U4936 ( .A(matrix_mul_2D_1__0__0_), .ZN(n11114) );
  INV_X1 U4937 ( .A(n55600), .ZN(n11115) );
  INV_X1 U4938 ( .A(n11115), .ZN(n11116) );
  BUF_X1 U4939 ( .A(n27384), .Z(n11117) );
  BUF_X1 U4940 ( .A(n27385), .Z(n11118) );
  BUF_X1 U4941 ( .A(n27386), .Z(n11119) );
  BUF_X1 U4942 ( .A(n27387), .Z(n11120) );
  BUF_X1 U4943 ( .A(n27388), .Z(n11121) );
  BUF_X1 U4944 ( .A(n27389), .Z(n11122) );
  BUF_X1 U4945 ( .A(n11126), .Z(n11123) );
  INV_X1 U4946 ( .A(matrix_mul_2D_0__7__14_), .ZN(n11124) );
  INV_X1 U4947 ( .A(n5531), .ZN(n11125) );
  INV_X1 U4948 ( .A(n11125), .ZN(n11126) );
  BUF_X1 U4949 ( .A(n11130), .Z(n11127) );
  INV_X1 U4950 ( .A(matrix_mul_2D_0__7__13_), .ZN(n11128) );
  INV_X1 U4951 ( .A(n5532), .ZN(n11129) );
  INV_X1 U4952 ( .A(n11129), .ZN(n11130) );
  BUF_X1 U4953 ( .A(n11134), .Z(n11131) );
  INV_X1 U4954 ( .A(matrix_mul_2D_0__7__12_), .ZN(n11132) );
  INV_X1 U4955 ( .A(n5533), .ZN(n11133) );
  INV_X1 U4956 ( .A(n11133), .ZN(n11134) );
  BUF_X1 U4957 ( .A(n11138), .Z(n11135) );
  INV_X1 U4958 ( .A(matrix_mul_2D_0__7__11_), .ZN(n11136) );
  INV_X1 U4959 ( .A(n5534), .ZN(n11137) );
  INV_X1 U4960 ( .A(n11137), .ZN(n11138) );
  BUF_X1 U4961 ( .A(n11142), .Z(n11139) );
  INV_X1 U4962 ( .A(matrix_mul_2D_0__7__10_), .ZN(n11140) );
  INV_X1 U4963 ( .A(n5535), .ZN(n11141) );
  INV_X1 U4964 ( .A(n11141), .ZN(n11142) );
  BUF_X1 U4965 ( .A(n11146), .Z(n11143) );
  INV_X1 U4966 ( .A(matrix_mul_2D_0__7__9_), .ZN(n11144) );
  INV_X1 U4967 ( .A(n5536), .ZN(n11145) );
  INV_X1 U4968 ( .A(n11145), .ZN(n11146) );
  BUF_X1 U4969 ( .A(n11150), .Z(n11147) );
  INV_X1 U4970 ( .A(matrix_mul_2D_0__7__8_), .ZN(n11148) );
  INV_X1 U4971 ( .A(n5537), .ZN(n11149) );
  INV_X1 U4972 ( .A(n11149), .ZN(n11150) );
  BUF_X1 U4973 ( .A(n11154), .Z(n11151) );
  INV_X1 U4974 ( .A(matrix_mul_2D_0__7__7_), .ZN(n11152) );
  INV_X1 U4975 ( .A(n5538), .ZN(n11153) );
  INV_X1 U4976 ( .A(n11153), .ZN(n11154) );
  BUF_X1 U4977 ( .A(n11158), .Z(n11155) );
  INV_X1 U4978 ( .A(matrix_mul_2D_0__7__6_), .ZN(n11156) );
  INV_X1 U4979 ( .A(n5539), .ZN(n11157) );
  INV_X1 U4980 ( .A(n11157), .ZN(n11158) );
  BUF_X1 U4981 ( .A(n11162), .Z(n11159) );
  INV_X1 U4982 ( .A(matrix_mul_2D_0__7__5_), .ZN(n11160) );
  INV_X1 U4983 ( .A(n5540), .ZN(n11161) );
  INV_X1 U4984 ( .A(n11161), .ZN(n11162) );
  BUF_X1 U4985 ( .A(n11166), .Z(n11163) );
  INV_X1 U4986 ( .A(matrix_mul_2D_0__7__4_), .ZN(n11164) );
  INV_X1 U4987 ( .A(n5541), .ZN(n11165) );
  INV_X1 U4988 ( .A(n11165), .ZN(n11166) );
  BUF_X1 U4989 ( .A(n11170), .Z(n11167) );
  INV_X1 U4990 ( .A(matrix_mul_2D_0__7__3_), .ZN(n11168) );
  INV_X1 U4991 ( .A(n5542), .ZN(n11169) );
  INV_X1 U4992 ( .A(n11169), .ZN(n11170) );
  BUF_X1 U4993 ( .A(n11174), .Z(n11171) );
  INV_X1 U4994 ( .A(matrix_mul_2D_0__7__2_), .ZN(n11172) );
  INV_X1 U4995 ( .A(n5543), .ZN(n11173) );
  INV_X1 U4996 ( .A(n11173), .ZN(n11174) );
  BUF_X1 U4997 ( .A(n11178), .Z(n11175) );
  INV_X1 U4998 ( .A(matrix_mul_2D_0__7__1_), .ZN(n11176) );
  INV_X1 U4999 ( .A(n5544), .ZN(n11177) );
  INV_X1 U5000 ( .A(n11177), .ZN(n11178) );
  BUF_X1 U5001 ( .A(n11183), .Z(n11179) );
  INV_X1 U5002 ( .A(n1970), .ZN(n11180) );
  INV_X1 U5003 ( .A(n11180), .ZN(n11181) );
  INV_X1 U5004 ( .A(n5545), .ZN(n11182) );
  INV_X1 U5005 ( .A(n11182), .ZN(n11183) );
  BUF_X1 U5006 ( .A(n27378), .Z(n11184) );
  BUF_X1 U5007 ( .A(n27379), .Z(n11185) );
  BUF_X1 U5008 ( .A(n273801), .Z(n11186) );
  BUF_X1 U5009 ( .A(n27381), .Z(n11187) );
  BUF_X1 U5010 ( .A(n27382), .Z(n11188) );
  BUF_X1 U5011 ( .A(n27383), .Z(n11189) );
  BUF_X1 U5012 ( .A(n11194), .Z(n11190) );
  INV_X1 U5013 ( .A(n1941), .ZN(n11191) );
  INV_X1 U5014 ( .A(n11191), .ZN(n11192) );
  INV_X1 U5015 ( .A(n55160), .ZN(n11193) );
  INV_X1 U5016 ( .A(n11193), .ZN(n11194) );
  BUF_X1 U5017 ( .A(n11199), .Z(n11195) );
  INV_X1 U5018 ( .A(n1942), .ZN(n11196) );
  INV_X1 U5019 ( .A(n11196), .ZN(n11197) );
  INV_X1 U5020 ( .A(n55170), .ZN(n11198) );
  INV_X1 U5021 ( .A(n11198), .ZN(n11199) );
  BUF_X1 U5022 ( .A(n11204), .Z(n11200) );
  INV_X1 U5023 ( .A(n1943), .ZN(n11201) );
  INV_X1 U5024 ( .A(n11201), .ZN(n11202) );
  INV_X1 U5025 ( .A(n55180), .ZN(n11203) );
  INV_X1 U5026 ( .A(n11203), .ZN(n11204) );
  BUF_X1 U5027 ( .A(n11209), .Z(n11205) );
  INV_X1 U5028 ( .A(n1944), .ZN(n11206) );
  INV_X1 U5029 ( .A(n11206), .ZN(n11207) );
  INV_X1 U5030 ( .A(n55190), .ZN(n11208) );
  INV_X1 U5031 ( .A(n11208), .ZN(n11209) );
  BUF_X1 U5032 ( .A(n11214), .Z(n11210) );
  INV_X1 U5033 ( .A(n1945), .ZN(n11211) );
  INV_X1 U5034 ( .A(n11211), .ZN(n11212) );
  INV_X1 U5035 ( .A(n55200), .ZN(n11213) );
  INV_X1 U5036 ( .A(n11213), .ZN(n11214) );
  BUF_X1 U5037 ( .A(n11219), .Z(n11215) );
  INV_X1 U5038 ( .A(n1946), .ZN(n11216) );
  INV_X1 U5039 ( .A(n11216), .ZN(n11217) );
  INV_X1 U5040 ( .A(n55210), .ZN(n11218) );
  INV_X1 U5041 ( .A(n11218), .ZN(n11219) );
  BUF_X1 U5042 ( .A(n11224), .Z(n11220) );
  INV_X1 U5043 ( .A(n1947), .ZN(n11221) );
  INV_X1 U5044 ( .A(n11221), .ZN(n11222) );
  INV_X1 U5045 ( .A(n55220), .ZN(n11223) );
  INV_X1 U5046 ( .A(n11223), .ZN(n11224) );
  BUF_X1 U5047 ( .A(n11229), .Z(n11225) );
  INV_X1 U5048 ( .A(n1948), .ZN(n11226) );
  INV_X1 U5049 ( .A(n11226), .ZN(n11227) );
  INV_X1 U5050 ( .A(n55230), .ZN(n11228) );
  INV_X1 U5051 ( .A(n11228), .ZN(n11229) );
  BUF_X1 U5052 ( .A(n11234), .Z(n11230) );
  INV_X1 U5053 ( .A(n1949), .ZN(n11231) );
  INV_X1 U5054 ( .A(n11231), .ZN(n11232) );
  INV_X1 U5055 ( .A(n55240), .ZN(n11233) );
  INV_X1 U5056 ( .A(n11233), .ZN(n11234) );
  BUF_X1 U5057 ( .A(n11239), .Z(n11235) );
  INV_X1 U5058 ( .A(n1950), .ZN(n11236) );
  INV_X1 U5059 ( .A(n11236), .ZN(n11237) );
  INV_X1 U5060 ( .A(n55250), .ZN(n11238) );
  INV_X1 U5061 ( .A(n11238), .ZN(n11239) );
  BUF_X1 U5062 ( .A(n11244), .Z(n11240) );
  INV_X1 U5063 ( .A(n1951), .ZN(n11241) );
  INV_X1 U5064 ( .A(n11241), .ZN(n11242) );
  INV_X1 U5065 ( .A(n55260), .ZN(n11243) );
  INV_X1 U5066 ( .A(n11243), .ZN(n11244) );
  BUF_X1 U5067 ( .A(n11249), .Z(n11245) );
  INV_X1 U5068 ( .A(n1952), .ZN(n11246) );
  INV_X1 U5069 ( .A(n11246), .ZN(n11247) );
  INV_X1 U5070 ( .A(n55270), .ZN(n11248) );
  INV_X1 U5071 ( .A(n11248), .ZN(n11249) );
  BUF_X1 U5072 ( .A(n11254), .Z(n11250) );
  INV_X1 U5073 ( .A(n1953), .ZN(n11251) );
  INV_X1 U5074 ( .A(n11251), .ZN(n11252) );
  INV_X1 U5075 ( .A(n5528), .ZN(n11253) );
  INV_X1 U5076 ( .A(n11253), .ZN(n11254) );
  BUF_X1 U5077 ( .A(n11259), .Z(n11255) );
  INV_X1 U5078 ( .A(n1954), .ZN(n11256) );
  INV_X1 U5079 ( .A(n11256), .ZN(n11257) );
  INV_X1 U5080 ( .A(n5529), .ZN(n11258) );
  INV_X1 U5081 ( .A(n11258), .ZN(n11259) );
  BUF_X1 U5082 ( .A(n11263), .Z(n11260) );
  INV_X1 U5083 ( .A(matrix_mul_2D_0__6__0_), .ZN(n11261) );
  INV_X1 U5084 ( .A(n5530), .ZN(n11262) );
  INV_X1 U5085 ( .A(n11262), .ZN(n11263) );
  BUF_X1 U5086 ( .A(n27372), .Z(n11264) );
  BUF_X1 U5087 ( .A(n27373), .Z(n11265) );
  BUF_X1 U5088 ( .A(n27374), .Z(n11266) );
  BUF_X1 U5089 ( .A(n27375), .Z(n11267) );
  BUF_X1 U5090 ( .A(n27376), .Z(n11268) );
  BUF_X1 U5091 ( .A(n27377), .Z(n11269) );
  BUF_X1 U5092 ( .A(n11273), .Z(n11270) );
  INV_X1 U5093 ( .A(matrix_mul_2D_0__5__14_), .ZN(n11271) );
  INV_X1 U5094 ( .A(n5501), .ZN(n11272) );
  INV_X1 U5095 ( .A(n11272), .ZN(n11273) );
  BUF_X1 U5096 ( .A(n11277), .Z(n11274) );
  INV_X1 U5097 ( .A(matrix_mul_2D_0__5__13_), .ZN(n11275) );
  INV_X1 U5098 ( .A(n5502), .ZN(n11276) );
  INV_X1 U5099 ( .A(n11276), .ZN(n11277) );
  BUF_X1 U5100 ( .A(n11281), .Z(n11278) );
  INV_X1 U5101 ( .A(matrix_mul_2D_0__5__12_), .ZN(n11279) );
  INV_X1 U5102 ( .A(n5503), .ZN(n11280) );
  INV_X1 U5103 ( .A(n11280), .ZN(n11281) );
  BUF_X1 U5104 ( .A(n11285), .Z(n11282) );
  INV_X1 U5105 ( .A(matrix_mul_2D_0__5__11_), .ZN(n11283) );
  INV_X1 U5106 ( .A(n5504), .ZN(n11284) );
  INV_X1 U5107 ( .A(n11284), .ZN(n11285) );
  BUF_X1 U5108 ( .A(n11289), .Z(n11286) );
  INV_X1 U5109 ( .A(matrix_mul_2D_0__5__10_), .ZN(n11287) );
  INV_X1 U5110 ( .A(n5505), .ZN(n11288) );
  INV_X1 U5111 ( .A(n11288), .ZN(n11289) );
  BUF_X1 U5112 ( .A(n11293), .Z(n11290) );
  INV_X1 U5113 ( .A(matrix_mul_2D_0__5__9_), .ZN(n11291) );
  INV_X1 U5114 ( .A(n5506), .ZN(n11292) );
  INV_X1 U5115 ( .A(n11292), .ZN(n11293) );
  BUF_X1 U5116 ( .A(n11297), .Z(n11294) );
  INV_X1 U5117 ( .A(matrix_mul_2D_0__5__8_), .ZN(n11295) );
  INV_X1 U5118 ( .A(n55070), .ZN(n11296) );
  INV_X1 U5119 ( .A(n11296), .ZN(n11297) );
  BUF_X1 U5120 ( .A(n11301), .Z(n11298) );
  INV_X1 U5121 ( .A(matrix_mul_2D_0__5__7_), .ZN(n11299) );
  INV_X1 U5122 ( .A(n55080), .ZN(n11300) );
  INV_X1 U5123 ( .A(n11300), .ZN(n11301) );
  BUF_X1 U5124 ( .A(n11305), .Z(n11302) );
  INV_X1 U5125 ( .A(matrix_mul_2D_0__5__6_), .ZN(n11303) );
  INV_X1 U5126 ( .A(n55090), .ZN(n11304) );
  INV_X1 U5127 ( .A(n11304), .ZN(n11305) );
  BUF_X1 U5128 ( .A(n11309), .Z(n11306) );
  INV_X1 U5129 ( .A(matrix_mul_2D_0__5__5_), .ZN(n11307) );
  INV_X1 U5130 ( .A(n55100), .ZN(n11308) );
  INV_X1 U5131 ( .A(n11308), .ZN(n11309) );
  BUF_X1 U5132 ( .A(n11313), .Z(n11310) );
  INV_X1 U5133 ( .A(matrix_mul_2D_0__5__4_), .ZN(n11311) );
  INV_X1 U5134 ( .A(n55110), .ZN(n11312) );
  INV_X1 U5135 ( .A(n11312), .ZN(n11313) );
  BUF_X1 U5136 ( .A(n11317), .Z(n11314) );
  INV_X1 U5137 ( .A(matrix_mul_2D_0__5__3_), .ZN(n11315) );
  INV_X1 U5138 ( .A(n55120), .ZN(n11316) );
  INV_X1 U5139 ( .A(n11316), .ZN(n11317) );
  BUF_X1 U5140 ( .A(n11321), .Z(n11318) );
  INV_X1 U5141 ( .A(matrix_mul_2D_0__5__2_), .ZN(n11319) );
  INV_X1 U5142 ( .A(n55130), .ZN(n11320) );
  INV_X1 U5143 ( .A(n11320), .ZN(n11321) );
  BUF_X1 U5144 ( .A(n11325), .Z(n11322) );
  INV_X1 U5145 ( .A(matrix_mul_2D_0__5__1_), .ZN(n11323) );
  INV_X1 U5146 ( .A(n55140), .ZN(n11324) );
  INV_X1 U5147 ( .A(n11324), .ZN(n11325) );
  BUF_X1 U5148 ( .A(n11330), .Z(n11326) );
  INV_X1 U5149 ( .A(n1940), .ZN(n11327) );
  INV_X1 U5150 ( .A(n11327), .ZN(n11328) );
  INV_X1 U5151 ( .A(n55150), .ZN(n11329) );
  INV_X1 U5152 ( .A(n11329), .ZN(n11330) );
  BUF_X1 U5153 ( .A(n27366), .Z(n11331) );
  BUF_X1 U5154 ( .A(n27367), .Z(n11332) );
  BUF_X1 U5155 ( .A(n27368), .Z(n11333) );
  BUF_X1 U5156 ( .A(n27369), .Z(n11334) );
  BUF_X1 U5157 ( .A(n273701), .Z(n11335) );
  BUF_X1 U5158 ( .A(n27371), .Z(n11336) );
  BUF_X1 U5159 ( .A(n11341), .Z(n11337) );
  INV_X1 U5160 ( .A(n1905), .ZN(n11338) );
  INV_X1 U5161 ( .A(n11338), .ZN(n11339) );
  INV_X1 U5162 ( .A(n54860), .ZN(n11340) );
  INV_X1 U5163 ( .A(n11340), .ZN(n11341) );
  BUF_X1 U5164 ( .A(n11346), .Z(n11342) );
  INV_X1 U5165 ( .A(n1906), .ZN(n11343) );
  INV_X1 U5166 ( .A(n11343), .ZN(n11344) );
  INV_X1 U5167 ( .A(n54870), .ZN(n11345) );
  INV_X1 U5168 ( .A(n11345), .ZN(n11346) );
  BUF_X1 U5169 ( .A(n11351), .Z(n11347) );
  INV_X1 U5170 ( .A(n1907), .ZN(n11348) );
  INV_X1 U5171 ( .A(n11348), .ZN(n11349) );
  INV_X1 U5172 ( .A(n54880), .ZN(n11350) );
  INV_X1 U5173 ( .A(n11350), .ZN(n11351) );
  BUF_X1 U5174 ( .A(n11356), .Z(n11352) );
  INV_X1 U5175 ( .A(n1908), .ZN(n11353) );
  INV_X1 U5176 ( .A(n11353), .ZN(n11354) );
  INV_X1 U5177 ( .A(n54890), .ZN(n11355) );
  INV_X1 U5178 ( .A(n11355), .ZN(n11356) );
  BUF_X1 U5179 ( .A(n11361), .Z(n11357) );
  INV_X1 U5180 ( .A(n1909), .ZN(n11358) );
  INV_X1 U5181 ( .A(n11358), .ZN(n11359) );
  INV_X1 U5182 ( .A(n5490), .ZN(n11360) );
  INV_X1 U5183 ( .A(n11360), .ZN(n11361) );
  BUF_X1 U5184 ( .A(n11366), .Z(n11362) );
  INV_X1 U5185 ( .A(n1910), .ZN(n11363) );
  INV_X1 U5186 ( .A(n11363), .ZN(n11364) );
  INV_X1 U5187 ( .A(n5491), .ZN(n11365) );
  INV_X1 U5188 ( .A(n11365), .ZN(n11366) );
  BUF_X1 U5189 ( .A(n11371), .Z(n11367) );
  INV_X1 U5190 ( .A(n1911), .ZN(n11368) );
  INV_X1 U5191 ( .A(n11368), .ZN(n11369) );
  INV_X1 U5192 ( .A(n5492), .ZN(n11370) );
  INV_X1 U5193 ( .A(n11370), .ZN(n11371) );
  BUF_X1 U5194 ( .A(n11376), .Z(n11372) );
  INV_X1 U5195 ( .A(n1912), .ZN(n11373) );
  INV_X1 U5196 ( .A(n11373), .ZN(n11374) );
  INV_X1 U5197 ( .A(n5493), .ZN(n11375) );
  INV_X1 U5198 ( .A(n11375), .ZN(n11376) );
  BUF_X1 U5199 ( .A(n11381), .Z(n11377) );
  INV_X1 U5200 ( .A(n1913), .ZN(n11378) );
  INV_X1 U5201 ( .A(n11378), .ZN(n11379) );
  INV_X1 U5202 ( .A(n5494), .ZN(n11380) );
  INV_X1 U5203 ( .A(n11380), .ZN(n11381) );
  BUF_X1 U5204 ( .A(n11386), .Z(n11382) );
  INV_X1 U5205 ( .A(n1914), .ZN(n11383) );
  INV_X1 U5206 ( .A(n11383), .ZN(n11384) );
  INV_X1 U5207 ( .A(n5495), .ZN(n11385) );
  INV_X1 U5208 ( .A(n11385), .ZN(n11386) );
  BUF_X1 U5209 ( .A(n11391), .Z(n11387) );
  INV_X1 U5210 ( .A(n1915), .ZN(n11388) );
  INV_X1 U5211 ( .A(n11388), .ZN(n11389) );
  INV_X1 U5212 ( .A(n5496), .ZN(n11390) );
  INV_X1 U5213 ( .A(n11390), .ZN(n11391) );
  BUF_X1 U5214 ( .A(n11396), .Z(n11392) );
  INV_X1 U5215 ( .A(n1916), .ZN(n11393) );
  INV_X1 U5216 ( .A(n11393), .ZN(n11394) );
  INV_X1 U5217 ( .A(n5497), .ZN(n11395) );
  INV_X1 U5218 ( .A(n11395), .ZN(n11396) );
  BUF_X1 U5219 ( .A(n11401), .Z(n11397) );
  INV_X1 U5220 ( .A(n1917), .ZN(n11398) );
  INV_X1 U5221 ( .A(n11398), .ZN(n11399) );
  INV_X1 U5222 ( .A(n5498), .ZN(n11400) );
  INV_X1 U5223 ( .A(n11400), .ZN(n11401) );
  BUF_X1 U5224 ( .A(n11406), .Z(n11402) );
  INV_X1 U5225 ( .A(n1918), .ZN(n11403) );
  INV_X1 U5226 ( .A(n11403), .ZN(n11404) );
  INV_X1 U5227 ( .A(n5499), .ZN(n11405) );
  INV_X1 U5228 ( .A(n11405), .ZN(n11406) );
  BUF_X1 U5229 ( .A(n11410), .Z(n11407) );
  INV_X1 U5230 ( .A(matrix_mul_2D_0__4__0_), .ZN(n11408) );
  INV_X1 U5231 ( .A(n5500), .ZN(n11409) );
  INV_X1 U5232 ( .A(n11409), .ZN(n11410) );
  BUF_X1 U5233 ( .A(n273601), .Z(n11411) );
  BUF_X1 U5234 ( .A(n27361), .Z(n11412) );
  BUF_X1 U5235 ( .A(n27362), .Z(n11413) );
  BUF_X1 U5236 ( .A(n27363), .Z(n11414) );
  BUF_X1 U5237 ( .A(n27364), .Z(n11415) );
  BUF_X1 U5238 ( .A(n27365), .Z(n11416) );
  BUF_X1 U5239 ( .A(n11421), .Z(n11417) );
  INV_X1 U5240 ( .A(n1890), .ZN(n11418) );
  INV_X1 U5241 ( .A(n11418), .ZN(n11419) );
  INV_X1 U5242 ( .A(n5471), .ZN(n11420) );
  INV_X1 U5243 ( .A(n11420), .ZN(n11421) );
  BUF_X1 U5244 ( .A(n11426), .Z(n11422) );
  INV_X1 U5245 ( .A(n1891), .ZN(n11423) );
  INV_X1 U5246 ( .A(n11423), .ZN(n11424) );
  INV_X1 U5247 ( .A(n5472), .ZN(n11425) );
  INV_X1 U5248 ( .A(n11425), .ZN(n11426) );
  BUF_X1 U5249 ( .A(n11431), .Z(n11427) );
  INV_X1 U5250 ( .A(n1892), .ZN(n11428) );
  INV_X1 U5251 ( .A(n11428), .ZN(n11429) );
  INV_X1 U5252 ( .A(n5473), .ZN(n11430) );
  INV_X1 U5253 ( .A(n11430), .ZN(n11431) );
  BUF_X1 U5254 ( .A(n11436), .Z(n11432) );
  INV_X1 U5255 ( .A(n1893), .ZN(n11433) );
  INV_X1 U5256 ( .A(n11433), .ZN(n11434) );
  INV_X1 U5257 ( .A(n54740), .ZN(n11435) );
  INV_X1 U5258 ( .A(n11435), .ZN(n11436) );
  BUF_X1 U5259 ( .A(n11441), .Z(n11437) );
  INV_X1 U5260 ( .A(n1894), .ZN(n11438) );
  INV_X1 U5261 ( .A(n11438), .ZN(n11439) );
  INV_X1 U5262 ( .A(n54750), .ZN(n11440) );
  INV_X1 U5263 ( .A(n11440), .ZN(n11441) );
  BUF_X1 U5264 ( .A(n11446), .Z(n11442) );
  INV_X1 U5265 ( .A(n1895), .ZN(n11443) );
  INV_X1 U5266 ( .A(n11443), .ZN(n11444) );
  INV_X1 U5267 ( .A(n54760), .ZN(n11445) );
  INV_X1 U5268 ( .A(n11445), .ZN(n11446) );
  BUF_X1 U5269 ( .A(n11451), .Z(n11447) );
  INV_X1 U5270 ( .A(n1896), .ZN(n11448) );
  INV_X1 U5271 ( .A(n11448), .ZN(n11449) );
  INV_X1 U5272 ( .A(n54770), .ZN(n11450) );
  INV_X1 U5273 ( .A(n11450), .ZN(n11451) );
  BUF_X1 U5274 ( .A(n11456), .Z(n11452) );
  INV_X1 U5275 ( .A(n1897), .ZN(n11453) );
  INV_X1 U5276 ( .A(n11453), .ZN(n11454) );
  INV_X1 U5277 ( .A(n54780), .ZN(n11455) );
  INV_X1 U5278 ( .A(n11455), .ZN(n11456) );
  BUF_X1 U5279 ( .A(n11461), .Z(n11457) );
  INV_X1 U5280 ( .A(n1898), .ZN(n11458) );
  INV_X1 U5281 ( .A(n11458), .ZN(n11459) );
  INV_X1 U5282 ( .A(n54790), .ZN(n11460) );
  INV_X1 U5283 ( .A(n11460), .ZN(n11461) );
  BUF_X1 U5284 ( .A(n11466), .Z(n11462) );
  INV_X1 U5285 ( .A(n1899), .ZN(n11463) );
  INV_X1 U5286 ( .A(n11463), .ZN(n11464) );
  INV_X1 U5287 ( .A(n54800), .ZN(n11465) );
  INV_X1 U5288 ( .A(n11465), .ZN(n11466) );
  BUF_X1 U5289 ( .A(n11471), .Z(n11467) );
  INV_X1 U5290 ( .A(n1900), .ZN(n11468) );
  INV_X1 U5291 ( .A(n11468), .ZN(n11469) );
  INV_X1 U5292 ( .A(n54810), .ZN(n11470) );
  INV_X1 U5293 ( .A(n11470), .ZN(n11471) );
  BUF_X1 U5294 ( .A(n11476), .Z(n11472) );
  INV_X1 U5295 ( .A(n1901), .ZN(n11473) );
  INV_X1 U5296 ( .A(n11473), .ZN(n11474) );
  INV_X1 U5297 ( .A(n54820), .ZN(n11475) );
  INV_X1 U5298 ( .A(n11475), .ZN(n11476) );
  BUF_X1 U5299 ( .A(n11481), .Z(n11477) );
  INV_X1 U5300 ( .A(n1902), .ZN(n11478) );
  INV_X1 U5301 ( .A(n11478), .ZN(n11479) );
  INV_X1 U5302 ( .A(n54830), .ZN(n11480) );
  INV_X1 U5303 ( .A(n11480), .ZN(n11481) );
  BUF_X1 U5304 ( .A(n11486), .Z(n11482) );
  INV_X1 U5305 ( .A(n1903), .ZN(n11483) );
  INV_X1 U5306 ( .A(n11483), .ZN(n11484) );
  INV_X1 U5307 ( .A(n54840), .ZN(n11485) );
  INV_X1 U5308 ( .A(n11485), .ZN(n11486) );
  BUF_X1 U5309 ( .A(n11490), .Z(n11487) );
  INV_X1 U5310 ( .A(matrix_mul_2D_0__3__0_), .ZN(n11488) );
  INV_X1 U5311 ( .A(n54850), .ZN(n11489) );
  INV_X1 U5312 ( .A(n11489), .ZN(n11490) );
  BUF_X1 U5313 ( .A(n27354), .Z(n11491) );
  BUF_X1 U5314 ( .A(n27355), .Z(n11492) );
  BUF_X1 U5315 ( .A(n27356), .Z(n11493) );
  BUF_X1 U5316 ( .A(n27357), .Z(n11494) );
  BUF_X1 U5317 ( .A(n27358), .Z(n11495) );
  BUF_X1 U5318 ( .A(n27359), .Z(n11496) );
  BUF_X1 U5319 ( .A(n11501), .Z(n11497) );
  INV_X1 U5320 ( .A(n1875), .ZN(n11498) );
  INV_X1 U5321 ( .A(n11498), .ZN(n11499) );
  INV_X1 U5322 ( .A(n5456), .ZN(n11500) );
  INV_X1 U5323 ( .A(n11500), .ZN(n11501) );
  BUF_X1 U5324 ( .A(n11506), .Z(n11502) );
  INV_X1 U5325 ( .A(n1876), .ZN(n11503) );
  INV_X1 U5326 ( .A(n11503), .ZN(n11504) );
  INV_X1 U5327 ( .A(n5457), .ZN(n11505) );
  INV_X1 U5328 ( .A(n11505), .ZN(n11506) );
  BUF_X1 U5329 ( .A(n11511), .Z(n11507) );
  INV_X1 U5330 ( .A(n1877), .ZN(n11508) );
  INV_X1 U5331 ( .A(n11508), .ZN(n11509) );
  INV_X1 U5332 ( .A(n5458), .ZN(n11510) );
  INV_X1 U5333 ( .A(n11510), .ZN(n11511) );
  BUF_X1 U5334 ( .A(n11516), .Z(n11512) );
  INV_X1 U5335 ( .A(n1878), .ZN(n11513) );
  INV_X1 U5336 ( .A(n11513), .ZN(n11514) );
  INV_X1 U5337 ( .A(n5459), .ZN(n11515) );
  INV_X1 U5338 ( .A(n11515), .ZN(n11516) );
  BUF_X1 U5339 ( .A(n11521), .Z(n11517) );
  INV_X1 U5340 ( .A(n1879), .ZN(n11518) );
  INV_X1 U5341 ( .A(n11518), .ZN(n11519) );
  INV_X1 U5342 ( .A(n5460), .ZN(n11520) );
  INV_X1 U5343 ( .A(n11520), .ZN(n11521) );
  BUF_X1 U5344 ( .A(n11526), .Z(n11522) );
  INV_X1 U5345 ( .A(n1880), .ZN(n11523) );
  INV_X1 U5346 ( .A(n11523), .ZN(n11524) );
  INV_X1 U5347 ( .A(n5461), .ZN(n11525) );
  INV_X1 U5348 ( .A(n11525), .ZN(n11526) );
  BUF_X1 U5349 ( .A(n11531), .Z(n11527) );
  INV_X1 U5350 ( .A(n1881), .ZN(n11528) );
  INV_X1 U5351 ( .A(n11528), .ZN(n11529) );
  INV_X1 U5352 ( .A(n5462), .ZN(n11530) );
  INV_X1 U5353 ( .A(n11530), .ZN(n11531) );
  BUF_X1 U5354 ( .A(n11536), .Z(n11532) );
  INV_X1 U5355 ( .A(n1882), .ZN(n11533) );
  INV_X1 U5356 ( .A(n11533), .ZN(n11534) );
  INV_X1 U5357 ( .A(n5463), .ZN(n11535) );
  INV_X1 U5358 ( .A(n11535), .ZN(n11536) );
  BUF_X1 U5359 ( .A(n11541), .Z(n11537) );
  INV_X1 U5360 ( .A(n1883), .ZN(n11538) );
  INV_X1 U5361 ( .A(n11538), .ZN(n11539) );
  INV_X1 U5362 ( .A(n5464), .ZN(n11540) );
  INV_X1 U5363 ( .A(n11540), .ZN(n11541) );
  BUF_X1 U5364 ( .A(n11546), .Z(n11542) );
  INV_X1 U5365 ( .A(n1884), .ZN(n11543) );
  INV_X1 U5366 ( .A(n11543), .ZN(n11544) );
  INV_X1 U5367 ( .A(n5465), .ZN(n11545) );
  INV_X1 U5368 ( .A(n11545), .ZN(n11546) );
  BUF_X1 U5369 ( .A(n11551), .Z(n11547) );
  INV_X1 U5370 ( .A(n1885), .ZN(n11548) );
  INV_X1 U5371 ( .A(n11548), .ZN(n11549) );
  INV_X1 U5372 ( .A(n5466), .ZN(n11550) );
  INV_X1 U5373 ( .A(n11550), .ZN(n11551) );
  BUF_X1 U5374 ( .A(n11556), .Z(n11552) );
  INV_X1 U5375 ( .A(n1886), .ZN(n11553) );
  INV_X1 U5376 ( .A(n11553), .ZN(n11554) );
  INV_X1 U5377 ( .A(n5467), .ZN(n11555) );
  INV_X1 U5378 ( .A(n11555), .ZN(n11556) );
  BUF_X1 U5379 ( .A(n11561), .Z(n11557) );
  INV_X1 U5380 ( .A(n1887), .ZN(n11558) );
  INV_X1 U5381 ( .A(n11558), .ZN(n11559) );
  INV_X1 U5382 ( .A(n5468), .ZN(n11560) );
  INV_X1 U5383 ( .A(n11560), .ZN(n11561) );
  BUF_X1 U5384 ( .A(n11566), .Z(n11562) );
  INV_X1 U5385 ( .A(n1888), .ZN(n11563) );
  INV_X1 U5386 ( .A(n11563), .ZN(n11564) );
  INV_X1 U5387 ( .A(n5469), .ZN(n11565) );
  INV_X1 U5388 ( .A(n11565), .ZN(n11566) );
  BUF_X1 U5389 ( .A(n11570), .Z(n11567) );
  INV_X1 U5390 ( .A(matrix_mul_2D_0__2__0_), .ZN(n11568) );
  INV_X1 U5391 ( .A(n5470), .ZN(n11569) );
  INV_X1 U5392 ( .A(n11569), .ZN(n11570) );
  BUF_X1 U5393 ( .A(n27348), .Z(n11571) );
  BUF_X1 U5394 ( .A(n27349), .Z(n11572) );
  BUF_X1 U5395 ( .A(n273501), .Z(n11573) );
  BUF_X1 U5396 ( .A(n27351), .Z(n11574) );
  BUF_X1 U5397 ( .A(n27352), .Z(n11575) );
  BUF_X1 U5398 ( .A(n27353), .Z(n11576) );
  BUF_X1 U5399 ( .A(n11581), .Z(n11577) );
  INV_X1 U5400 ( .A(n1860), .ZN(n11578) );
  INV_X1 U5401 ( .A(n11578), .ZN(n11579) );
  INV_X1 U5402 ( .A(n5441), .ZN(n11580) );
  INV_X1 U5403 ( .A(n11580), .ZN(n11581) );
  BUF_X1 U5404 ( .A(n11586), .Z(n11582) );
  INV_X1 U5405 ( .A(n1861), .ZN(n11583) );
  INV_X1 U5406 ( .A(n11583), .ZN(n11584) );
  INV_X1 U5407 ( .A(n5442), .ZN(n11585) );
  INV_X1 U5408 ( .A(n11585), .ZN(n11586) );
  BUF_X1 U5409 ( .A(n11591), .Z(n11587) );
  INV_X1 U5410 ( .A(n1862), .ZN(n11588) );
  INV_X1 U5411 ( .A(n11588), .ZN(n11589) );
  INV_X1 U5412 ( .A(n5443), .ZN(n11590) );
  INV_X1 U5413 ( .A(n11590), .ZN(n11591) );
  BUF_X1 U5414 ( .A(n11596), .Z(n11592) );
  INV_X1 U5415 ( .A(n1863), .ZN(n11593) );
  INV_X1 U5416 ( .A(n11593), .ZN(n11594) );
  INV_X1 U5417 ( .A(n5444), .ZN(n11595) );
  INV_X1 U5418 ( .A(n11595), .ZN(n11596) );
  BUF_X1 U5419 ( .A(n11601), .Z(n11597) );
  INV_X1 U5420 ( .A(n1864), .ZN(n11598) );
  INV_X1 U5421 ( .A(n11598), .ZN(n11599) );
  INV_X1 U5422 ( .A(n5445), .ZN(n11600) );
  INV_X1 U5423 ( .A(n11600), .ZN(n11601) );
  BUF_X1 U5424 ( .A(n11606), .Z(n11602) );
  INV_X1 U5425 ( .A(n1865), .ZN(n11603) );
  INV_X1 U5426 ( .A(n11603), .ZN(n11604) );
  INV_X1 U5427 ( .A(n5446), .ZN(n11605) );
  INV_X1 U5428 ( .A(n11605), .ZN(n11606) );
  BUF_X1 U5429 ( .A(n11611), .Z(n11607) );
  INV_X1 U5430 ( .A(n1866), .ZN(n11608) );
  INV_X1 U5431 ( .A(n11608), .ZN(n11609) );
  INV_X1 U5432 ( .A(n5447), .ZN(n11610) );
  INV_X1 U5433 ( .A(n11610), .ZN(n11611) );
  BUF_X1 U5434 ( .A(n11616), .Z(n11612) );
  INV_X1 U5435 ( .A(n1867), .ZN(n11613) );
  INV_X1 U5436 ( .A(n11613), .ZN(n11614) );
  INV_X1 U5437 ( .A(n5448), .ZN(n11615) );
  INV_X1 U5438 ( .A(n11615), .ZN(n11616) );
  BUF_X1 U5439 ( .A(n11621), .Z(n11617) );
  INV_X1 U5440 ( .A(n1868), .ZN(n11618) );
  INV_X1 U5441 ( .A(n11618), .ZN(n11619) );
  INV_X1 U5442 ( .A(n5449), .ZN(n11620) );
  INV_X1 U5443 ( .A(n11620), .ZN(n11621) );
  BUF_X1 U5444 ( .A(n11626), .Z(n11622) );
  INV_X1 U5445 ( .A(n1869), .ZN(n11623) );
  INV_X1 U5446 ( .A(n11623), .ZN(n11624) );
  INV_X1 U5447 ( .A(n5450), .ZN(n11625) );
  INV_X1 U5448 ( .A(n11625), .ZN(n11626) );
  BUF_X1 U5449 ( .A(n11631), .Z(n11627) );
  INV_X1 U5450 ( .A(n1870), .ZN(n11628) );
  INV_X1 U5451 ( .A(n11628), .ZN(n11629) );
  INV_X1 U5452 ( .A(n5451), .ZN(n11630) );
  INV_X1 U5453 ( .A(n11630), .ZN(n11631) );
  BUF_X1 U5454 ( .A(n11636), .Z(n11632) );
  INV_X1 U5455 ( .A(n1871), .ZN(n11633) );
  INV_X1 U5456 ( .A(n11633), .ZN(n11634) );
  INV_X1 U5457 ( .A(n5452), .ZN(n11635) );
  INV_X1 U5458 ( .A(n11635), .ZN(n11636) );
  BUF_X1 U5459 ( .A(n11641), .Z(n11637) );
  INV_X1 U5460 ( .A(n1872), .ZN(n11638) );
  INV_X1 U5461 ( .A(n11638), .ZN(n11639) );
  INV_X1 U5462 ( .A(n5453), .ZN(n11640) );
  INV_X1 U5463 ( .A(n11640), .ZN(n11641) );
  BUF_X1 U5464 ( .A(n11646), .Z(n11642) );
  INV_X1 U5465 ( .A(n1873), .ZN(n11643) );
  INV_X1 U5466 ( .A(n11643), .ZN(n11644) );
  INV_X1 U5467 ( .A(n5454), .ZN(n11645) );
  INV_X1 U5468 ( .A(n11645), .ZN(n11646) );
  BUF_X1 U5469 ( .A(n11650), .Z(n11647) );
  INV_X1 U5470 ( .A(matrix_mul_2D_0__1__0_), .ZN(n11648) );
  INV_X1 U5471 ( .A(n5455), .ZN(n11649) );
  INV_X1 U5472 ( .A(n11649), .ZN(n11650) );
  BUF_X1 U5473 ( .A(n27342), .Z(n11651) );
  BUF_X1 U5474 ( .A(n27343), .Z(n11652) );
  BUF_X1 U5475 ( .A(n27344), .Z(n11653) );
  BUF_X1 U5476 ( .A(n27345), .Z(n11654) );
  BUF_X1 U5477 ( .A(n27346), .Z(n11655) );
  BUF_X1 U5478 ( .A(n27347), .Z(n11656) );
  INV_X1 U5479 ( .A(n1844), .ZN(n11854) );
  BUF_X1 U5480 ( .A(n11855), .Z(n11657) );
  INV_X1 U5481 ( .A(n6386), .ZN(n11658) );
  INV_X1 U5482 ( .A(n11658), .ZN(n11659) );
  INV_X1 U5483 ( .A(n1843), .ZN(n11861) );
  BUF_X1 U5484 ( .A(n11862), .Z(n11660) );
  INV_X1 U5485 ( .A(n6387), .ZN(n11661) );
  INV_X1 U5486 ( .A(n11661), .ZN(n11662) );
  INV_X1 U5487 ( .A(n1842), .ZN(n11868) );
  BUF_X1 U5488 ( .A(n11869), .Z(n11663) );
  INV_X1 U5489 ( .A(n6388), .ZN(n11664) );
  INV_X1 U5490 ( .A(n11664), .ZN(n11665) );
  INV_X1 U5491 ( .A(n1841), .ZN(n11875) );
  BUF_X1 U5492 ( .A(n11876), .Z(n11666) );
  INV_X1 U5493 ( .A(n6389), .ZN(n11667) );
  INV_X1 U5494 ( .A(n11667), .ZN(n11668) );
  INV_X1 U5495 ( .A(n1840), .ZN(n11882) );
  BUF_X1 U5496 ( .A(n11883), .Z(n11669) );
  INV_X1 U5497 ( .A(n6390), .ZN(n11670) );
  INV_X1 U5498 ( .A(n11670), .ZN(n11671) );
  INV_X1 U5499 ( .A(n1839), .ZN(n11889) );
  BUF_X1 U5500 ( .A(n11890), .Z(n11672) );
  INV_X1 U5501 ( .A(n6391), .ZN(n11673) );
  INV_X1 U5502 ( .A(n11673), .ZN(n11674) );
  INV_X1 U5503 ( .A(n1838), .ZN(n11896) );
  BUF_X1 U5504 ( .A(n11897), .Z(n11675) );
  INV_X1 U5505 ( .A(n6392), .ZN(n11676) );
  INV_X1 U5506 ( .A(n11676), .ZN(n11677) );
  INV_X1 U5507 ( .A(n1837), .ZN(n11903) );
  BUF_X1 U5508 ( .A(n11904), .Z(n11678) );
  INV_X1 U5509 ( .A(n6393), .ZN(n11679) );
  INV_X1 U5510 ( .A(n11679), .ZN(n11680) );
  INV_X1 U5511 ( .A(n1836), .ZN(n11910) );
  BUF_X1 U5512 ( .A(n11911), .Z(n11681) );
  INV_X1 U5513 ( .A(n6394), .ZN(n11682) );
  INV_X1 U5514 ( .A(n11682), .ZN(n11683) );
  INV_X1 U5515 ( .A(n1835), .ZN(n11917) );
  BUF_X1 U5516 ( .A(n11918), .Z(n11684) );
  INV_X1 U5517 ( .A(n6395), .ZN(n11685) );
  INV_X1 U5518 ( .A(n11685), .ZN(n11686) );
  INV_X1 U5519 ( .A(n1834), .ZN(n11924) );
  BUF_X1 U5520 ( .A(n11925), .Z(n11687) );
  INV_X1 U5521 ( .A(n63960), .ZN(n11688) );
  INV_X1 U5522 ( .A(n11688), .ZN(n11689) );
  INV_X1 U5523 ( .A(n1833), .ZN(n11931) );
  BUF_X1 U5524 ( .A(n11932), .Z(n11690) );
  INV_X1 U5525 ( .A(n63970), .ZN(n11691) );
  INV_X1 U5526 ( .A(n11691), .ZN(n11692) );
  INV_X1 U5527 ( .A(n1832), .ZN(n11938) );
  BUF_X1 U5528 ( .A(n11939), .Z(n11693) );
  INV_X1 U5529 ( .A(n63980), .ZN(n11694) );
  INV_X1 U5530 ( .A(n11694), .ZN(n11695) );
  INV_X1 U5531 ( .A(n1831), .ZN(n11945) );
  BUF_X1 U5532 ( .A(n11946), .Z(n11696) );
  INV_X1 U5533 ( .A(n63990), .ZN(n11697) );
  INV_X1 U5534 ( .A(n11697), .ZN(n11698) );
  INV_X1 U5535 ( .A(n1830), .ZN(n11952) );
  BUF_X1 U5536 ( .A(n11953), .Z(n11699) );
  INV_X1 U5537 ( .A(n64000), .ZN(n11700) );
  INV_X1 U5538 ( .A(n11700), .ZN(n11701) );
  INV_X1 U5539 ( .A(n1829), .ZN(n11959) );
  BUF_X1 U5540 ( .A(n11960), .Z(n11702) );
  INV_X1 U5541 ( .A(n64010), .ZN(n11703) );
  INV_X1 U5542 ( .A(n11703), .ZN(n11704) );
  INV_X1 U5543 ( .A(n1828), .ZN(n11966) );
  BUF_X1 U5544 ( .A(n11967), .Z(n11705) );
  INV_X1 U5545 ( .A(n64020), .ZN(n11706) );
  INV_X1 U5546 ( .A(n11706), .ZN(n11707) );
  INV_X1 U5547 ( .A(n1827), .ZN(n11973) );
  BUF_X1 U5548 ( .A(n11974), .Z(n11708) );
  INV_X1 U5549 ( .A(n64030), .ZN(n11709) );
  INV_X1 U5550 ( .A(n11709), .ZN(n11710) );
  INV_X1 U5551 ( .A(n1826), .ZN(n11980) );
  BUF_X1 U5552 ( .A(n11981), .Z(n11711) );
  INV_X1 U5553 ( .A(n64040), .ZN(n11712) );
  INV_X1 U5554 ( .A(n11712), .ZN(n11713) );
  INV_X1 U5555 ( .A(n1825), .ZN(n11987) );
  BUF_X1 U5556 ( .A(n11988), .Z(n11714) );
  INV_X1 U5557 ( .A(n64050), .ZN(n11715) );
  INV_X1 U5558 ( .A(n11715), .ZN(n11716) );
  INV_X1 U5559 ( .A(n1824), .ZN(n11994) );
  BUF_X1 U5560 ( .A(n11995), .Z(n11717) );
  INV_X1 U5561 ( .A(n64060), .ZN(n11718) );
  INV_X1 U5562 ( .A(n11718), .ZN(n11719) );
  INV_X1 U5563 ( .A(n1823), .ZN(n12001) );
  BUF_X1 U5564 ( .A(n12002), .Z(n11720) );
  INV_X1 U5565 ( .A(n64070), .ZN(n11721) );
  INV_X1 U5566 ( .A(n11721), .ZN(n11722) );
  INV_X1 U5567 ( .A(n1822), .ZN(n12008) );
  BUF_X1 U5568 ( .A(n12009), .Z(n11723) );
  INV_X1 U5569 ( .A(n64080), .ZN(n11724) );
  INV_X1 U5570 ( .A(n11724), .ZN(n11725) );
  INV_X1 U5571 ( .A(n1821), .ZN(n12015) );
  BUF_X1 U5572 ( .A(n12016), .Z(n11726) );
  INV_X1 U5573 ( .A(n64090), .ZN(n11727) );
  INV_X1 U5574 ( .A(n11727), .ZN(n11728) );
  INV_X1 U5575 ( .A(n1820), .ZN(n12022) );
  BUF_X1 U5576 ( .A(n12023), .Z(n11729) );
  INV_X1 U5577 ( .A(n64100), .ZN(n11730) );
  INV_X1 U5578 ( .A(n11730), .ZN(n11731) );
  INV_X1 U5579 ( .A(n1819), .ZN(n12029) );
  BUF_X1 U5580 ( .A(n12030), .Z(n11732) );
  INV_X1 U5581 ( .A(n64110), .ZN(n11733) );
  INV_X1 U5582 ( .A(n11733), .ZN(n11734) );
  INV_X1 U5583 ( .A(n1818), .ZN(n12036) );
  BUF_X1 U5584 ( .A(n12037), .Z(n11735) );
  INV_X1 U5585 ( .A(n6412), .ZN(n11736) );
  INV_X1 U5586 ( .A(n11736), .ZN(n11737) );
  INV_X1 U5587 ( .A(n1817), .ZN(n12043) );
  BUF_X1 U5588 ( .A(n12044), .Z(n11738) );
  INV_X1 U5589 ( .A(n6413), .ZN(n11739) );
  INV_X1 U5590 ( .A(n11739), .ZN(n11740) );
  INV_X1 U5591 ( .A(n1816), .ZN(n12050) );
  BUF_X1 U5592 ( .A(n12051), .Z(n11741) );
  INV_X1 U5593 ( .A(n6414), .ZN(n11742) );
  INV_X1 U5594 ( .A(n11742), .ZN(n11743) );
  INV_X1 U5595 ( .A(n1815), .ZN(n12057) );
  BUF_X1 U5596 ( .A(n12058), .Z(n11744) );
  INV_X1 U5597 ( .A(n6415), .ZN(n11745) );
  INV_X1 U5598 ( .A(n11745), .ZN(n11746) );
  INV_X1 U5599 ( .A(n1814), .ZN(n12064) );
  BUF_X1 U5600 ( .A(n12065), .Z(n11747) );
  INV_X1 U5601 ( .A(n6416), .ZN(n11748) );
  INV_X1 U5602 ( .A(n11748), .ZN(n11749) );
  INV_X1 U5603 ( .A(n1813), .ZN(n12071) );
  BUF_X1 U5604 ( .A(n12072), .Z(n11750) );
  INV_X1 U5605 ( .A(n6417), .ZN(n11751) );
  INV_X1 U5606 ( .A(n11751), .ZN(n11752) );
  INV_X1 U5607 ( .A(n1812), .ZN(n12078) );
  BUF_X1 U5608 ( .A(n12079), .Z(n11753) );
  INV_X1 U5609 ( .A(n6418), .ZN(n11754) );
  INV_X1 U5610 ( .A(n11754), .ZN(n11755) );
  INV_X1 U5611 ( .A(n1811), .ZN(n12085) );
  BUF_X1 U5612 ( .A(n12086), .Z(n11756) );
  INV_X1 U5613 ( .A(n6419), .ZN(n11757) );
  INV_X1 U5614 ( .A(n11757), .ZN(n11758) );
  INV_X1 U5615 ( .A(n1810), .ZN(n12092) );
  BUF_X1 U5616 ( .A(n12093), .Z(n11759) );
  INV_X1 U5617 ( .A(n6420), .ZN(n11760) );
  INV_X1 U5618 ( .A(n11760), .ZN(n11761) );
  INV_X1 U5619 ( .A(n1809), .ZN(n12099) );
  BUF_X1 U5620 ( .A(n12100), .Z(n11762) );
  INV_X1 U5621 ( .A(n6421), .ZN(n11763) );
  INV_X1 U5622 ( .A(n11763), .ZN(n11764) );
  INV_X1 U5623 ( .A(n1808), .ZN(n12106) );
  BUF_X1 U5624 ( .A(n12107), .Z(n11765) );
  INV_X1 U5625 ( .A(n6422), .ZN(n11766) );
  INV_X1 U5626 ( .A(n11766), .ZN(n11767) );
  INV_X1 U5627 ( .A(n1807), .ZN(n12113) );
  BUF_X1 U5628 ( .A(n12114), .Z(n11768) );
  INV_X1 U5629 ( .A(n6423), .ZN(n11769) );
  INV_X1 U5630 ( .A(n11769), .ZN(n11770) );
  INV_X1 U5631 ( .A(n1806), .ZN(n12120) );
  BUF_X1 U5632 ( .A(n12121), .Z(n11771) );
  INV_X1 U5633 ( .A(n6424), .ZN(n11772) );
  INV_X1 U5634 ( .A(n11772), .ZN(n11773) );
  INV_X1 U5635 ( .A(n1805), .ZN(n12127) );
  BUF_X1 U5636 ( .A(n12128), .Z(n11774) );
  INV_X1 U5637 ( .A(n6425), .ZN(n11775) );
  INV_X1 U5638 ( .A(n11775), .ZN(n11776) );
  INV_X1 U5639 ( .A(n1804), .ZN(n12134) );
  BUF_X1 U5640 ( .A(n12135), .Z(n11777) );
  INV_X1 U5641 ( .A(n6426), .ZN(n11778) );
  INV_X1 U5642 ( .A(n11778), .ZN(n11779) );
  INV_X1 U5643 ( .A(n1803), .ZN(n12141) );
  BUF_X1 U5644 ( .A(n12142), .Z(n11780) );
  INV_X1 U5645 ( .A(n6427), .ZN(n11781) );
  INV_X1 U5646 ( .A(n11781), .ZN(n11782) );
  INV_X1 U5647 ( .A(n1802), .ZN(n12148) );
  BUF_X1 U5648 ( .A(n12149), .Z(n11783) );
  INV_X1 U5649 ( .A(n6428), .ZN(n11784) );
  INV_X1 U5650 ( .A(n11784), .ZN(n11785) );
  INV_X1 U5651 ( .A(n1801), .ZN(n12155) );
  BUF_X1 U5652 ( .A(n12156), .Z(n11786) );
  INV_X1 U5653 ( .A(n64290), .ZN(n11787) );
  INV_X1 U5654 ( .A(n11787), .ZN(n11788) );
  INV_X1 U5655 ( .A(n1800), .ZN(n12162) );
  BUF_X1 U5656 ( .A(n12163), .Z(n11789) );
  INV_X1 U5657 ( .A(n64300), .ZN(n11790) );
  INV_X1 U5658 ( .A(n11790), .ZN(n11791) );
  INV_X1 U5659 ( .A(n1799), .ZN(n12169) );
  BUF_X1 U5660 ( .A(n12170), .Z(n11792) );
  INV_X1 U5661 ( .A(n64310), .ZN(n11793) );
  INV_X1 U5662 ( .A(n11793), .ZN(n11794) );
  INV_X1 U5663 ( .A(n1798), .ZN(n12176) );
  BUF_X1 U5664 ( .A(n12177), .Z(n11795) );
  INV_X1 U5665 ( .A(n64320), .ZN(n11796) );
  INV_X1 U5666 ( .A(n11796), .ZN(n11797) );
  INV_X1 U5667 ( .A(n1797), .ZN(n12183) );
  BUF_X1 U5668 ( .A(n12184), .Z(n11798) );
  INV_X1 U5669 ( .A(n64330), .ZN(n11799) );
  INV_X1 U5670 ( .A(n11799), .ZN(n11800) );
  INV_X1 U5671 ( .A(n1796), .ZN(n12190) );
  BUF_X1 U5672 ( .A(n12191), .Z(n11801) );
  INV_X1 U5673 ( .A(n64340), .ZN(n11802) );
  INV_X1 U5674 ( .A(n11802), .ZN(n11803) );
  INV_X1 U5675 ( .A(n1795), .ZN(n12197) );
  BUF_X1 U5676 ( .A(n12198), .Z(n11804) );
  INV_X1 U5677 ( .A(n64350), .ZN(n11805) );
  INV_X1 U5678 ( .A(n11805), .ZN(n11806) );
  INV_X1 U5679 ( .A(n1794), .ZN(n12204) );
  BUF_X1 U5680 ( .A(n12205), .Z(n11807) );
  INV_X1 U5681 ( .A(n64360), .ZN(n11808) );
  INV_X1 U5682 ( .A(n11808), .ZN(n11809) );
  INV_X1 U5683 ( .A(n1793), .ZN(n12211) );
  BUF_X1 U5684 ( .A(n12212), .Z(n11810) );
  INV_X1 U5685 ( .A(n64370), .ZN(n11811) );
  INV_X1 U5686 ( .A(n11811), .ZN(n11812) );
  INV_X1 U5687 ( .A(n1792), .ZN(n12218) );
  BUF_X1 U5688 ( .A(n12219), .Z(n11813) );
  INV_X1 U5689 ( .A(n64380), .ZN(n11814) );
  INV_X1 U5690 ( .A(n11814), .ZN(n11815) );
  INV_X1 U5691 ( .A(n1791), .ZN(n12225) );
  BUF_X1 U5692 ( .A(n12226), .Z(n11816) );
  INV_X1 U5693 ( .A(n64390), .ZN(n11817) );
  INV_X1 U5694 ( .A(n11817), .ZN(n11818) );
  INV_X1 U5695 ( .A(n1790), .ZN(n12232) );
  BUF_X1 U5696 ( .A(n12233), .Z(n11819) );
  INV_X1 U5697 ( .A(n64400), .ZN(n11820) );
  INV_X1 U5698 ( .A(n11820), .ZN(n11821) );
  INV_X1 U5699 ( .A(n1789), .ZN(n12239) );
  BUF_X1 U5700 ( .A(n12240), .Z(n11822) );
  INV_X1 U5701 ( .A(n64410), .ZN(n11823) );
  INV_X1 U5702 ( .A(n11823), .ZN(n11824) );
  INV_X1 U5703 ( .A(n1788), .ZN(n12246) );
  BUF_X1 U5704 ( .A(n12247), .Z(n11825) );
  INV_X1 U5705 ( .A(n64420), .ZN(n11826) );
  INV_X1 U5706 ( .A(n11826), .ZN(n11827) );
  INV_X1 U5707 ( .A(n1787), .ZN(n12253) );
  BUF_X1 U5708 ( .A(n12254), .Z(n11828) );
  INV_X1 U5709 ( .A(n64430), .ZN(n11829) );
  INV_X1 U5710 ( .A(n11829), .ZN(n11830) );
  INV_X1 U5711 ( .A(n1786), .ZN(n12260) );
  BUF_X1 U5712 ( .A(n12261), .Z(n11831) );
  INV_X1 U5713 ( .A(n64440), .ZN(n11832) );
  INV_X1 U5714 ( .A(n11832), .ZN(n11833) );
  INV_X1 U5715 ( .A(n1785), .ZN(n12267) );
  BUF_X1 U5716 ( .A(n12268), .Z(n11834) );
  INV_X1 U5717 ( .A(n64450), .ZN(n11835) );
  INV_X1 U5718 ( .A(n11835), .ZN(n11836) );
  INV_X1 U5719 ( .A(n1784), .ZN(n12274) );
  BUF_X1 U5720 ( .A(n12275), .Z(n11837) );
  INV_X1 U5721 ( .A(n64460), .ZN(n11838) );
  INV_X1 U5722 ( .A(n11838), .ZN(n11839) );
  INV_X1 U5723 ( .A(n1783), .ZN(n12281) );
  BUF_X1 U5724 ( .A(n12282), .Z(n11840) );
  INV_X1 U5725 ( .A(n64470), .ZN(n11841) );
  INV_X1 U5726 ( .A(n11841), .ZN(n11842) );
  INV_X1 U5727 ( .A(n1782), .ZN(n12288) );
  BUF_X1 U5728 ( .A(n12289), .Z(n11843) );
  INV_X1 U5729 ( .A(n64480), .ZN(n11844) );
  INV_X1 U5730 ( .A(n11844), .ZN(n11845) );
  INV_X1 U5731 ( .A(n1781), .ZN(n12295) );
  BUF_X1 U5732 ( .A(n12296), .Z(n11846) );
  INV_X1 U5733 ( .A(n64490), .ZN(n11847) );
  INV_X1 U5734 ( .A(n11847), .ZN(n11848) );
  BUF_X1 U5735 ( .A(n11851), .Z(n11849) );
  INV_X1 U5736 ( .A(n11853), .ZN(n11850) );
  INV_X1 U5737 ( .A(n11850), .ZN(n11851) );
  INV_X1 U5738 ( .A(n6897), .ZN(n11852) );
  INV_X1 U5739 ( .A(n11852), .ZN(n11853) );
  INV_X1 U5740 ( .A(n11854), .ZN(n11855) );
  BUF_X1 U5741 ( .A(n11858), .Z(n11856) );
  INV_X1 U5742 ( .A(n11860), .ZN(n11857) );
  INV_X1 U5743 ( .A(n11857), .ZN(n11858) );
  INV_X1 U5744 ( .A(n6896), .ZN(n11859) );
  INV_X1 U5745 ( .A(n11859), .ZN(n11860) );
  INV_X1 U5746 ( .A(n11861), .ZN(n11862) );
  BUF_X1 U5747 ( .A(n11865), .Z(n11863) );
  INV_X1 U5748 ( .A(n11867), .ZN(n11864) );
  INV_X1 U5749 ( .A(n11864), .ZN(n11865) );
  INV_X1 U5750 ( .A(n6895), .ZN(n11866) );
  INV_X1 U5751 ( .A(n11866), .ZN(n11867) );
  INV_X1 U5752 ( .A(n11868), .ZN(n11869) );
  BUF_X1 U5753 ( .A(n11872), .Z(n11870) );
  INV_X1 U5754 ( .A(n11874), .ZN(n11871) );
  INV_X1 U5755 ( .A(n11871), .ZN(n11872) );
  INV_X1 U5756 ( .A(n68940), .ZN(n11873) );
  INV_X1 U5757 ( .A(n11873), .ZN(n11874) );
  INV_X1 U5758 ( .A(n11875), .ZN(n11876) );
  BUF_X1 U5759 ( .A(n11879), .Z(n11877) );
  INV_X1 U5760 ( .A(n11881), .ZN(n11878) );
  INV_X1 U5761 ( .A(n11878), .ZN(n11879) );
  INV_X1 U5762 ( .A(n68930), .ZN(n11880) );
  INV_X1 U5763 ( .A(n11880), .ZN(n11881) );
  INV_X1 U5764 ( .A(n11882), .ZN(n11883) );
  BUF_X1 U5765 ( .A(n11886), .Z(n11884) );
  INV_X1 U5766 ( .A(n11888), .ZN(n11885) );
  INV_X1 U5767 ( .A(n11885), .ZN(n11886) );
  INV_X1 U5768 ( .A(n68920), .ZN(n11887) );
  INV_X1 U5769 ( .A(n11887), .ZN(n11888) );
  INV_X1 U5770 ( .A(n11889), .ZN(n11890) );
  BUF_X1 U5771 ( .A(n11893), .Z(n11891) );
  INV_X1 U5772 ( .A(n11895), .ZN(n11892) );
  INV_X1 U5773 ( .A(n11892), .ZN(n11893) );
  INV_X1 U5774 ( .A(n68910), .ZN(n11894) );
  INV_X1 U5775 ( .A(n11894), .ZN(n11895) );
  INV_X1 U5776 ( .A(n11896), .ZN(n11897) );
  BUF_X1 U5777 ( .A(n11900), .Z(n11898) );
  INV_X1 U5778 ( .A(n11902), .ZN(n11899) );
  INV_X1 U5779 ( .A(n11899), .ZN(n11900) );
  INV_X1 U5780 ( .A(n68900), .ZN(n11901) );
  INV_X1 U5781 ( .A(n11901), .ZN(n11902) );
  INV_X1 U5782 ( .A(n11903), .ZN(n11904) );
  BUF_X1 U5783 ( .A(n11907), .Z(n11905) );
  INV_X1 U5784 ( .A(n11909), .ZN(n11906) );
  INV_X1 U5785 ( .A(n11906), .ZN(n11907) );
  INV_X1 U5786 ( .A(n68890), .ZN(n11908) );
  INV_X1 U5787 ( .A(n11908), .ZN(n11909) );
  INV_X1 U5788 ( .A(n11910), .ZN(n11911) );
  BUF_X1 U5789 ( .A(n11914), .Z(n11912) );
  INV_X1 U5790 ( .A(n11916), .ZN(n11913) );
  INV_X1 U5791 ( .A(n11913), .ZN(n11914) );
  INV_X1 U5792 ( .A(n68880), .ZN(n11915) );
  INV_X1 U5793 ( .A(n11915), .ZN(n11916) );
  INV_X1 U5794 ( .A(n11917), .ZN(n11918) );
  BUF_X1 U5795 ( .A(n11921), .Z(n11919) );
  INV_X1 U5796 ( .A(n11923), .ZN(n11920) );
  INV_X1 U5797 ( .A(n11920), .ZN(n11921) );
  INV_X1 U5798 ( .A(n68870), .ZN(n11922) );
  INV_X1 U5799 ( .A(n11922), .ZN(n11923) );
  INV_X1 U5800 ( .A(n11924), .ZN(n11925) );
  BUF_X1 U5801 ( .A(n11928), .Z(n11926) );
  INV_X1 U5802 ( .A(n11930), .ZN(n11927) );
  INV_X1 U5803 ( .A(n11927), .ZN(n11928) );
  INV_X1 U5804 ( .A(n68860), .ZN(n11929) );
  INV_X1 U5805 ( .A(n11929), .ZN(n11930) );
  INV_X1 U5806 ( .A(n11931), .ZN(n11932) );
  BUF_X1 U5807 ( .A(n11935), .Z(n11933) );
  INV_X1 U5808 ( .A(n11937), .ZN(n11934) );
  INV_X1 U5809 ( .A(n11934), .ZN(n11935) );
  INV_X1 U5810 ( .A(n68850), .ZN(n11936) );
  INV_X1 U5811 ( .A(n11936), .ZN(n11937) );
  INV_X1 U5812 ( .A(n11938), .ZN(n11939) );
  BUF_X1 U5813 ( .A(n11942), .Z(n11940) );
  INV_X1 U5814 ( .A(n11944), .ZN(n11941) );
  INV_X1 U5815 ( .A(n11941), .ZN(n11942) );
  INV_X1 U5816 ( .A(n68840), .ZN(n11943) );
  INV_X1 U5817 ( .A(n11943), .ZN(n11944) );
  INV_X1 U5818 ( .A(n11945), .ZN(n11946) );
  BUF_X1 U5819 ( .A(n11949), .Z(n11947) );
  INV_X1 U5820 ( .A(n11951), .ZN(n11948) );
  INV_X1 U5821 ( .A(n11948), .ZN(n11949) );
  INV_X1 U5822 ( .A(n68830), .ZN(n11950) );
  INV_X1 U5823 ( .A(n11950), .ZN(n11951) );
  INV_X1 U5824 ( .A(n11952), .ZN(n11953) );
  BUF_X1 U5825 ( .A(n11956), .Z(n11954) );
  INV_X1 U5826 ( .A(n11958), .ZN(n11955) );
  INV_X1 U5827 ( .A(n11955), .ZN(n11956) );
  INV_X1 U5828 ( .A(n68820), .ZN(n11957) );
  INV_X1 U5829 ( .A(n11957), .ZN(n11958) );
  INV_X1 U5830 ( .A(n11959), .ZN(n11960) );
  BUF_X1 U5831 ( .A(n11963), .Z(n11961) );
  INV_X1 U5832 ( .A(n11965), .ZN(n11962) );
  INV_X1 U5833 ( .A(n11962), .ZN(n11963) );
  INV_X1 U5834 ( .A(n68810), .ZN(n11964) );
  INV_X1 U5835 ( .A(n11964), .ZN(n11965) );
  INV_X1 U5836 ( .A(n11966), .ZN(n11967) );
  BUF_X1 U5837 ( .A(n11970), .Z(n11968) );
  INV_X1 U5838 ( .A(n11972), .ZN(n11969) );
  INV_X1 U5839 ( .A(n11969), .ZN(n11970) );
  INV_X1 U5840 ( .A(n68800), .ZN(n11971) );
  INV_X1 U5841 ( .A(n11971), .ZN(n11972) );
  INV_X1 U5842 ( .A(n11973), .ZN(n11974) );
  BUF_X1 U5843 ( .A(n11977), .Z(n11975) );
  INV_X1 U5844 ( .A(n11979), .ZN(n11976) );
  INV_X1 U5845 ( .A(n11976), .ZN(n11977) );
  INV_X1 U5846 ( .A(n68790), .ZN(n11978) );
  INV_X1 U5847 ( .A(n11978), .ZN(n11979) );
  INV_X1 U5848 ( .A(n11980), .ZN(n11981) );
  BUF_X1 U5849 ( .A(n11984), .Z(n11982) );
  INV_X1 U5850 ( .A(n11986), .ZN(n11983) );
  INV_X1 U5851 ( .A(n11983), .ZN(n11984) );
  INV_X1 U5852 ( .A(n68780), .ZN(n11985) );
  INV_X1 U5853 ( .A(n11985), .ZN(n11986) );
  INV_X1 U5854 ( .A(n11987), .ZN(n11988) );
  BUF_X1 U5855 ( .A(n11991), .Z(n11989) );
  INV_X1 U5856 ( .A(n11993), .ZN(n11990) );
  INV_X1 U5857 ( .A(n11990), .ZN(n11991) );
  INV_X1 U5858 ( .A(n68770), .ZN(n11992) );
  INV_X1 U5859 ( .A(n11992), .ZN(n11993) );
  INV_X1 U5860 ( .A(n11994), .ZN(n11995) );
  BUF_X1 U5861 ( .A(n11998), .Z(n11996) );
  INV_X1 U5862 ( .A(n12000), .ZN(n11997) );
  INV_X1 U5863 ( .A(n11997), .ZN(n11998) );
  INV_X1 U5864 ( .A(n68760), .ZN(n11999) );
  INV_X1 U5865 ( .A(n11999), .ZN(n12000) );
  INV_X1 U5866 ( .A(n12001), .ZN(n12002) );
  BUF_X1 U5867 ( .A(n12005), .Z(n12003) );
  INV_X1 U5868 ( .A(n12007), .ZN(n12004) );
  INV_X1 U5869 ( .A(n12004), .ZN(n12005) );
  INV_X1 U5870 ( .A(n68750), .ZN(n12006) );
  INV_X1 U5871 ( .A(n12006), .ZN(n12007) );
  INV_X1 U5872 ( .A(n12008), .ZN(n12009) );
  BUF_X1 U5873 ( .A(n12012), .Z(n12010) );
  INV_X1 U5874 ( .A(n12014), .ZN(n12011) );
  INV_X1 U5875 ( .A(n12011), .ZN(n12012) );
  INV_X1 U5876 ( .A(n68740), .ZN(n12013) );
  INV_X1 U5877 ( .A(n12013), .ZN(n12014) );
  INV_X1 U5878 ( .A(n12015), .ZN(n12016) );
  BUF_X1 U5879 ( .A(n12019), .Z(n12017) );
  INV_X1 U5880 ( .A(n12021), .ZN(n12018) );
  INV_X1 U5881 ( .A(n12018), .ZN(n12019) );
  INV_X1 U5882 ( .A(n6873), .ZN(n12020) );
  INV_X1 U5883 ( .A(n12020), .ZN(n12021) );
  INV_X1 U5884 ( .A(n12022), .ZN(n12023) );
  BUF_X1 U5885 ( .A(n12026), .Z(n12024) );
  INV_X1 U5886 ( .A(n12028), .ZN(n12025) );
  INV_X1 U5887 ( .A(n12025), .ZN(n12026) );
  INV_X1 U5888 ( .A(n6872), .ZN(n12027) );
  INV_X1 U5889 ( .A(n12027), .ZN(n12028) );
  INV_X1 U5890 ( .A(n12029), .ZN(n12030) );
  BUF_X1 U5891 ( .A(n12033), .Z(n12031) );
  INV_X1 U5892 ( .A(n12035), .ZN(n12032) );
  INV_X1 U5893 ( .A(n12032), .ZN(n12033) );
  INV_X1 U5894 ( .A(n6871), .ZN(n12034) );
  INV_X1 U5895 ( .A(n12034), .ZN(n12035) );
  INV_X1 U5896 ( .A(n12036), .ZN(n12037) );
  BUF_X1 U5897 ( .A(n12040), .Z(n12038) );
  INV_X1 U5898 ( .A(n12042), .ZN(n12039) );
  INV_X1 U5899 ( .A(n12039), .ZN(n12040) );
  INV_X1 U5900 ( .A(n6870), .ZN(n12041) );
  INV_X1 U5901 ( .A(n12041), .ZN(n12042) );
  INV_X1 U5902 ( .A(n12043), .ZN(n12044) );
  BUF_X1 U5903 ( .A(n12047), .Z(n12045) );
  INV_X1 U5904 ( .A(n12049), .ZN(n12046) );
  INV_X1 U5905 ( .A(n12046), .ZN(n12047) );
  INV_X1 U5906 ( .A(n6869), .ZN(n12048) );
  INV_X1 U5907 ( .A(n12048), .ZN(n12049) );
  INV_X1 U5908 ( .A(n12050), .ZN(n12051) );
  BUF_X1 U5909 ( .A(n12054), .Z(n12052) );
  INV_X1 U5910 ( .A(n12056), .ZN(n12053) );
  INV_X1 U5911 ( .A(n12053), .ZN(n12054) );
  INV_X1 U5912 ( .A(n6868), .ZN(n12055) );
  INV_X1 U5913 ( .A(n12055), .ZN(n12056) );
  INV_X1 U5914 ( .A(n12057), .ZN(n12058) );
  BUF_X1 U5915 ( .A(n12061), .Z(n12059) );
  INV_X1 U5916 ( .A(n12063), .ZN(n12060) );
  INV_X1 U5917 ( .A(n12060), .ZN(n12061) );
  INV_X1 U5918 ( .A(n6867), .ZN(n12062) );
  INV_X1 U5919 ( .A(n12062), .ZN(n12063) );
  INV_X1 U5920 ( .A(n12064), .ZN(n12065) );
  BUF_X1 U5921 ( .A(n12068), .Z(n12066) );
  INV_X1 U5922 ( .A(n12070), .ZN(n12067) );
  INV_X1 U5923 ( .A(n12067), .ZN(n12068) );
  INV_X1 U5924 ( .A(n6866), .ZN(n12069) );
  INV_X1 U5925 ( .A(n12069), .ZN(n12070) );
  INV_X1 U5926 ( .A(n12071), .ZN(n12072) );
  BUF_X1 U5927 ( .A(n12075), .Z(n12073) );
  INV_X1 U5928 ( .A(n12077), .ZN(n12074) );
  INV_X1 U5929 ( .A(n12074), .ZN(n12075) );
  INV_X1 U5930 ( .A(n6865), .ZN(n12076) );
  INV_X1 U5931 ( .A(n12076), .ZN(n12077) );
  INV_X1 U5932 ( .A(n12078), .ZN(n12079) );
  BUF_X1 U5933 ( .A(n12082), .Z(n12080) );
  INV_X1 U5934 ( .A(n12084), .ZN(n12081) );
  INV_X1 U5935 ( .A(n12081), .ZN(n12082) );
  INV_X1 U5936 ( .A(n6864), .ZN(n12083) );
  INV_X1 U5937 ( .A(n12083), .ZN(n12084) );
  INV_X1 U5938 ( .A(n12085), .ZN(n12086) );
  BUF_X1 U5939 ( .A(n12089), .Z(n12087) );
  INV_X1 U5940 ( .A(n12091), .ZN(n12088) );
  INV_X1 U5941 ( .A(n12088), .ZN(n12089) );
  INV_X1 U5942 ( .A(n6863), .ZN(n12090) );
  INV_X1 U5943 ( .A(n12090), .ZN(n12091) );
  INV_X1 U5944 ( .A(n12092), .ZN(n12093) );
  BUF_X1 U5945 ( .A(n12096), .Z(n12094) );
  INV_X1 U5946 ( .A(n12098), .ZN(n12095) );
  INV_X1 U5947 ( .A(n12095), .ZN(n12096) );
  INV_X1 U5948 ( .A(n6862), .ZN(n12097) );
  INV_X1 U5949 ( .A(n12097), .ZN(n12098) );
  INV_X1 U5950 ( .A(n12099), .ZN(n12100) );
  BUF_X1 U5951 ( .A(n12103), .Z(n12101) );
  INV_X1 U5952 ( .A(n12105), .ZN(n12102) );
  INV_X1 U5953 ( .A(n12102), .ZN(n12103) );
  INV_X1 U5954 ( .A(n6861), .ZN(n12104) );
  INV_X1 U5955 ( .A(n12104), .ZN(n12105) );
  INV_X1 U5956 ( .A(n12106), .ZN(n12107) );
  BUF_X1 U5957 ( .A(n12110), .Z(n12108) );
  INV_X1 U5958 ( .A(n12112), .ZN(n12109) );
  INV_X1 U5959 ( .A(n12109), .ZN(n12110) );
  INV_X1 U5960 ( .A(n6860), .ZN(n12111) );
  INV_X1 U5961 ( .A(n12111), .ZN(n12112) );
  INV_X1 U5962 ( .A(n12113), .ZN(n12114) );
  BUF_X1 U5963 ( .A(n12117), .Z(n12115) );
  INV_X1 U5964 ( .A(n12119), .ZN(n12116) );
  INV_X1 U5965 ( .A(n12116), .ZN(n12117) );
  INV_X1 U5966 ( .A(n6859), .ZN(n12118) );
  INV_X1 U5967 ( .A(n12118), .ZN(n12119) );
  INV_X1 U5968 ( .A(n12120), .ZN(n12121) );
  BUF_X1 U5969 ( .A(n12124), .Z(n12122) );
  INV_X1 U5970 ( .A(n12126), .ZN(n12123) );
  INV_X1 U5971 ( .A(n12123), .ZN(n12124) );
  INV_X1 U5972 ( .A(n6858), .ZN(n12125) );
  INV_X1 U5973 ( .A(n12125), .ZN(n12126) );
  INV_X1 U5974 ( .A(n12127), .ZN(n12128) );
  BUF_X1 U5975 ( .A(n12131), .Z(n12129) );
  INV_X1 U5976 ( .A(n12133), .ZN(n12130) );
  INV_X1 U5977 ( .A(n12130), .ZN(n12131) );
  INV_X1 U5978 ( .A(n6857), .ZN(n12132) );
  INV_X1 U5979 ( .A(n12132), .ZN(n12133) );
  INV_X1 U5980 ( .A(n12134), .ZN(n12135) );
  BUF_X1 U5981 ( .A(n12138), .Z(n12136) );
  INV_X1 U5982 ( .A(n12140), .ZN(n12137) );
  INV_X1 U5983 ( .A(n12137), .ZN(n12138) );
  INV_X1 U5984 ( .A(n68560), .ZN(n12139) );
  INV_X1 U5985 ( .A(n12139), .ZN(n12140) );
  INV_X1 U5986 ( .A(n12141), .ZN(n12142) );
  BUF_X1 U5987 ( .A(n12145), .Z(n12143) );
  INV_X1 U5988 ( .A(n12147), .ZN(n12144) );
  INV_X1 U5989 ( .A(n12144), .ZN(n12145) );
  INV_X1 U5990 ( .A(n68550), .ZN(n12146) );
  INV_X1 U5991 ( .A(n12146), .ZN(n12147) );
  INV_X1 U5992 ( .A(n12148), .ZN(n12149) );
  BUF_X1 U5993 ( .A(n12152), .Z(n12150) );
  INV_X1 U5994 ( .A(n12154), .ZN(n12151) );
  INV_X1 U5995 ( .A(n12151), .ZN(n12152) );
  INV_X1 U5996 ( .A(n68540), .ZN(n12153) );
  INV_X1 U5997 ( .A(n12153), .ZN(n12154) );
  INV_X1 U5998 ( .A(n12155), .ZN(n12156) );
  BUF_X1 U5999 ( .A(n12159), .Z(n12157) );
  INV_X1 U6000 ( .A(n12161), .ZN(n12158) );
  INV_X1 U6001 ( .A(n12158), .ZN(n12159) );
  INV_X1 U6002 ( .A(n68530), .ZN(n12160) );
  INV_X1 U6003 ( .A(n12160), .ZN(n12161) );
  INV_X1 U6004 ( .A(n12162), .ZN(n12163) );
  BUF_X1 U6005 ( .A(n12166), .Z(n12164) );
  INV_X1 U6006 ( .A(n12168), .ZN(n12165) );
  INV_X1 U6007 ( .A(n12165), .ZN(n12166) );
  INV_X1 U6008 ( .A(n68520), .ZN(n12167) );
  INV_X1 U6009 ( .A(n12167), .ZN(n12168) );
  INV_X1 U6010 ( .A(n12169), .ZN(n12170) );
  BUF_X1 U6011 ( .A(n12173), .Z(n12171) );
  INV_X1 U6012 ( .A(n12175), .ZN(n12172) );
  INV_X1 U6013 ( .A(n12172), .ZN(n12173) );
  INV_X1 U6014 ( .A(n68510), .ZN(n12174) );
  INV_X1 U6015 ( .A(n12174), .ZN(n12175) );
  INV_X1 U6016 ( .A(n12176), .ZN(n12177) );
  BUF_X1 U6017 ( .A(n12180), .Z(n12178) );
  INV_X1 U6018 ( .A(n12182), .ZN(n12179) );
  INV_X1 U6019 ( .A(n12179), .ZN(n12180) );
  INV_X1 U6020 ( .A(n68500), .ZN(n12181) );
  INV_X1 U6021 ( .A(n12181), .ZN(n12182) );
  INV_X1 U6022 ( .A(n12183), .ZN(n12184) );
  BUF_X1 U6023 ( .A(n12187), .Z(n12185) );
  INV_X1 U6024 ( .A(n12189), .ZN(n12186) );
  INV_X1 U6025 ( .A(n12186), .ZN(n12187) );
  INV_X1 U6026 ( .A(n68490), .ZN(n12188) );
  INV_X1 U6027 ( .A(n12188), .ZN(n12189) );
  INV_X1 U6028 ( .A(n12190), .ZN(n12191) );
  BUF_X1 U6029 ( .A(n12194), .Z(n12192) );
  INV_X1 U6030 ( .A(n12196), .ZN(n12193) );
  INV_X1 U6031 ( .A(n12193), .ZN(n12194) );
  INV_X1 U6032 ( .A(n68480), .ZN(n12195) );
  INV_X1 U6033 ( .A(n12195), .ZN(n12196) );
  INV_X1 U6034 ( .A(n12197), .ZN(n12198) );
  BUF_X1 U6035 ( .A(n12201), .Z(n12199) );
  INV_X1 U6036 ( .A(n12203), .ZN(n12200) );
  INV_X1 U6037 ( .A(n12200), .ZN(n12201) );
  INV_X1 U6038 ( .A(n68470), .ZN(n12202) );
  INV_X1 U6039 ( .A(n12202), .ZN(n12203) );
  INV_X1 U6040 ( .A(n12204), .ZN(n12205) );
  BUF_X1 U6041 ( .A(n12208), .Z(n12206) );
  INV_X1 U6042 ( .A(n12210), .ZN(n12207) );
  INV_X1 U6043 ( .A(n12207), .ZN(n12208) );
  INV_X1 U6044 ( .A(n68460), .ZN(n12209) );
  INV_X1 U6045 ( .A(n12209), .ZN(n12210) );
  INV_X1 U6046 ( .A(n12211), .ZN(n12212) );
  BUF_X1 U6047 ( .A(n12215), .Z(n12213) );
  INV_X1 U6048 ( .A(n12217), .ZN(n12214) );
  INV_X1 U6049 ( .A(n12214), .ZN(n12215) );
  INV_X1 U6050 ( .A(n68450), .ZN(n12216) );
  INV_X1 U6051 ( .A(n12216), .ZN(n12217) );
  INV_X1 U6052 ( .A(n12218), .ZN(n12219) );
  BUF_X1 U6053 ( .A(n12222), .Z(n12220) );
  INV_X1 U6054 ( .A(n12224), .ZN(n12221) );
  INV_X1 U6055 ( .A(n12221), .ZN(n12222) );
  INV_X1 U6056 ( .A(n68440), .ZN(n12223) );
  INV_X1 U6057 ( .A(n12223), .ZN(n12224) );
  INV_X1 U6058 ( .A(n12225), .ZN(n12226) );
  BUF_X1 U6059 ( .A(n12229), .Z(n12227) );
  INV_X1 U6060 ( .A(n12231), .ZN(n12228) );
  INV_X1 U6061 ( .A(n12228), .ZN(n12229) );
  INV_X1 U6062 ( .A(n68430), .ZN(n12230) );
  INV_X1 U6063 ( .A(n12230), .ZN(n12231) );
  INV_X1 U6064 ( .A(n12232), .ZN(n12233) );
  BUF_X1 U6065 ( .A(n12236), .Z(n12234) );
  INV_X1 U6066 ( .A(n12238), .ZN(n12235) );
  INV_X1 U6067 ( .A(n12235), .ZN(n12236) );
  INV_X1 U6068 ( .A(n68420), .ZN(n12237) );
  INV_X1 U6069 ( .A(n12237), .ZN(n12238) );
  INV_X1 U6070 ( .A(n12239), .ZN(n12240) );
  BUF_X1 U6071 ( .A(n12243), .Z(n12241) );
  INV_X1 U6072 ( .A(n12245), .ZN(n12242) );
  INV_X1 U6073 ( .A(n12242), .ZN(n12243) );
  INV_X1 U6074 ( .A(n68410), .ZN(n12244) );
  INV_X1 U6075 ( .A(n12244), .ZN(n12245) );
  INV_X1 U6076 ( .A(n12246), .ZN(n12247) );
  BUF_X1 U6077 ( .A(n12250), .Z(n12248) );
  INV_X1 U6078 ( .A(n12252), .ZN(n12249) );
  INV_X1 U6079 ( .A(n12249), .ZN(n12250) );
  INV_X1 U6080 ( .A(n6840), .ZN(n12251) );
  INV_X1 U6081 ( .A(n12251), .ZN(n12252) );
  INV_X1 U6082 ( .A(n12253), .ZN(n12254) );
  BUF_X1 U6083 ( .A(n12257), .Z(n12255) );
  INV_X1 U6084 ( .A(n12259), .ZN(n12256) );
  INV_X1 U6085 ( .A(n12256), .ZN(n12257) );
  INV_X1 U6086 ( .A(n6839), .ZN(n12258) );
  INV_X1 U6087 ( .A(n12258), .ZN(n12259) );
  INV_X1 U6088 ( .A(n12260), .ZN(n12261) );
  BUF_X1 U6089 ( .A(n12264), .Z(n12262) );
  INV_X1 U6090 ( .A(n12266), .ZN(n12263) );
  INV_X1 U6091 ( .A(n12263), .ZN(n12264) );
  INV_X1 U6092 ( .A(n6838), .ZN(n12265) );
  INV_X1 U6093 ( .A(n12265), .ZN(n12266) );
  INV_X1 U6094 ( .A(n12267), .ZN(n12268) );
  BUF_X1 U6095 ( .A(n12271), .Z(n12269) );
  INV_X1 U6096 ( .A(n12273), .ZN(n12270) );
  INV_X1 U6097 ( .A(n12270), .ZN(n12271) );
  INV_X1 U6098 ( .A(n6837), .ZN(n12272) );
  INV_X1 U6099 ( .A(n12272), .ZN(n12273) );
  INV_X1 U6100 ( .A(n12274), .ZN(n12275) );
  BUF_X1 U6101 ( .A(n12278), .Z(n12276) );
  INV_X1 U6102 ( .A(n12280), .ZN(n12277) );
  INV_X1 U6103 ( .A(n12277), .ZN(n12278) );
  INV_X1 U6104 ( .A(n6836), .ZN(n12279) );
  INV_X1 U6105 ( .A(n12279), .ZN(n12280) );
  INV_X1 U6106 ( .A(n12281), .ZN(n12282) );
  BUF_X1 U6107 ( .A(n12285), .Z(n12283) );
  INV_X1 U6108 ( .A(n12287), .ZN(n12284) );
  INV_X1 U6109 ( .A(n12284), .ZN(n12285) );
  INV_X1 U6110 ( .A(n6835), .ZN(n12286) );
  INV_X1 U6111 ( .A(n12286), .ZN(n12287) );
  INV_X1 U6112 ( .A(n12288), .ZN(n12289) );
  BUF_X1 U6113 ( .A(n12292), .Z(n12290) );
  INV_X1 U6114 ( .A(n12294), .ZN(n12291) );
  INV_X1 U6115 ( .A(n12291), .ZN(n12292) );
  INV_X1 U6116 ( .A(n6834), .ZN(n12293) );
  INV_X1 U6117 ( .A(n12293), .ZN(n12294) );
  INV_X1 U6118 ( .A(n12295), .ZN(n12296) );
  BUF_X1 U6119 ( .A(n12299), .Z(n12297) );
  INV_X1 U6120 ( .A(n12301), .ZN(n12298) );
  INV_X1 U6121 ( .A(n12298), .ZN(n12299) );
  INV_X1 U6122 ( .A(n6833), .ZN(n12300) );
  INV_X1 U6123 ( .A(n12300), .ZN(n12301) );
  BUF_X1 U6124 ( .A(n12304), .Z(n12302) );
  INV_X1 U6125 ( .A(n12306), .ZN(n12303) );
  INV_X1 U6126 ( .A(n12303), .ZN(n12304) );
  INV_X1 U6127 ( .A(n6832), .ZN(n12305) );
  INV_X1 U6128 ( .A(n12305), .ZN(n12306) );
  BUF_X1 U6129 ( .A(n12309), .Z(n12307) );
  INV_X1 U6130 ( .A(n12311), .ZN(n12308) );
  INV_X1 U6131 ( .A(n12308), .ZN(n12309) );
  INV_X1 U6132 ( .A(n6831), .ZN(n12310) );
  INV_X1 U6133 ( .A(n12310), .ZN(n12311) );
  BUF_X1 U6134 ( .A(n12314), .Z(n12312) );
  INV_X1 U6135 ( .A(n12316), .ZN(n12313) );
  INV_X1 U6136 ( .A(n12313), .ZN(n12314) );
  INV_X1 U6137 ( .A(n6830), .ZN(n12315) );
  INV_X1 U6138 ( .A(n12315), .ZN(n12316) );
  BUF_X1 U6139 ( .A(n12319), .Z(n12317) );
  INV_X1 U6140 ( .A(n12321), .ZN(n12318) );
  INV_X1 U6141 ( .A(n12318), .ZN(n12319) );
  INV_X1 U6142 ( .A(n6829), .ZN(n12320) );
  INV_X1 U6143 ( .A(n12320), .ZN(n12321) );
  BUF_X1 U6144 ( .A(n12324), .Z(n12322) );
  INV_X1 U6145 ( .A(n12326), .ZN(n12323) );
  INV_X1 U6146 ( .A(n12323), .ZN(n12324) );
  INV_X1 U6147 ( .A(n6828), .ZN(n12325) );
  INV_X1 U6148 ( .A(n12325), .ZN(n12326) );
  BUF_X1 U6149 ( .A(n12329), .Z(n12327) );
  INV_X1 U6150 ( .A(n12331), .ZN(n12328) );
  INV_X1 U6151 ( .A(n12328), .ZN(n12329) );
  INV_X1 U6152 ( .A(n6827), .ZN(n12330) );
  INV_X1 U6153 ( .A(n12330), .ZN(n12331) );
  BUF_X1 U6154 ( .A(n12334), .Z(n12332) );
  INV_X1 U6155 ( .A(n12336), .ZN(n12333) );
  INV_X1 U6156 ( .A(n12333), .ZN(n12334) );
  INV_X1 U6157 ( .A(n6826), .ZN(n12335) );
  INV_X1 U6158 ( .A(n12335), .ZN(n12336) );
  BUF_X1 U6159 ( .A(n12339), .Z(n12337) );
  INV_X1 U6160 ( .A(n12341), .ZN(n12338) );
  INV_X1 U6161 ( .A(n12338), .ZN(n12339) );
  INV_X1 U6162 ( .A(n6825), .ZN(n12340) );
  INV_X1 U6163 ( .A(n12340), .ZN(n12341) );
  BUF_X1 U6164 ( .A(n12344), .Z(n12342) );
  INV_X1 U6165 ( .A(n12346), .ZN(n12343) );
  INV_X1 U6166 ( .A(n12343), .ZN(n12344) );
  INV_X1 U6167 ( .A(n6824), .ZN(n12345) );
  INV_X1 U6168 ( .A(n12345), .ZN(n12346) );
  BUF_X1 U6169 ( .A(n12349), .Z(n12347) );
  INV_X1 U6170 ( .A(n12351), .ZN(n12348) );
  INV_X1 U6171 ( .A(n12348), .ZN(n12349) );
  INV_X1 U6172 ( .A(n6823), .ZN(n12350) );
  INV_X1 U6173 ( .A(n12350), .ZN(n12351) );
  BUF_X1 U6174 ( .A(n12354), .Z(n12352) );
  INV_X1 U6175 ( .A(n12356), .ZN(n12353) );
  INV_X1 U6176 ( .A(n12353), .ZN(n12354) );
  INV_X1 U6177 ( .A(n6822), .ZN(n12355) );
  INV_X1 U6178 ( .A(n12355), .ZN(n12356) );
  BUF_X1 U6179 ( .A(n12359), .Z(n12357) );
  INV_X1 U6180 ( .A(n12361), .ZN(n12358) );
  INV_X1 U6181 ( .A(n12358), .ZN(n12359) );
  INV_X1 U6182 ( .A(n6821), .ZN(n12360) );
  INV_X1 U6183 ( .A(n12360), .ZN(n12361) );
  BUF_X1 U6184 ( .A(n12364), .Z(n12362) );
  INV_X1 U6185 ( .A(n12366), .ZN(n12363) );
  INV_X1 U6186 ( .A(n12363), .ZN(n12364) );
  INV_X1 U6187 ( .A(n6820), .ZN(n12365) );
  INV_X1 U6188 ( .A(n12365), .ZN(n12366) );
  BUF_X1 U6189 ( .A(n12369), .Z(n12367) );
  INV_X1 U6190 ( .A(n12371), .ZN(n12368) );
  INV_X1 U6191 ( .A(n12368), .ZN(n12369) );
  INV_X1 U6192 ( .A(n6819), .ZN(n12370) );
  INV_X1 U6193 ( .A(n12370), .ZN(n12371) );
  BUF_X1 U6194 ( .A(n12374), .Z(n12372) );
  INV_X1 U6195 ( .A(n12376), .ZN(n12373) );
  INV_X1 U6196 ( .A(n12373), .ZN(n12374) );
  INV_X1 U6197 ( .A(n6818), .ZN(n12375) );
  INV_X1 U6198 ( .A(n12375), .ZN(n12376) );
  BUF_X1 U6199 ( .A(n12379), .Z(n12377) );
  INV_X1 U6200 ( .A(n12381), .ZN(n12378) );
  INV_X1 U6201 ( .A(n12378), .ZN(n12379) );
  INV_X1 U6202 ( .A(n6817), .ZN(n12380) );
  INV_X1 U6203 ( .A(n12380), .ZN(n12381) );
  BUF_X1 U6204 ( .A(n12384), .Z(n12382) );
  INV_X1 U6205 ( .A(n12386), .ZN(n12383) );
  INV_X1 U6206 ( .A(n12383), .ZN(n12384) );
  INV_X1 U6207 ( .A(n6816), .ZN(n12385) );
  INV_X1 U6208 ( .A(n12385), .ZN(n12386) );
  BUF_X1 U6209 ( .A(n12389), .Z(n12387) );
  INV_X1 U6210 ( .A(n12391), .ZN(n12388) );
  INV_X1 U6211 ( .A(n12388), .ZN(n12389) );
  INV_X1 U6212 ( .A(n6815), .ZN(n12390) );
  INV_X1 U6213 ( .A(n12390), .ZN(n12391) );
  BUF_X1 U6214 ( .A(n12394), .Z(n12392) );
  INV_X1 U6215 ( .A(n12396), .ZN(n12393) );
  INV_X1 U6216 ( .A(n12393), .ZN(n12394) );
  INV_X1 U6217 ( .A(n6814), .ZN(n12395) );
  INV_X1 U6218 ( .A(n12395), .ZN(n12396) );
  BUF_X1 U6219 ( .A(n12399), .Z(n12397) );
  INV_X1 U6220 ( .A(n12401), .ZN(n12398) );
  INV_X1 U6221 ( .A(n12398), .ZN(n12399) );
  INV_X1 U6222 ( .A(n6813), .ZN(n12400) );
  INV_X1 U6223 ( .A(n12400), .ZN(n12401) );
  BUF_X1 U6224 ( .A(n12404), .Z(n12402) );
  INV_X1 U6225 ( .A(n12406), .ZN(n12403) );
  INV_X1 U6226 ( .A(n12403), .ZN(n12404) );
  INV_X1 U6227 ( .A(n6812), .ZN(n12405) );
  INV_X1 U6228 ( .A(n12405), .ZN(n12406) );
  BUF_X1 U6229 ( .A(n12409), .Z(n12407) );
  INV_X1 U6230 ( .A(n12411), .ZN(n12408) );
  INV_X1 U6231 ( .A(n12408), .ZN(n12409) );
  INV_X1 U6232 ( .A(n6811), .ZN(n12410) );
  INV_X1 U6233 ( .A(n12410), .ZN(n12411) );
  BUF_X1 U6234 ( .A(n12414), .Z(n12412) );
  INV_X1 U6235 ( .A(n12416), .ZN(n12413) );
  INV_X1 U6236 ( .A(n12413), .ZN(n12414) );
  INV_X1 U6237 ( .A(n6810), .ZN(n12415) );
  INV_X1 U6238 ( .A(n12415), .ZN(n12416) );
  BUF_X1 U6239 ( .A(n12419), .Z(n12417) );
  INV_X1 U6240 ( .A(n12421), .ZN(n12418) );
  INV_X1 U6241 ( .A(n12418), .ZN(n12419) );
  INV_X1 U6242 ( .A(n6809), .ZN(n12420) );
  INV_X1 U6243 ( .A(n12420), .ZN(n12421) );
  BUF_X1 U6244 ( .A(n12424), .Z(n12422) );
  INV_X1 U6245 ( .A(n12426), .ZN(n12423) );
  INV_X1 U6246 ( .A(n12423), .ZN(n12424) );
  INV_X1 U6247 ( .A(n6808), .ZN(n12425) );
  INV_X1 U6248 ( .A(n12425), .ZN(n12426) );
  BUF_X1 U6249 ( .A(n12429), .Z(n12427) );
  INV_X1 U6250 ( .A(n12431), .ZN(n12428) );
  INV_X1 U6251 ( .A(n12428), .ZN(n12429) );
  INV_X1 U6252 ( .A(n6807), .ZN(n12430) );
  INV_X1 U6253 ( .A(n12430), .ZN(n12431) );
  BUF_X1 U6254 ( .A(n12434), .Z(n12432) );
  INV_X1 U6255 ( .A(n12436), .ZN(n12433) );
  INV_X1 U6256 ( .A(n12433), .ZN(n12434) );
  INV_X1 U6257 ( .A(n6806), .ZN(n12435) );
  INV_X1 U6258 ( .A(n12435), .ZN(n12436) );
  BUF_X1 U6259 ( .A(n12439), .Z(n12437) );
  INV_X1 U6260 ( .A(n12441), .ZN(n12438) );
  INV_X1 U6261 ( .A(n12438), .ZN(n12439) );
  INV_X1 U6262 ( .A(n6805), .ZN(n12440) );
  INV_X1 U6263 ( .A(n12440), .ZN(n12441) );
  BUF_X1 U6264 ( .A(n12444), .Z(n12442) );
  INV_X1 U6265 ( .A(n12446), .ZN(n12443) );
  INV_X1 U6266 ( .A(n12443), .ZN(n12444) );
  INV_X1 U6267 ( .A(n6804), .ZN(n12445) );
  INV_X1 U6268 ( .A(n12445), .ZN(n12446) );
  BUF_X1 U6269 ( .A(n12449), .Z(n12447) );
  INV_X1 U6270 ( .A(n12451), .ZN(n12448) );
  INV_X1 U6271 ( .A(n12448), .ZN(n12449) );
  INV_X1 U6272 ( .A(n6803), .ZN(n12450) );
  INV_X1 U6273 ( .A(n12450), .ZN(n12451) );
  BUF_X1 U6274 ( .A(n12454), .Z(n12452) );
  INV_X1 U6275 ( .A(n12456), .ZN(n12453) );
  INV_X1 U6276 ( .A(n12453), .ZN(n12454) );
  INV_X1 U6277 ( .A(n68020), .ZN(n12455) );
  INV_X1 U6278 ( .A(n12455), .ZN(n12456) );
  BUF_X1 U6279 ( .A(n12459), .Z(n12457) );
  INV_X1 U6280 ( .A(n12461), .ZN(n12458) );
  INV_X1 U6281 ( .A(n12458), .ZN(n12459) );
  INV_X1 U6282 ( .A(n68010), .ZN(n12460) );
  INV_X1 U6283 ( .A(n12460), .ZN(n12461) );
  BUF_X1 U6284 ( .A(n12464), .Z(n12462) );
  INV_X1 U6285 ( .A(n12466), .ZN(n12463) );
  INV_X1 U6286 ( .A(n12463), .ZN(n12464) );
  INV_X1 U6287 ( .A(n68000), .ZN(n12465) );
  INV_X1 U6288 ( .A(n12465), .ZN(n12466) );
  BUF_X1 U6289 ( .A(n12469), .Z(n12467) );
  INV_X1 U6290 ( .A(n12471), .ZN(n12468) );
  INV_X1 U6291 ( .A(n12468), .ZN(n12469) );
  INV_X1 U6292 ( .A(n67990), .ZN(n12470) );
  INV_X1 U6293 ( .A(n12470), .ZN(n12471) );
  BUF_X1 U6294 ( .A(n12474), .Z(n12472) );
  INV_X1 U6295 ( .A(n12476), .ZN(n12473) );
  INV_X1 U6296 ( .A(n12473), .ZN(n12474) );
  INV_X1 U6297 ( .A(n67980), .ZN(n12475) );
  INV_X1 U6298 ( .A(n12475), .ZN(n12476) );
  BUF_X1 U6299 ( .A(n12479), .Z(n12477) );
  INV_X1 U6300 ( .A(n12481), .ZN(n12478) );
  INV_X1 U6301 ( .A(n12478), .ZN(n12479) );
  INV_X1 U6302 ( .A(n67970), .ZN(n12480) );
  INV_X1 U6303 ( .A(n12480), .ZN(n12481) );
  BUF_X1 U6304 ( .A(n12484), .Z(n12482) );
  INV_X1 U6305 ( .A(n12486), .ZN(n12483) );
  INV_X1 U6306 ( .A(n12483), .ZN(n12484) );
  INV_X1 U6307 ( .A(n67960), .ZN(n12485) );
  INV_X1 U6308 ( .A(n12485), .ZN(n12486) );
  BUF_X1 U6309 ( .A(n12489), .Z(n12487) );
  INV_X1 U6310 ( .A(n12491), .ZN(n12488) );
  INV_X1 U6311 ( .A(n12488), .ZN(n12489) );
  INV_X1 U6312 ( .A(n67950), .ZN(n12490) );
  INV_X1 U6313 ( .A(n12490), .ZN(n12491) );
  BUF_X1 U6314 ( .A(n12494), .Z(n12492) );
  INV_X1 U6315 ( .A(n12496), .ZN(n12493) );
  INV_X1 U6316 ( .A(n12493), .ZN(n12494) );
  INV_X1 U6317 ( .A(n67940), .ZN(n12495) );
  INV_X1 U6318 ( .A(n12495), .ZN(n12496) );
  BUF_X1 U6319 ( .A(n12499), .Z(n12497) );
  INV_X1 U6320 ( .A(n12501), .ZN(n12498) );
  INV_X1 U6321 ( .A(n12498), .ZN(n12499) );
  INV_X1 U6322 ( .A(n67930), .ZN(n12500) );
  INV_X1 U6323 ( .A(n12500), .ZN(n12501) );
  BUF_X1 U6324 ( .A(n12504), .Z(n12502) );
  INV_X1 U6325 ( .A(n12506), .ZN(n12503) );
  INV_X1 U6326 ( .A(n12503), .ZN(n12504) );
  INV_X1 U6327 ( .A(n67920), .ZN(n12505) );
  INV_X1 U6328 ( .A(n12505), .ZN(n12506) );
  BUF_X1 U6329 ( .A(n12509), .Z(n12507) );
  INV_X1 U6330 ( .A(n12511), .ZN(n12508) );
  INV_X1 U6331 ( .A(n12508), .ZN(n12509) );
  INV_X1 U6332 ( .A(n67910), .ZN(n12510) );
  INV_X1 U6333 ( .A(n12510), .ZN(n12511) );
  BUF_X1 U6334 ( .A(n12514), .Z(n12512) );
  INV_X1 U6335 ( .A(n12516), .ZN(n12513) );
  INV_X1 U6336 ( .A(n12513), .ZN(n12514) );
  INV_X1 U6337 ( .A(n67900), .ZN(n12515) );
  INV_X1 U6338 ( .A(n12515), .ZN(n12516) );
  BUF_X1 U6339 ( .A(n12519), .Z(n12517) );
  INV_X1 U6340 ( .A(n12521), .ZN(n12518) );
  INV_X1 U6341 ( .A(n12518), .ZN(n12519) );
  INV_X1 U6342 ( .A(n67890), .ZN(n12520) );
  INV_X1 U6343 ( .A(n12520), .ZN(n12521) );
  BUF_X1 U6344 ( .A(n12524), .Z(n12522) );
  INV_X1 U6345 ( .A(n12526), .ZN(n12523) );
  INV_X1 U6346 ( .A(n12523), .ZN(n12524) );
  INV_X1 U6347 ( .A(n67880), .ZN(n12525) );
  INV_X1 U6348 ( .A(n12525), .ZN(n12526) );
  BUF_X1 U6349 ( .A(n12529), .Z(n12527) );
  INV_X1 U6350 ( .A(n12531), .ZN(n12528) );
  INV_X1 U6351 ( .A(n12528), .ZN(n12529) );
  INV_X1 U6352 ( .A(n67870), .ZN(n12530) );
  INV_X1 U6353 ( .A(n12530), .ZN(n12531) );
  BUF_X1 U6354 ( .A(n12534), .Z(n12532) );
  INV_X1 U6355 ( .A(n12536), .ZN(n12533) );
  INV_X1 U6356 ( .A(n12533), .ZN(n12534) );
  INV_X1 U6357 ( .A(n67860), .ZN(n12535) );
  INV_X1 U6358 ( .A(n12535), .ZN(n12536) );
  BUF_X1 U6359 ( .A(n12539), .Z(n12537) );
  INV_X1 U6360 ( .A(n12541), .ZN(n12538) );
  INV_X1 U6361 ( .A(n12538), .ZN(n12539) );
  INV_X1 U6362 ( .A(n67850), .ZN(n12540) );
  INV_X1 U6363 ( .A(n12540), .ZN(n12541) );
  BUF_X1 U6364 ( .A(n12544), .Z(n12542) );
  INV_X1 U6365 ( .A(n12546), .ZN(n12543) );
  INV_X1 U6366 ( .A(n12543), .ZN(n12544) );
  INV_X1 U6367 ( .A(n67840), .ZN(n12545) );
  INV_X1 U6368 ( .A(n12545), .ZN(n12546) );
  BUF_X1 U6369 ( .A(n12549), .Z(n12547) );
  INV_X1 U6370 ( .A(n12551), .ZN(n12548) );
  INV_X1 U6371 ( .A(n12548), .ZN(n12549) );
  INV_X1 U6372 ( .A(n67830), .ZN(n12550) );
  INV_X1 U6373 ( .A(n12550), .ZN(n12551) );
  BUF_X1 U6374 ( .A(n12554), .Z(n12552) );
  INV_X1 U6375 ( .A(n12556), .ZN(n12553) );
  INV_X1 U6376 ( .A(n12553), .ZN(n12554) );
  INV_X1 U6377 ( .A(n67820), .ZN(n12555) );
  INV_X1 U6378 ( .A(n12555), .ZN(n12556) );
  BUF_X1 U6379 ( .A(n12559), .Z(n12557) );
  INV_X1 U6380 ( .A(n12561), .ZN(n12558) );
  INV_X1 U6381 ( .A(n12558), .ZN(n12559) );
  INV_X1 U6382 ( .A(n6781), .ZN(n12560) );
  INV_X1 U6383 ( .A(n12560), .ZN(n12561) );
  BUF_X1 U6384 ( .A(n12564), .Z(n12562) );
  INV_X1 U6385 ( .A(n12566), .ZN(n12563) );
  INV_X1 U6386 ( .A(n12563), .ZN(n12564) );
  INV_X1 U6387 ( .A(n6780), .ZN(n12565) );
  INV_X1 U6388 ( .A(n12565), .ZN(n12566) );
  BUF_X1 U6389 ( .A(n12569), .Z(n12567) );
  INV_X1 U6390 ( .A(n12571), .ZN(n12568) );
  INV_X1 U6391 ( .A(n12568), .ZN(n12569) );
  INV_X1 U6392 ( .A(n6779), .ZN(n12570) );
  INV_X1 U6393 ( .A(n12570), .ZN(n12571) );
  BUF_X1 U6394 ( .A(n12574), .Z(n12572) );
  INV_X1 U6395 ( .A(n12576), .ZN(n12573) );
  INV_X1 U6396 ( .A(n12573), .ZN(n12574) );
  INV_X1 U6397 ( .A(n6778), .ZN(n12575) );
  INV_X1 U6398 ( .A(n12575), .ZN(n12576) );
  BUF_X1 U6399 ( .A(n12579), .Z(n12577) );
  INV_X1 U6400 ( .A(n12581), .ZN(n12578) );
  INV_X1 U6401 ( .A(n12578), .ZN(n12579) );
  INV_X1 U6402 ( .A(n6777), .ZN(n12580) );
  INV_X1 U6403 ( .A(n12580), .ZN(n12581) );
  BUF_X1 U6404 ( .A(n12584), .Z(n12582) );
  INV_X1 U6405 ( .A(n12586), .ZN(n12583) );
  INV_X1 U6406 ( .A(n12583), .ZN(n12584) );
  INV_X1 U6407 ( .A(n6776), .ZN(n12585) );
  INV_X1 U6408 ( .A(n12585), .ZN(n12586) );
  BUF_X1 U6409 ( .A(n12589), .Z(n12587) );
  INV_X1 U6410 ( .A(n12591), .ZN(n12588) );
  INV_X1 U6411 ( .A(n12588), .ZN(n12589) );
  INV_X1 U6412 ( .A(n6775), .ZN(n12590) );
  INV_X1 U6413 ( .A(n12590), .ZN(n12591) );
  BUF_X1 U6414 ( .A(n12594), .Z(n12592) );
  INV_X1 U6415 ( .A(n12596), .ZN(n12593) );
  INV_X1 U6416 ( .A(n12593), .ZN(n12594) );
  INV_X1 U6417 ( .A(n6774), .ZN(n12595) );
  INV_X1 U6418 ( .A(n12595), .ZN(n12596) );
  BUF_X1 U6419 ( .A(n12599), .Z(n12597) );
  INV_X1 U6420 ( .A(n12601), .ZN(n12598) );
  INV_X1 U6421 ( .A(n12598), .ZN(n12599) );
  INV_X1 U6422 ( .A(n6773), .ZN(n12600) );
  INV_X1 U6423 ( .A(n12600), .ZN(n12601) );
  BUF_X1 U6424 ( .A(n12604), .Z(n12602) );
  INV_X1 U6425 ( .A(n12606), .ZN(n12603) );
  INV_X1 U6426 ( .A(n12603), .ZN(n12604) );
  INV_X1 U6427 ( .A(n6772), .ZN(n12605) );
  INV_X1 U6428 ( .A(n12605), .ZN(n12606) );
  BUF_X1 U6429 ( .A(n12609), .Z(n12607) );
  INV_X1 U6430 ( .A(n12611), .ZN(n12608) );
  INV_X1 U6431 ( .A(n12608), .ZN(n12609) );
  INV_X1 U6432 ( .A(n6771), .ZN(n12610) );
  INV_X1 U6433 ( .A(n12610), .ZN(n12611) );
  BUF_X1 U6434 ( .A(n12614), .Z(n12612) );
  INV_X1 U6435 ( .A(n12616), .ZN(n12613) );
  INV_X1 U6436 ( .A(n12613), .ZN(n12614) );
  INV_X1 U6437 ( .A(n6770), .ZN(n12615) );
  INV_X1 U6438 ( .A(n12615), .ZN(n12616) );
  BUF_X1 U6439 ( .A(n12619), .Z(n12617) );
  INV_X1 U6440 ( .A(n12621), .ZN(n12618) );
  INV_X1 U6441 ( .A(n12618), .ZN(n12619) );
  INV_X1 U6442 ( .A(n6769), .ZN(n12620) );
  INV_X1 U6443 ( .A(n12620), .ZN(n12621) );
  BUF_X1 U6444 ( .A(n12624), .Z(n12622) );
  INV_X1 U6445 ( .A(n12626), .ZN(n12623) );
  INV_X1 U6446 ( .A(n12623), .ZN(n12624) );
  INV_X1 U6447 ( .A(n6768), .ZN(n12625) );
  INV_X1 U6448 ( .A(n12625), .ZN(n12626) );
  BUF_X1 U6449 ( .A(n12629), .Z(n12627) );
  INV_X1 U6450 ( .A(n12631), .ZN(n12628) );
  INV_X1 U6451 ( .A(n12628), .ZN(n12629) );
  INV_X1 U6452 ( .A(n6767), .ZN(n12630) );
  INV_X1 U6453 ( .A(n12630), .ZN(n12631) );
  BUF_X1 U6454 ( .A(n12634), .Z(n12632) );
  INV_X1 U6455 ( .A(n12636), .ZN(n12633) );
  INV_X1 U6456 ( .A(n12633), .ZN(n12634) );
  INV_X1 U6457 ( .A(n6766), .ZN(n12635) );
  INV_X1 U6458 ( .A(n12635), .ZN(n12636) );
  BUF_X1 U6459 ( .A(n12639), .Z(n12637) );
  INV_X1 U6460 ( .A(n12641), .ZN(n12638) );
  INV_X1 U6461 ( .A(n12638), .ZN(n12639) );
  INV_X1 U6462 ( .A(n6765), .ZN(n12640) );
  INV_X1 U6463 ( .A(n12640), .ZN(n12641) );
  BUF_X1 U6464 ( .A(n12644), .Z(n12642) );
  INV_X1 U6465 ( .A(n12646), .ZN(n12643) );
  INV_X1 U6466 ( .A(n12643), .ZN(n12644) );
  INV_X1 U6467 ( .A(n67640), .ZN(n12645) );
  INV_X1 U6468 ( .A(n12645), .ZN(n12646) );
  BUF_X1 U6469 ( .A(n12649), .Z(n12647) );
  INV_X1 U6470 ( .A(n12651), .ZN(n12648) );
  INV_X1 U6471 ( .A(n12648), .ZN(n12649) );
  INV_X1 U6472 ( .A(n67630), .ZN(n12650) );
  INV_X1 U6473 ( .A(n12650), .ZN(n12651) );
  BUF_X1 U6474 ( .A(n12654), .Z(n12652) );
  INV_X1 U6475 ( .A(n12656), .ZN(n12653) );
  INV_X1 U6476 ( .A(n12653), .ZN(n12654) );
  INV_X1 U6477 ( .A(n67620), .ZN(n12655) );
  INV_X1 U6478 ( .A(n12655), .ZN(n12656) );
  BUF_X1 U6479 ( .A(n12659), .Z(n12657) );
  INV_X1 U6480 ( .A(n12661), .ZN(n12658) );
  INV_X1 U6481 ( .A(n12658), .ZN(n12659) );
  INV_X1 U6482 ( .A(n67610), .ZN(n12660) );
  INV_X1 U6483 ( .A(n12660), .ZN(n12661) );
  BUF_X1 U6484 ( .A(n12664), .Z(n12662) );
  INV_X1 U6485 ( .A(n12666), .ZN(n12663) );
  INV_X1 U6486 ( .A(n12663), .ZN(n12664) );
  INV_X1 U6487 ( .A(n67600), .ZN(n12665) );
  INV_X1 U6488 ( .A(n12665), .ZN(n12666) );
  BUF_X1 U6489 ( .A(n12669), .Z(n12667) );
  INV_X1 U6490 ( .A(n12671), .ZN(n12668) );
  INV_X1 U6491 ( .A(n12668), .ZN(n12669) );
  INV_X1 U6492 ( .A(n67590), .ZN(n12670) );
  INV_X1 U6493 ( .A(n12670), .ZN(n12671) );
  BUF_X1 U6494 ( .A(n12674), .Z(n12672) );
  INV_X1 U6495 ( .A(n12676), .ZN(n12673) );
  INV_X1 U6496 ( .A(n12673), .ZN(n12674) );
  INV_X1 U6497 ( .A(n67580), .ZN(n12675) );
  INV_X1 U6498 ( .A(n12675), .ZN(n12676) );
  BUF_X1 U6499 ( .A(n12679), .Z(n12677) );
  INV_X1 U6500 ( .A(n12681), .ZN(n12678) );
  INV_X1 U6501 ( .A(n12678), .ZN(n12679) );
  INV_X1 U6502 ( .A(n67570), .ZN(n12680) );
  INV_X1 U6503 ( .A(n12680), .ZN(n12681) );
  BUF_X1 U6504 ( .A(n12684), .Z(n12682) );
  INV_X1 U6505 ( .A(n12686), .ZN(n12683) );
  INV_X1 U6506 ( .A(n12683), .ZN(n12684) );
  INV_X1 U6507 ( .A(n67560), .ZN(n12685) );
  INV_X1 U6508 ( .A(n12685), .ZN(n12686) );
  BUF_X1 U6509 ( .A(n12689), .Z(n12687) );
  INV_X1 U6510 ( .A(n12691), .ZN(n12688) );
  INV_X1 U6511 ( .A(n12688), .ZN(n12689) );
  INV_X1 U6512 ( .A(n67550), .ZN(n12690) );
  INV_X1 U6513 ( .A(n12690), .ZN(n12691) );
  BUF_X1 U6514 ( .A(n12694), .Z(n12692) );
  INV_X1 U6515 ( .A(n12696), .ZN(n12693) );
  INV_X1 U6516 ( .A(n12693), .ZN(n12694) );
  INV_X1 U6517 ( .A(n67540), .ZN(n12695) );
  INV_X1 U6518 ( .A(n12695), .ZN(n12696) );
  BUF_X1 U6519 ( .A(n12699), .Z(n12697) );
  INV_X1 U6520 ( .A(n12701), .ZN(n12698) );
  INV_X1 U6521 ( .A(n12698), .ZN(n12699) );
  INV_X1 U6522 ( .A(n67530), .ZN(n12700) );
  INV_X1 U6523 ( .A(n12700), .ZN(n12701) );
  BUF_X1 U6524 ( .A(n12704), .Z(n12702) );
  INV_X1 U6525 ( .A(n12706), .ZN(n12703) );
  INV_X1 U6526 ( .A(n12703), .ZN(n12704) );
  INV_X1 U6527 ( .A(n67520), .ZN(n12705) );
  INV_X1 U6528 ( .A(n12705), .ZN(n12706) );
  BUF_X1 U6529 ( .A(n12709), .Z(n12707) );
  INV_X1 U6530 ( .A(n12711), .ZN(n12708) );
  INV_X1 U6531 ( .A(n12708), .ZN(n12709) );
  INV_X1 U6532 ( .A(n67510), .ZN(n12710) );
  INV_X1 U6533 ( .A(n12710), .ZN(n12711) );
  BUF_X1 U6534 ( .A(n12714), .Z(n12712) );
  INV_X1 U6535 ( .A(n12716), .ZN(n12713) );
  INV_X1 U6536 ( .A(n12713), .ZN(n12714) );
  INV_X1 U6537 ( .A(n67500), .ZN(n12715) );
  INV_X1 U6538 ( .A(n12715), .ZN(n12716) );
  BUF_X1 U6539 ( .A(n12719), .Z(n12717) );
  INV_X1 U6540 ( .A(n12721), .ZN(n12718) );
  INV_X1 U6541 ( .A(n12718), .ZN(n12719) );
  INV_X1 U6542 ( .A(n67490), .ZN(n12720) );
  INV_X1 U6543 ( .A(n12720), .ZN(n12721) );
  BUF_X1 U6544 ( .A(n12724), .Z(n12722) );
  INV_X1 U6545 ( .A(n12726), .ZN(n12723) );
  INV_X1 U6546 ( .A(n12723), .ZN(n12724) );
  INV_X1 U6547 ( .A(n6748), .ZN(n12725) );
  INV_X1 U6548 ( .A(n12725), .ZN(n12726) );
  BUF_X1 U6549 ( .A(n12729), .Z(n12727) );
  INV_X1 U6550 ( .A(n12731), .ZN(n12728) );
  INV_X1 U6551 ( .A(n12728), .ZN(n12729) );
  INV_X1 U6552 ( .A(n6747), .ZN(n12730) );
  INV_X1 U6553 ( .A(n12730), .ZN(n12731) );
  BUF_X1 U6554 ( .A(n12734), .Z(n12732) );
  INV_X1 U6555 ( .A(n12736), .ZN(n12733) );
  INV_X1 U6556 ( .A(n12733), .ZN(n12734) );
  INV_X1 U6557 ( .A(n6746), .ZN(n12735) );
  INV_X1 U6558 ( .A(n12735), .ZN(n12736) );
  BUF_X1 U6559 ( .A(n12739), .Z(n12737) );
  INV_X1 U6560 ( .A(n12741), .ZN(n12738) );
  INV_X1 U6561 ( .A(n12738), .ZN(n12739) );
  INV_X1 U6562 ( .A(n6745), .ZN(n12740) );
  INV_X1 U6563 ( .A(n12740), .ZN(n12741) );
  BUF_X1 U6564 ( .A(n12744), .Z(n12742) );
  INV_X1 U6565 ( .A(n12746), .ZN(n12743) );
  INV_X1 U6566 ( .A(n12743), .ZN(n12744) );
  INV_X1 U6567 ( .A(n6744), .ZN(n12745) );
  INV_X1 U6568 ( .A(n12745), .ZN(n12746) );
  BUF_X1 U6569 ( .A(n12749), .Z(n12747) );
  INV_X1 U6570 ( .A(n12751), .ZN(n12748) );
  INV_X1 U6571 ( .A(n12748), .ZN(n12749) );
  INV_X1 U6572 ( .A(n6743), .ZN(n12750) );
  INV_X1 U6573 ( .A(n12750), .ZN(n12751) );
  BUF_X1 U6574 ( .A(n12754), .Z(n12752) );
  INV_X1 U6575 ( .A(n12756), .ZN(n12753) );
  INV_X1 U6576 ( .A(n12753), .ZN(n12754) );
  INV_X1 U6577 ( .A(n6742), .ZN(n12755) );
  INV_X1 U6578 ( .A(n12755), .ZN(n12756) );
  BUF_X1 U6579 ( .A(n12759), .Z(n12757) );
  INV_X1 U6580 ( .A(n12761), .ZN(n12758) );
  INV_X1 U6581 ( .A(n12758), .ZN(n12759) );
  INV_X1 U6582 ( .A(n6741), .ZN(n12760) );
  INV_X1 U6583 ( .A(n12760), .ZN(n12761) );
  BUF_X1 U6584 ( .A(n12764), .Z(n12762) );
  INV_X1 U6585 ( .A(n12766), .ZN(n12763) );
  INV_X1 U6586 ( .A(n12763), .ZN(n12764) );
  INV_X1 U6587 ( .A(n6740), .ZN(n12765) );
  INV_X1 U6588 ( .A(n12765), .ZN(n12766) );
  BUF_X1 U6589 ( .A(n12769), .Z(n12767) );
  INV_X1 U6590 ( .A(n12771), .ZN(n12768) );
  INV_X1 U6591 ( .A(n12768), .ZN(n12769) );
  INV_X1 U6592 ( .A(n6739), .ZN(n12770) );
  INV_X1 U6593 ( .A(n12770), .ZN(n12771) );
  BUF_X1 U6594 ( .A(n12774), .Z(n12772) );
  INV_X1 U6595 ( .A(n12776), .ZN(n12773) );
  INV_X1 U6596 ( .A(n12773), .ZN(n12774) );
  INV_X1 U6597 ( .A(n6738), .ZN(n12775) );
  INV_X1 U6598 ( .A(n12775), .ZN(n12776) );
  BUF_X1 U6599 ( .A(n12779), .Z(n12777) );
  INV_X1 U6600 ( .A(n12781), .ZN(n12778) );
  INV_X1 U6601 ( .A(n12778), .ZN(n12779) );
  INV_X1 U6602 ( .A(n6737), .ZN(n12780) );
  INV_X1 U6603 ( .A(n12780), .ZN(n12781) );
  BUF_X1 U6604 ( .A(n12784), .Z(n12782) );
  INV_X1 U6605 ( .A(n12786), .ZN(n12783) );
  INV_X1 U6606 ( .A(n12783), .ZN(n12784) );
  INV_X1 U6607 ( .A(n6736), .ZN(n12785) );
  INV_X1 U6608 ( .A(n12785), .ZN(n12786) );
  BUF_X1 U6609 ( .A(n12789), .Z(n12787) );
  INV_X1 U6610 ( .A(n12791), .ZN(n12788) );
  INV_X1 U6611 ( .A(n12788), .ZN(n12789) );
  INV_X1 U6612 ( .A(n6735), .ZN(n12790) );
  INV_X1 U6613 ( .A(n12790), .ZN(n12791) );
  BUF_X1 U6614 ( .A(n12794), .Z(n12792) );
  INV_X1 U6615 ( .A(n12796), .ZN(n12793) );
  INV_X1 U6616 ( .A(n12793), .ZN(n12794) );
  INV_X1 U6617 ( .A(n6734), .ZN(n12795) );
  INV_X1 U6618 ( .A(n12795), .ZN(n12796) );
  BUF_X1 U6619 ( .A(n12799), .Z(n12797) );
  INV_X1 U6620 ( .A(n12801), .ZN(n12798) );
  INV_X1 U6621 ( .A(n12798), .ZN(n12799) );
  INV_X1 U6622 ( .A(n6733), .ZN(n12800) );
  INV_X1 U6623 ( .A(n12800), .ZN(n12801) );
  BUF_X1 U6624 ( .A(n12804), .Z(n12802) );
  INV_X1 U6625 ( .A(n12806), .ZN(n12803) );
  INV_X1 U6626 ( .A(n12803), .ZN(n12804) );
  INV_X1 U6627 ( .A(n6732), .ZN(n12805) );
  INV_X1 U6628 ( .A(n12805), .ZN(n12806) );
  BUF_X1 U6629 ( .A(n12809), .Z(n12807) );
  INV_X1 U6630 ( .A(n12811), .ZN(n12808) );
  INV_X1 U6631 ( .A(n12808), .ZN(n12809) );
  INV_X1 U6632 ( .A(n6731), .ZN(n12810) );
  INV_X1 U6633 ( .A(n12810), .ZN(n12811) );
  BUF_X1 U6634 ( .A(n12814), .Z(n12812) );
  INV_X1 U6635 ( .A(n12816), .ZN(n12813) );
  INV_X1 U6636 ( .A(n12813), .ZN(n12814) );
  INV_X1 U6637 ( .A(n6730), .ZN(n12815) );
  INV_X1 U6638 ( .A(n12815), .ZN(n12816) );
  BUF_X1 U6639 ( .A(n12819), .Z(n12817) );
  INV_X1 U6640 ( .A(n12821), .ZN(n12818) );
  INV_X1 U6641 ( .A(n12818), .ZN(n12819) );
  INV_X1 U6642 ( .A(n6729), .ZN(n12820) );
  INV_X1 U6643 ( .A(n12820), .ZN(n12821) );
  BUF_X1 U6644 ( .A(n12824), .Z(n12822) );
  INV_X1 U6645 ( .A(n12826), .ZN(n12823) );
  INV_X1 U6646 ( .A(n12823), .ZN(n12824) );
  INV_X1 U6647 ( .A(n6728), .ZN(n12825) );
  INV_X1 U6648 ( .A(n12825), .ZN(n12826) );
  BUF_X1 U6649 ( .A(n12829), .Z(n12827) );
  INV_X1 U6650 ( .A(n12831), .ZN(n12828) );
  INV_X1 U6651 ( .A(n12828), .ZN(n12829) );
  INV_X1 U6652 ( .A(n6727), .ZN(n12830) );
  INV_X1 U6653 ( .A(n12830), .ZN(n12831) );
  BUF_X1 U6654 ( .A(n12834), .Z(n12832) );
  INV_X1 U6655 ( .A(n12836), .ZN(n12833) );
  INV_X1 U6656 ( .A(n12833), .ZN(n12834) );
  INV_X1 U6657 ( .A(n6726), .ZN(n12835) );
  INV_X1 U6658 ( .A(n12835), .ZN(n12836) );
  BUF_X1 U6659 ( .A(n12839), .Z(n12837) );
  INV_X1 U6660 ( .A(n12841), .ZN(n12838) );
  INV_X1 U6661 ( .A(n12838), .ZN(n12839) );
  INV_X1 U6662 ( .A(n6725), .ZN(n12840) );
  INV_X1 U6663 ( .A(n12840), .ZN(n12841) );
  BUF_X1 U6664 ( .A(n12844), .Z(n12842) );
  INV_X1 U6665 ( .A(n12846), .ZN(n12843) );
  INV_X1 U6666 ( .A(n12843), .ZN(n12844) );
  INV_X1 U6667 ( .A(n6724), .ZN(n12845) );
  INV_X1 U6668 ( .A(n12845), .ZN(n12846) );
  BUF_X1 U6669 ( .A(n12849), .Z(n12847) );
  INV_X1 U6670 ( .A(n12851), .ZN(n12848) );
  INV_X1 U6671 ( .A(n12848), .ZN(n12849) );
  INV_X1 U6672 ( .A(n6723), .ZN(n12850) );
  INV_X1 U6673 ( .A(n12850), .ZN(n12851) );
  BUF_X1 U6674 ( .A(n12854), .Z(n12852) );
  INV_X1 U6675 ( .A(n12856), .ZN(n12853) );
  INV_X1 U6676 ( .A(n12853), .ZN(n12854) );
  INV_X1 U6677 ( .A(n6722), .ZN(n12855) );
  INV_X1 U6678 ( .A(n12855), .ZN(n12856) );
  BUF_X1 U6679 ( .A(n12859), .Z(n12857) );
  INV_X1 U6680 ( .A(n12861), .ZN(n12858) );
  INV_X1 U6681 ( .A(n12858), .ZN(n12859) );
  INV_X1 U6682 ( .A(n6721), .ZN(n12860) );
  INV_X1 U6683 ( .A(n12860), .ZN(n12861) );
  BUF_X1 U6684 ( .A(n12864), .Z(n12862) );
  INV_X1 U6685 ( .A(n12866), .ZN(n12863) );
  INV_X1 U6686 ( .A(n12863), .ZN(n12864) );
  INV_X1 U6687 ( .A(n67200), .ZN(n12865) );
  INV_X1 U6688 ( .A(n12865), .ZN(n12866) );
  BUF_X1 U6689 ( .A(n12869), .Z(n12867) );
  INV_X1 U6690 ( .A(n12871), .ZN(n12868) );
  INV_X1 U6691 ( .A(n12868), .ZN(n12869) );
  INV_X1 U6692 ( .A(n67190), .ZN(n12870) );
  INV_X1 U6693 ( .A(n12870), .ZN(n12871) );
  BUF_X1 U6694 ( .A(n12874), .Z(n12872) );
  INV_X1 U6695 ( .A(n12876), .ZN(n12873) );
  INV_X1 U6696 ( .A(n12873), .ZN(n12874) );
  INV_X1 U6697 ( .A(n67180), .ZN(n12875) );
  INV_X1 U6698 ( .A(n12875), .ZN(n12876) );
  BUF_X1 U6699 ( .A(n12879), .Z(n12877) );
  INV_X1 U6700 ( .A(n12881), .ZN(n12878) );
  INV_X1 U6701 ( .A(n12878), .ZN(n12879) );
  INV_X1 U6702 ( .A(n67170), .ZN(n12880) );
  INV_X1 U6703 ( .A(n12880), .ZN(n12881) );
  BUF_X1 U6704 ( .A(n12884), .Z(n12882) );
  INV_X1 U6705 ( .A(n12886), .ZN(n12883) );
  INV_X1 U6706 ( .A(n12883), .ZN(n12884) );
  INV_X1 U6707 ( .A(n67160), .ZN(n12885) );
  INV_X1 U6708 ( .A(n12885), .ZN(n12886) );
  BUF_X1 U6709 ( .A(n12889), .Z(n12887) );
  INV_X1 U6710 ( .A(n12891), .ZN(n12888) );
  INV_X1 U6711 ( .A(n12888), .ZN(n12889) );
  INV_X1 U6712 ( .A(n67150), .ZN(n12890) );
  INV_X1 U6713 ( .A(n12890), .ZN(n12891) );
  BUF_X1 U6714 ( .A(n12894), .Z(n12892) );
  INV_X1 U6715 ( .A(n12896), .ZN(n12893) );
  INV_X1 U6716 ( .A(n12893), .ZN(n12894) );
  INV_X1 U6717 ( .A(n67140), .ZN(n12895) );
  INV_X1 U6718 ( .A(n12895), .ZN(n12896) );
  BUF_X1 U6719 ( .A(n12899), .Z(n12897) );
  INV_X1 U6720 ( .A(n12901), .ZN(n12898) );
  INV_X1 U6721 ( .A(n12898), .ZN(n12899) );
  INV_X1 U6722 ( .A(n67130), .ZN(n12900) );
  INV_X1 U6723 ( .A(n12900), .ZN(n12901) );
  BUF_X1 U6724 ( .A(n12904), .Z(n12902) );
  INV_X1 U6725 ( .A(n12906), .ZN(n12903) );
  INV_X1 U6726 ( .A(n12903), .ZN(n12904) );
  INV_X1 U6727 ( .A(n67120), .ZN(n12905) );
  INV_X1 U6728 ( .A(n12905), .ZN(n12906) );
  BUF_X1 U6729 ( .A(n12909), .Z(n12907) );
  INV_X1 U6730 ( .A(n12911), .ZN(n12908) );
  INV_X1 U6731 ( .A(n12908), .ZN(n12909) );
  INV_X1 U6732 ( .A(n67110), .ZN(n12910) );
  INV_X1 U6733 ( .A(n12910), .ZN(n12911) );
  BUF_X1 U6734 ( .A(n12914), .Z(n12912) );
  INV_X1 U6735 ( .A(n12916), .ZN(n12913) );
  INV_X1 U6736 ( .A(n12913), .ZN(n12914) );
  INV_X1 U6737 ( .A(n67100), .ZN(n12915) );
  INV_X1 U6738 ( .A(n12915), .ZN(n12916) );
  BUF_X1 U6739 ( .A(n12919), .Z(n12917) );
  INV_X1 U6740 ( .A(n12921), .ZN(n12918) );
  INV_X1 U6741 ( .A(n12918), .ZN(n12919) );
  INV_X1 U6742 ( .A(n67090), .ZN(n12920) );
  INV_X1 U6743 ( .A(n12920), .ZN(n12921) );
  BUF_X1 U6744 ( .A(n12924), .Z(n12922) );
  INV_X1 U6745 ( .A(n12926), .ZN(n12923) );
  INV_X1 U6746 ( .A(n12923), .ZN(n12924) );
  INV_X1 U6747 ( .A(n67080), .ZN(n12925) );
  INV_X1 U6748 ( .A(n12925), .ZN(n12926) );
  BUF_X1 U6749 ( .A(n12929), .Z(n12927) );
  INV_X1 U6750 ( .A(n12931), .ZN(n12928) );
  INV_X1 U6751 ( .A(n12928), .ZN(n12929) );
  INV_X1 U6752 ( .A(n67070), .ZN(n12930) );
  INV_X1 U6753 ( .A(n12930), .ZN(n12931) );
  BUF_X1 U6754 ( .A(n12934), .Z(n12932) );
  INV_X1 U6755 ( .A(n12936), .ZN(n12933) );
  INV_X1 U6756 ( .A(n12933), .ZN(n12934) );
  INV_X1 U6757 ( .A(n67060), .ZN(n12935) );
  INV_X1 U6758 ( .A(n12935), .ZN(n12936) );
  BUF_X1 U6759 ( .A(n12939), .Z(n12937) );
  INV_X1 U6760 ( .A(n12941), .ZN(n12938) );
  INV_X1 U6761 ( .A(n12938), .ZN(n12939) );
  INV_X1 U6762 ( .A(n67050), .ZN(n12940) );
  INV_X1 U6763 ( .A(n12940), .ZN(n12941) );
  BUF_X1 U6764 ( .A(n12944), .Z(n12942) );
  INV_X1 U6765 ( .A(n12946), .ZN(n12943) );
  INV_X1 U6766 ( .A(n12943), .ZN(n12944) );
  INV_X1 U6767 ( .A(n67040), .ZN(n12945) );
  INV_X1 U6768 ( .A(n12945), .ZN(n12946) );
  BUF_X1 U6769 ( .A(n12949), .Z(n12947) );
  INV_X1 U6770 ( .A(n12951), .ZN(n12948) );
  INV_X1 U6771 ( .A(n12948), .ZN(n12949) );
  INV_X1 U6772 ( .A(n67030), .ZN(n12950) );
  INV_X1 U6773 ( .A(n12950), .ZN(n12951) );
  BUF_X1 U6774 ( .A(n12954), .Z(n12952) );
  INV_X1 U6775 ( .A(n12956), .ZN(n12953) );
  INV_X1 U6776 ( .A(n12953), .ZN(n12954) );
  INV_X1 U6777 ( .A(n67020), .ZN(n12955) );
  INV_X1 U6778 ( .A(n12955), .ZN(n12956) );
  BUF_X1 U6779 ( .A(n12959), .Z(n12957) );
  INV_X1 U6780 ( .A(n12961), .ZN(n12958) );
  INV_X1 U6781 ( .A(n12958), .ZN(n12959) );
  INV_X1 U6782 ( .A(n67010), .ZN(n12960) );
  INV_X1 U6783 ( .A(n12960), .ZN(n12961) );
  BUF_X1 U6784 ( .A(n12964), .Z(n12962) );
  INV_X1 U6785 ( .A(n12966), .ZN(n12963) );
  INV_X1 U6786 ( .A(n12963), .ZN(n12964) );
  INV_X1 U6787 ( .A(n67000), .ZN(n12965) );
  INV_X1 U6788 ( .A(n12965), .ZN(n12966) );
  BUF_X1 U6789 ( .A(n12969), .Z(n12967) );
  INV_X1 U6790 ( .A(n12971), .ZN(n12968) );
  INV_X1 U6791 ( .A(n12968), .ZN(n12969) );
  INV_X1 U6792 ( .A(n6699), .ZN(n12970) );
  INV_X1 U6793 ( .A(n12970), .ZN(n12971) );
  BUF_X1 U6794 ( .A(n12974), .Z(n12972) );
  INV_X1 U6795 ( .A(n12976), .ZN(n12973) );
  INV_X1 U6796 ( .A(n12973), .ZN(n12974) );
  INV_X1 U6797 ( .A(n6698), .ZN(n12975) );
  INV_X1 U6798 ( .A(n12975), .ZN(n12976) );
  BUF_X1 U6799 ( .A(n12979), .Z(n12977) );
  INV_X1 U6800 ( .A(n12981), .ZN(n12978) );
  INV_X1 U6801 ( .A(n12978), .ZN(n12979) );
  INV_X1 U6802 ( .A(n6697), .ZN(n12980) );
  INV_X1 U6803 ( .A(n12980), .ZN(n12981) );
  BUF_X1 U6804 ( .A(n12984), .Z(n12982) );
  INV_X1 U6805 ( .A(n12986), .ZN(n12983) );
  INV_X1 U6806 ( .A(n12983), .ZN(n12984) );
  INV_X1 U6807 ( .A(n6696), .ZN(n12985) );
  INV_X1 U6808 ( .A(n12985), .ZN(n12986) );
  BUF_X1 U6809 ( .A(n12989), .Z(n12987) );
  INV_X1 U6810 ( .A(n12991), .ZN(n12988) );
  INV_X1 U6811 ( .A(n12988), .ZN(n12989) );
  INV_X1 U6812 ( .A(n6695), .ZN(n12990) );
  INV_X1 U6813 ( .A(n12990), .ZN(n12991) );
  BUF_X1 U6814 ( .A(n12994), .Z(n12992) );
  INV_X1 U6815 ( .A(n12996), .ZN(n12993) );
  INV_X1 U6816 ( .A(n12993), .ZN(n12994) );
  INV_X1 U6817 ( .A(n6694), .ZN(n12995) );
  INV_X1 U6818 ( .A(n12995), .ZN(n12996) );
  BUF_X1 U6819 ( .A(n12999), .Z(n12997) );
  INV_X1 U6820 ( .A(n13001), .ZN(n12998) );
  INV_X1 U6821 ( .A(n12998), .ZN(n12999) );
  INV_X1 U6822 ( .A(n6693), .ZN(n13000) );
  INV_X1 U6823 ( .A(n13000), .ZN(n13001) );
  BUF_X1 U6824 ( .A(n13004), .Z(n13002) );
  INV_X1 U6825 ( .A(n13006), .ZN(n13003) );
  INV_X1 U6826 ( .A(n13003), .ZN(n13004) );
  INV_X1 U6827 ( .A(n6692), .ZN(n13005) );
  INV_X1 U6828 ( .A(n13005), .ZN(n13006) );
  BUF_X1 U6829 ( .A(n13009), .Z(n13007) );
  INV_X1 U6830 ( .A(n13011), .ZN(n13008) );
  INV_X1 U6831 ( .A(n13008), .ZN(n13009) );
  INV_X1 U6832 ( .A(n6691), .ZN(n13010) );
  INV_X1 U6833 ( .A(n13010), .ZN(n13011) );
  BUF_X1 U6834 ( .A(n13014), .Z(n13012) );
  INV_X1 U6835 ( .A(n13016), .ZN(n13013) );
  INV_X1 U6836 ( .A(n13013), .ZN(n13014) );
  INV_X1 U6837 ( .A(n6690), .ZN(n13015) );
  INV_X1 U6838 ( .A(n13015), .ZN(n13016) );
  BUF_X1 U6839 ( .A(n13019), .Z(n13017) );
  INV_X1 U6840 ( .A(n13021), .ZN(n13018) );
  INV_X1 U6841 ( .A(n13018), .ZN(n13019) );
  INV_X1 U6842 ( .A(n6689), .ZN(n13020) );
  INV_X1 U6843 ( .A(n13020), .ZN(n13021) );
  BUF_X1 U6844 ( .A(n13024), .Z(n13022) );
  INV_X1 U6845 ( .A(n13026), .ZN(n13023) );
  INV_X1 U6846 ( .A(n13023), .ZN(n13024) );
  INV_X1 U6847 ( .A(n6688), .ZN(n13025) );
  INV_X1 U6848 ( .A(n13025), .ZN(n13026) );
  BUF_X1 U6849 ( .A(n13029), .Z(n13027) );
  INV_X1 U6850 ( .A(n13031), .ZN(n13028) );
  INV_X1 U6851 ( .A(n13028), .ZN(n13029) );
  INV_X1 U6852 ( .A(n6687), .ZN(n13030) );
  INV_X1 U6853 ( .A(n13030), .ZN(n13031) );
  BUF_X1 U6854 ( .A(n13034), .Z(n13032) );
  INV_X1 U6855 ( .A(n13036), .ZN(n13033) );
  INV_X1 U6856 ( .A(n13033), .ZN(n13034) );
  INV_X1 U6857 ( .A(n6686), .ZN(n13035) );
  INV_X1 U6858 ( .A(n13035), .ZN(n13036) );
  BUF_X1 U6859 ( .A(n13039), .Z(n13037) );
  INV_X1 U6860 ( .A(n13041), .ZN(n13038) );
  INV_X1 U6861 ( .A(n13038), .ZN(n13039) );
  INV_X1 U6862 ( .A(n6685), .ZN(n13040) );
  INV_X1 U6863 ( .A(n13040), .ZN(n13041) );
  BUF_X1 U6864 ( .A(n13044), .Z(n13042) );
  INV_X1 U6865 ( .A(n13046), .ZN(n13043) );
  INV_X1 U6866 ( .A(n13043), .ZN(n13044) );
  INV_X1 U6867 ( .A(n6684), .ZN(n13045) );
  INV_X1 U6868 ( .A(n13045), .ZN(n13046) );
  BUF_X1 U6869 ( .A(n13049), .Z(n13047) );
  INV_X1 U6870 ( .A(n13051), .ZN(n13048) );
  INV_X1 U6871 ( .A(n13048), .ZN(n13049) );
  INV_X1 U6872 ( .A(n6683), .ZN(n13050) );
  INV_X1 U6873 ( .A(n13050), .ZN(n13051) );
  BUF_X1 U6874 ( .A(n13054), .Z(n13052) );
  INV_X1 U6875 ( .A(n13056), .ZN(n13053) );
  INV_X1 U6876 ( .A(n13053), .ZN(n13054) );
  INV_X1 U6877 ( .A(n66820), .ZN(n13055) );
  INV_X1 U6878 ( .A(n13055), .ZN(n13056) );
  BUF_X1 U6879 ( .A(n13059), .Z(n13057) );
  INV_X1 U6880 ( .A(n13061), .ZN(n13058) );
  INV_X1 U6881 ( .A(n13058), .ZN(n13059) );
  INV_X1 U6882 ( .A(n66810), .ZN(n13060) );
  INV_X1 U6883 ( .A(n13060), .ZN(n13061) );
  BUF_X1 U6884 ( .A(n13064), .Z(n13062) );
  INV_X1 U6885 ( .A(n13066), .ZN(n13063) );
  INV_X1 U6886 ( .A(n13063), .ZN(n13064) );
  INV_X1 U6887 ( .A(n66800), .ZN(n13065) );
  INV_X1 U6888 ( .A(n13065), .ZN(n13066) );
  BUF_X1 U6889 ( .A(n13069), .Z(n13067) );
  INV_X1 U6890 ( .A(n13071), .ZN(n13068) );
  INV_X1 U6891 ( .A(n13068), .ZN(n13069) );
  INV_X1 U6892 ( .A(n66790), .ZN(n13070) );
  INV_X1 U6893 ( .A(n13070), .ZN(n13071) );
  BUF_X1 U6894 ( .A(n13074), .Z(n13072) );
  INV_X1 U6895 ( .A(n13076), .ZN(n13073) );
  INV_X1 U6896 ( .A(n13073), .ZN(n13074) );
  INV_X1 U6897 ( .A(n66780), .ZN(n13075) );
  INV_X1 U6898 ( .A(n13075), .ZN(n13076) );
  BUF_X1 U6899 ( .A(n13079), .Z(n13077) );
  INV_X1 U6900 ( .A(n13081), .ZN(n13078) );
  INV_X1 U6901 ( .A(n13078), .ZN(n13079) );
  INV_X1 U6902 ( .A(n66770), .ZN(n13080) );
  INV_X1 U6903 ( .A(n13080), .ZN(n13081) );
  BUF_X1 U6904 ( .A(n13084), .Z(n13082) );
  INV_X1 U6905 ( .A(n13086), .ZN(n13083) );
  INV_X1 U6906 ( .A(n13083), .ZN(n13084) );
  INV_X1 U6907 ( .A(n66760), .ZN(n13085) );
  INV_X1 U6908 ( .A(n13085), .ZN(n13086) );
  BUF_X1 U6909 ( .A(n13089), .Z(n13087) );
  INV_X1 U6910 ( .A(n13091), .ZN(n13088) );
  INV_X1 U6911 ( .A(n13088), .ZN(n13089) );
  INV_X1 U6912 ( .A(n66750), .ZN(n13090) );
  INV_X1 U6913 ( .A(n13090), .ZN(n13091) );
  BUF_X1 U6914 ( .A(n13094), .Z(n13092) );
  INV_X1 U6915 ( .A(n13096), .ZN(n13093) );
  INV_X1 U6916 ( .A(n13093), .ZN(n13094) );
  INV_X1 U6917 ( .A(n66740), .ZN(n13095) );
  INV_X1 U6918 ( .A(n13095), .ZN(n13096) );
  BUF_X1 U6919 ( .A(n13099), .Z(n13097) );
  INV_X1 U6920 ( .A(n13101), .ZN(n13098) );
  INV_X1 U6921 ( .A(n13098), .ZN(n13099) );
  INV_X1 U6922 ( .A(n66730), .ZN(n13100) );
  INV_X1 U6923 ( .A(n13100), .ZN(n13101) );
  BUF_X1 U6924 ( .A(n13104), .Z(n13102) );
  INV_X1 U6925 ( .A(n13106), .ZN(n13103) );
  INV_X1 U6926 ( .A(n13103), .ZN(n13104) );
  INV_X1 U6927 ( .A(n66720), .ZN(n13105) );
  INV_X1 U6928 ( .A(n13105), .ZN(n13106) );
  BUF_X1 U6929 ( .A(n13109), .Z(n13107) );
  INV_X1 U6930 ( .A(n13111), .ZN(n13108) );
  INV_X1 U6931 ( .A(n13108), .ZN(n13109) );
  INV_X1 U6932 ( .A(n66710), .ZN(n13110) );
  INV_X1 U6933 ( .A(n13110), .ZN(n13111) );
  BUF_X1 U6934 ( .A(n13114), .Z(n13112) );
  INV_X1 U6935 ( .A(n13116), .ZN(n13113) );
  INV_X1 U6936 ( .A(n13113), .ZN(n13114) );
  INV_X1 U6937 ( .A(n66700), .ZN(n13115) );
  INV_X1 U6938 ( .A(n13115), .ZN(n13116) );
  BUF_X1 U6939 ( .A(n13119), .Z(n13117) );
  INV_X1 U6940 ( .A(n13121), .ZN(n13118) );
  INV_X1 U6941 ( .A(n13118), .ZN(n13119) );
  INV_X1 U6942 ( .A(n66690), .ZN(n13120) );
  INV_X1 U6943 ( .A(n13120), .ZN(n13121) );
  BUF_X1 U6944 ( .A(n13124), .Z(n13122) );
  INV_X1 U6945 ( .A(n13126), .ZN(n13123) );
  INV_X1 U6946 ( .A(n13123), .ZN(n13124) );
  INV_X1 U6947 ( .A(n66680), .ZN(n13125) );
  INV_X1 U6948 ( .A(n13125), .ZN(n13126) );
  BUF_X1 U6949 ( .A(n13129), .Z(n13127) );
  INV_X1 U6950 ( .A(n13131), .ZN(n13128) );
  INV_X1 U6951 ( .A(n13128), .ZN(n13129) );
  INV_X1 U6952 ( .A(n66670), .ZN(n13130) );
  INV_X1 U6953 ( .A(n13130), .ZN(n13131) );
  BUF_X1 U6954 ( .A(n13134), .Z(n13132) );
  INV_X1 U6955 ( .A(n13136), .ZN(n13133) );
  INV_X1 U6956 ( .A(n13133), .ZN(n13134) );
  INV_X1 U6957 ( .A(n6666), .ZN(n13135) );
  INV_X1 U6958 ( .A(n13135), .ZN(n13136) );
  BUF_X1 U6959 ( .A(n13139), .Z(n13137) );
  INV_X1 U6960 ( .A(n13141), .ZN(n13138) );
  INV_X1 U6961 ( .A(n13138), .ZN(n13139) );
  INV_X1 U6962 ( .A(n6665), .ZN(n13140) );
  INV_X1 U6963 ( .A(n13140), .ZN(n13141) );
  BUF_X1 U6964 ( .A(n13144), .Z(n13142) );
  INV_X1 U6965 ( .A(n13146), .ZN(n13143) );
  INV_X1 U6966 ( .A(n13143), .ZN(n13144) );
  INV_X1 U6967 ( .A(n6664), .ZN(n13145) );
  INV_X1 U6968 ( .A(n13145), .ZN(n13146) );
  BUF_X1 U6969 ( .A(n13149), .Z(n13147) );
  INV_X1 U6970 ( .A(n13151), .ZN(n13148) );
  INV_X1 U6971 ( .A(n13148), .ZN(n13149) );
  INV_X1 U6972 ( .A(n6663), .ZN(n13150) );
  INV_X1 U6973 ( .A(n13150), .ZN(n13151) );
  BUF_X1 U6974 ( .A(n13154), .Z(n13152) );
  INV_X1 U6975 ( .A(n13156), .ZN(n13153) );
  INV_X1 U6976 ( .A(n13153), .ZN(n13154) );
  INV_X1 U6977 ( .A(n6662), .ZN(n13155) );
  INV_X1 U6978 ( .A(n13155), .ZN(n13156) );
  BUF_X1 U6979 ( .A(n13159), .Z(n13157) );
  INV_X1 U6980 ( .A(n13161), .ZN(n13158) );
  INV_X1 U6981 ( .A(n13158), .ZN(n13159) );
  INV_X1 U6982 ( .A(n6661), .ZN(n13160) );
  INV_X1 U6983 ( .A(n13160), .ZN(n13161) );
  BUF_X1 U6984 ( .A(n13164), .Z(n13162) );
  INV_X1 U6985 ( .A(n13166), .ZN(n13163) );
  INV_X1 U6986 ( .A(n13163), .ZN(n13164) );
  INV_X1 U6987 ( .A(n6660), .ZN(n13165) );
  INV_X1 U6988 ( .A(n13165), .ZN(n13166) );
  BUF_X1 U6989 ( .A(n13169), .Z(n13167) );
  INV_X1 U6990 ( .A(n13171), .ZN(n13168) );
  INV_X1 U6991 ( .A(n13168), .ZN(n13169) );
  INV_X1 U6992 ( .A(n6659), .ZN(n13170) );
  INV_X1 U6993 ( .A(n13170), .ZN(n13171) );
  BUF_X1 U6994 ( .A(n13174), .Z(n13172) );
  INV_X1 U6995 ( .A(n13176), .ZN(n13173) );
  INV_X1 U6996 ( .A(n13173), .ZN(n13174) );
  INV_X1 U6997 ( .A(n6658), .ZN(n13175) );
  INV_X1 U6998 ( .A(n13175), .ZN(n13176) );
  BUF_X1 U6999 ( .A(n13179), .Z(n13177) );
  INV_X1 U7000 ( .A(n13181), .ZN(n13178) );
  INV_X1 U7001 ( .A(n13178), .ZN(n13179) );
  INV_X1 U7002 ( .A(n6657), .ZN(n13180) );
  INV_X1 U7003 ( .A(n13180), .ZN(n13181) );
  BUF_X1 U7004 ( .A(n13184), .Z(n13182) );
  INV_X1 U7005 ( .A(n13186), .ZN(n13183) );
  INV_X1 U7006 ( .A(n13183), .ZN(n13184) );
  INV_X1 U7007 ( .A(n6656), .ZN(n13185) );
  INV_X1 U7008 ( .A(n13185), .ZN(n13186) );
  BUF_X1 U7009 ( .A(n13189), .Z(n13187) );
  INV_X1 U7010 ( .A(n13191), .ZN(n13188) );
  INV_X1 U7011 ( .A(n13188), .ZN(n13189) );
  INV_X1 U7012 ( .A(n6655), .ZN(n13190) );
  INV_X1 U7013 ( .A(n13190), .ZN(n13191) );
  BUF_X1 U7014 ( .A(n13194), .Z(n13192) );
  INV_X1 U7015 ( .A(n13196), .ZN(n13193) );
  INV_X1 U7016 ( .A(n13193), .ZN(n13194) );
  INV_X1 U7017 ( .A(n6654), .ZN(n13195) );
  INV_X1 U7018 ( .A(n13195), .ZN(n13196) );
  BUF_X1 U7019 ( .A(n13199), .Z(n13197) );
  INV_X1 U7020 ( .A(n13201), .ZN(n13198) );
  INV_X1 U7021 ( .A(n13198), .ZN(n13199) );
  INV_X1 U7022 ( .A(n6653), .ZN(n13200) );
  INV_X1 U7023 ( .A(n13200), .ZN(n13201) );
  BUF_X1 U7024 ( .A(n13204), .Z(n13202) );
  INV_X1 U7025 ( .A(n13206), .ZN(n13203) );
  INV_X1 U7026 ( .A(n13203), .ZN(n13204) );
  INV_X1 U7027 ( .A(n6652), .ZN(n13205) );
  INV_X1 U7028 ( .A(n13205), .ZN(n13206) );
  BUF_X1 U7029 ( .A(n13209), .Z(n13207) );
  INV_X1 U7030 ( .A(n13211), .ZN(n13208) );
  INV_X1 U7031 ( .A(n13208), .ZN(n13209) );
  INV_X1 U7032 ( .A(n6651), .ZN(n13210) );
  INV_X1 U7033 ( .A(n13210), .ZN(n13211) );
  BUF_X1 U7034 ( .A(n13214), .Z(n13212) );
  INV_X1 U7035 ( .A(n13216), .ZN(n13213) );
  INV_X1 U7036 ( .A(n13213), .ZN(n13214) );
  INV_X1 U7037 ( .A(n6650), .ZN(n13215) );
  INV_X1 U7038 ( .A(n13215), .ZN(n13216) );
  BUF_X1 U7039 ( .A(n13219), .Z(n13217) );
  INV_X1 U7040 ( .A(n13221), .ZN(n13218) );
  INV_X1 U7041 ( .A(n13218), .ZN(n13219) );
  INV_X1 U7042 ( .A(n6649), .ZN(n13220) );
  INV_X1 U7043 ( .A(n13220), .ZN(n13221) );
  BUF_X1 U7044 ( .A(n13224), .Z(n13222) );
  INV_X1 U7045 ( .A(n13226), .ZN(n13223) );
  INV_X1 U7046 ( .A(n13223), .ZN(n13224) );
  INV_X1 U7047 ( .A(n6648), .ZN(n13225) );
  INV_X1 U7048 ( .A(n13225), .ZN(n13226) );
  BUF_X1 U7049 ( .A(n13229), .Z(n13227) );
  INV_X1 U7050 ( .A(n13231), .ZN(n13228) );
  INV_X1 U7051 ( .A(n13228), .ZN(n13229) );
  INV_X1 U7052 ( .A(n6647), .ZN(n13230) );
  INV_X1 U7053 ( .A(n13230), .ZN(n13231) );
  BUF_X1 U7054 ( .A(n13234), .Z(n13232) );
  INV_X1 U7055 ( .A(n13236), .ZN(n13233) );
  INV_X1 U7056 ( .A(n13233), .ZN(n13234) );
  INV_X1 U7057 ( .A(n6646), .ZN(n13235) );
  INV_X1 U7058 ( .A(n13235), .ZN(n13236) );
  BUF_X1 U7059 ( .A(n13239), .Z(n13237) );
  INV_X1 U7060 ( .A(n13241), .ZN(n13238) );
  INV_X1 U7061 ( .A(n13238), .ZN(n13239) );
  INV_X1 U7062 ( .A(n6645), .ZN(n13240) );
  INV_X1 U7063 ( .A(n13240), .ZN(n13241) );
  BUF_X1 U7064 ( .A(n13244), .Z(n13242) );
  INV_X1 U7065 ( .A(n13246), .ZN(n13243) );
  INV_X1 U7066 ( .A(n13243), .ZN(n13244) );
  INV_X1 U7067 ( .A(n6644), .ZN(n13245) );
  INV_X1 U7068 ( .A(n13245), .ZN(n13246) );
  BUF_X1 U7069 ( .A(n13249), .Z(n13247) );
  INV_X1 U7070 ( .A(n13251), .ZN(n13248) );
  INV_X1 U7071 ( .A(n13248), .ZN(n13249) );
  INV_X1 U7072 ( .A(n6643), .ZN(n13250) );
  INV_X1 U7073 ( .A(n13250), .ZN(n13251) );
  BUF_X1 U7074 ( .A(n13254), .Z(n13252) );
  INV_X1 U7075 ( .A(n13256), .ZN(n13253) );
  INV_X1 U7076 ( .A(n13253), .ZN(n13254) );
  INV_X1 U7077 ( .A(n6642), .ZN(n13255) );
  INV_X1 U7078 ( .A(n13255), .ZN(n13256) );
  BUF_X1 U7079 ( .A(n13259), .Z(n13257) );
  INV_X1 U7080 ( .A(n13261), .ZN(n13258) );
  INV_X1 U7081 ( .A(n13258), .ZN(n13259) );
  INV_X1 U7082 ( .A(n6641), .ZN(n13260) );
  INV_X1 U7083 ( .A(n13260), .ZN(n13261) );
  BUF_X1 U7084 ( .A(n13264), .Z(n13262) );
  INV_X1 U7085 ( .A(n13266), .ZN(n13263) );
  INV_X1 U7086 ( .A(n13263), .ZN(n13264) );
  INV_X1 U7087 ( .A(n6640), .ZN(n13265) );
  INV_X1 U7088 ( .A(n13265), .ZN(n13266) );
  BUF_X1 U7089 ( .A(n13269), .Z(n13267) );
  INV_X1 U7090 ( .A(n13271), .ZN(n13268) );
  INV_X1 U7091 ( .A(n13268), .ZN(n13269) );
  INV_X1 U7092 ( .A(n6639), .ZN(n13270) );
  INV_X1 U7093 ( .A(n13270), .ZN(n13271) );
  BUF_X1 U7094 ( .A(n13274), .Z(n13272) );
  INV_X1 U7095 ( .A(n13276), .ZN(n13273) );
  INV_X1 U7096 ( .A(n13273), .ZN(n13274) );
  INV_X1 U7097 ( .A(n6638), .ZN(n13275) );
  INV_X1 U7098 ( .A(n13275), .ZN(n13276) );
  BUF_X1 U7099 ( .A(n13279), .Z(n13277) );
  INV_X1 U7100 ( .A(n13281), .ZN(n13278) );
  INV_X1 U7101 ( .A(n13278), .ZN(n13279) );
  INV_X1 U7102 ( .A(n6637), .ZN(n13280) );
  INV_X1 U7103 ( .A(n13280), .ZN(n13281) );
  BUF_X1 U7104 ( .A(n13284), .Z(n13282) );
  INV_X1 U7105 ( .A(n13286), .ZN(n13283) );
  INV_X1 U7106 ( .A(n13283), .ZN(n13284) );
  INV_X1 U7107 ( .A(n6636), .ZN(n13285) );
  INV_X1 U7108 ( .A(n13285), .ZN(n13286) );
  BUF_X1 U7109 ( .A(n13289), .Z(n13287) );
  INV_X1 U7110 ( .A(n13291), .ZN(n13288) );
  INV_X1 U7111 ( .A(n13288), .ZN(n13289) );
  INV_X1 U7112 ( .A(n6635), .ZN(n13290) );
  INV_X1 U7113 ( .A(n13290), .ZN(n13291) );
  BUF_X1 U7114 ( .A(n13294), .Z(n13292) );
  INV_X1 U7115 ( .A(n13296), .ZN(n13293) );
  INV_X1 U7116 ( .A(n13293), .ZN(n13294) );
  INV_X1 U7117 ( .A(n6634), .ZN(n13295) );
  INV_X1 U7118 ( .A(n13295), .ZN(n13296) );
  BUF_X1 U7119 ( .A(n13299), .Z(n13297) );
  INV_X1 U7120 ( .A(n13301), .ZN(n13298) );
  INV_X1 U7121 ( .A(n13298), .ZN(n13299) );
  INV_X1 U7122 ( .A(n6633), .ZN(n13300) );
  INV_X1 U7123 ( .A(n13300), .ZN(n13301) );
  BUF_X1 U7124 ( .A(n13304), .Z(n13302) );
  INV_X1 U7125 ( .A(n13306), .ZN(n13303) );
  INV_X1 U7126 ( .A(n13303), .ZN(n13304) );
  INV_X1 U7127 ( .A(n6632), .ZN(n13305) );
  INV_X1 U7128 ( .A(n13305), .ZN(n13306) );
  BUF_X1 U7129 ( .A(n13309), .Z(n13307) );
  INV_X1 U7130 ( .A(n13311), .ZN(n13308) );
  INV_X1 U7131 ( .A(n13308), .ZN(n13309) );
  INV_X1 U7132 ( .A(n6631), .ZN(n13310) );
  INV_X1 U7133 ( .A(n13310), .ZN(n13311) );
  BUF_X1 U7134 ( .A(n13314), .Z(n13312) );
  INV_X1 U7135 ( .A(n13316), .ZN(n13313) );
  INV_X1 U7136 ( .A(n13313), .ZN(n13314) );
  INV_X1 U7137 ( .A(n6630), .ZN(n13315) );
  INV_X1 U7138 ( .A(n13315), .ZN(n13316) );
  BUF_X1 U7139 ( .A(n13319), .Z(n13317) );
  INV_X1 U7140 ( .A(n13321), .ZN(n13318) );
  INV_X1 U7141 ( .A(n13318), .ZN(n13319) );
  INV_X1 U7142 ( .A(n6629), .ZN(n13320) );
  INV_X1 U7143 ( .A(n13320), .ZN(n13321) );
  BUF_X1 U7144 ( .A(n13324), .Z(n13322) );
  INV_X1 U7145 ( .A(n13326), .ZN(n13323) );
  INV_X1 U7146 ( .A(n13323), .ZN(n13324) );
  INV_X1 U7147 ( .A(n6628), .ZN(n13325) );
  INV_X1 U7148 ( .A(n13325), .ZN(n13326) );
  BUF_X1 U7149 ( .A(n13329), .Z(n13327) );
  INV_X1 U7150 ( .A(n13331), .ZN(n13328) );
  INV_X1 U7151 ( .A(n13328), .ZN(n13329) );
  INV_X1 U7152 ( .A(n6627), .ZN(n13330) );
  INV_X1 U7153 ( .A(n13330), .ZN(n13331) );
  BUF_X1 U7154 ( .A(n13334), .Z(n13332) );
  INV_X1 U7155 ( .A(n13336), .ZN(n13333) );
  INV_X1 U7156 ( .A(n13333), .ZN(n13334) );
  INV_X1 U7157 ( .A(n6626), .ZN(n13335) );
  INV_X1 U7158 ( .A(n13335), .ZN(n13336) );
  BUF_X1 U7159 ( .A(n13339), .Z(n13337) );
  INV_X1 U7160 ( .A(n13341), .ZN(n13338) );
  INV_X1 U7161 ( .A(n13338), .ZN(n13339) );
  INV_X1 U7162 ( .A(n6625), .ZN(n13340) );
  INV_X1 U7163 ( .A(n13340), .ZN(n13341) );
  BUF_X1 U7164 ( .A(n13344), .Z(n13342) );
  INV_X1 U7165 ( .A(n13346), .ZN(n13343) );
  INV_X1 U7166 ( .A(n13343), .ZN(n13344) );
  INV_X1 U7167 ( .A(n6624), .ZN(n13345) );
  INV_X1 U7168 ( .A(n13345), .ZN(n13346) );
  BUF_X1 U7169 ( .A(n13349), .Z(n13347) );
  INV_X1 U7170 ( .A(n13351), .ZN(n13348) );
  INV_X1 U7171 ( .A(n13348), .ZN(n13349) );
  INV_X1 U7172 ( .A(n6623), .ZN(n13350) );
  INV_X1 U7173 ( .A(n13350), .ZN(n13351) );
  BUF_X1 U7174 ( .A(n13354), .Z(n13352) );
  INV_X1 U7175 ( .A(n13356), .ZN(n13353) );
  INV_X1 U7176 ( .A(n13353), .ZN(n13354) );
  INV_X1 U7177 ( .A(n6622), .ZN(n13355) );
  INV_X1 U7178 ( .A(n13355), .ZN(n13356) );
  BUF_X1 U7179 ( .A(n13359), .Z(n13357) );
  INV_X1 U7180 ( .A(n13361), .ZN(n13358) );
  INV_X1 U7181 ( .A(n13358), .ZN(n13359) );
  INV_X1 U7182 ( .A(n6621), .ZN(n13360) );
  INV_X1 U7183 ( .A(n13360), .ZN(n13361) );
  BUF_X1 U7184 ( .A(n13364), .Z(n13362) );
  INV_X1 U7185 ( .A(n13366), .ZN(n13363) );
  INV_X1 U7186 ( .A(n13363), .ZN(n13364) );
  INV_X1 U7187 ( .A(n66200), .ZN(n13365) );
  INV_X1 U7188 ( .A(n13365), .ZN(n13366) );
  BUF_X1 U7189 ( .A(n13369), .Z(n13367) );
  INV_X1 U7190 ( .A(n13371), .ZN(n13368) );
  INV_X1 U7191 ( .A(n13368), .ZN(n13369) );
  INV_X1 U7192 ( .A(n66190), .ZN(n13370) );
  INV_X1 U7193 ( .A(n13370), .ZN(n13371) );
  BUF_X1 U7194 ( .A(n13374), .Z(n13372) );
  INV_X1 U7195 ( .A(n13376), .ZN(n13373) );
  INV_X1 U7196 ( .A(n13373), .ZN(n13374) );
  INV_X1 U7197 ( .A(n66180), .ZN(n13375) );
  INV_X1 U7198 ( .A(n13375), .ZN(n13376) );
  BUF_X1 U7199 ( .A(n13379), .Z(n13377) );
  INV_X1 U7200 ( .A(n13381), .ZN(n13378) );
  INV_X1 U7201 ( .A(n13378), .ZN(n13379) );
  INV_X1 U7202 ( .A(n66170), .ZN(n13380) );
  INV_X1 U7203 ( .A(n13380), .ZN(n13381) );
  BUF_X1 U7204 ( .A(n13384), .Z(n13382) );
  INV_X1 U7205 ( .A(n13386), .ZN(n13383) );
  INV_X1 U7206 ( .A(n13383), .ZN(n13384) );
  INV_X1 U7207 ( .A(n66160), .ZN(n13385) );
  INV_X1 U7208 ( .A(n13385), .ZN(n13386) );
  BUF_X1 U7209 ( .A(n13389), .Z(n13387) );
  INV_X1 U7210 ( .A(n13391), .ZN(n13388) );
  INV_X1 U7211 ( .A(n13388), .ZN(n13389) );
  INV_X1 U7212 ( .A(n66150), .ZN(n13390) );
  INV_X1 U7213 ( .A(n13390), .ZN(n13391) );
  BUF_X1 U7214 ( .A(n13394), .Z(n13392) );
  INV_X1 U7215 ( .A(n13396), .ZN(n13393) );
  INV_X1 U7216 ( .A(n13393), .ZN(n13394) );
  INV_X1 U7217 ( .A(n66140), .ZN(n13395) );
  INV_X1 U7218 ( .A(n13395), .ZN(n13396) );
  BUF_X1 U7219 ( .A(n13399), .Z(n13397) );
  INV_X1 U7220 ( .A(n13401), .ZN(n13398) );
  INV_X1 U7221 ( .A(n13398), .ZN(n13399) );
  INV_X1 U7222 ( .A(n66130), .ZN(n13400) );
  INV_X1 U7223 ( .A(n13400), .ZN(n13401) );
  BUF_X1 U7224 ( .A(n13404), .Z(n13402) );
  INV_X1 U7225 ( .A(n13406), .ZN(n13403) );
  INV_X1 U7226 ( .A(n13403), .ZN(n13404) );
  INV_X1 U7227 ( .A(n66120), .ZN(n13405) );
  INV_X1 U7228 ( .A(n13405), .ZN(n13406) );
  BUF_X1 U7229 ( .A(n13409), .Z(n13407) );
  INV_X1 U7230 ( .A(n13411), .ZN(n13408) );
  INV_X1 U7231 ( .A(n13408), .ZN(n13409) );
  INV_X1 U7232 ( .A(n66110), .ZN(n13410) );
  INV_X1 U7233 ( .A(n13410), .ZN(n13411) );
  BUF_X1 U7234 ( .A(n13414), .Z(n13412) );
  INV_X1 U7235 ( .A(n13416), .ZN(n13413) );
  INV_X1 U7236 ( .A(n13413), .ZN(n13414) );
  INV_X1 U7237 ( .A(n66100), .ZN(n13415) );
  INV_X1 U7238 ( .A(n13415), .ZN(n13416) );
  BUF_X1 U7239 ( .A(n13419), .Z(n13417) );
  INV_X1 U7240 ( .A(n13421), .ZN(n13418) );
  INV_X1 U7241 ( .A(n13418), .ZN(n13419) );
  INV_X1 U7242 ( .A(n66090), .ZN(n13420) );
  INV_X1 U7243 ( .A(n13420), .ZN(n13421) );
  BUF_X1 U7244 ( .A(n13424), .Z(n13422) );
  INV_X1 U7245 ( .A(n13426), .ZN(n13423) );
  INV_X1 U7246 ( .A(n13423), .ZN(n13424) );
  INV_X1 U7247 ( .A(n66080), .ZN(n13425) );
  INV_X1 U7248 ( .A(n13425), .ZN(n13426) );
  BUF_X1 U7249 ( .A(n13429), .Z(n13427) );
  INV_X1 U7250 ( .A(n13431), .ZN(n13428) );
  INV_X1 U7251 ( .A(n13428), .ZN(n13429) );
  INV_X1 U7252 ( .A(n66070), .ZN(n13430) );
  INV_X1 U7253 ( .A(n13430), .ZN(n13431) );
  BUF_X1 U7254 ( .A(n13434), .Z(n13432) );
  INV_X1 U7255 ( .A(n13436), .ZN(n13433) );
  INV_X1 U7256 ( .A(n13433), .ZN(n13434) );
  INV_X1 U7257 ( .A(n66060), .ZN(n13435) );
  INV_X1 U7258 ( .A(n13435), .ZN(n13436) );
  BUF_X1 U7259 ( .A(n13439), .Z(n13437) );
  INV_X1 U7260 ( .A(n13441), .ZN(n13438) );
  INV_X1 U7261 ( .A(n13438), .ZN(n13439) );
  INV_X1 U7262 ( .A(n66050), .ZN(n13440) );
  INV_X1 U7263 ( .A(n13440), .ZN(n13441) );
  BUF_X1 U7264 ( .A(n13444), .Z(n13442) );
  INV_X1 U7265 ( .A(n13446), .ZN(n13443) );
  INV_X1 U7266 ( .A(n13443), .ZN(n13444) );
  INV_X1 U7267 ( .A(n66040), .ZN(n13445) );
  INV_X1 U7268 ( .A(n13445), .ZN(n13446) );
  BUF_X1 U7269 ( .A(n13449), .Z(n13447) );
  INV_X1 U7270 ( .A(n13451), .ZN(n13448) );
  INV_X1 U7271 ( .A(n13448), .ZN(n13449) );
  INV_X1 U7272 ( .A(n66030), .ZN(n13450) );
  INV_X1 U7273 ( .A(n13450), .ZN(n13451) );
  BUF_X1 U7274 ( .A(n13454), .Z(n13452) );
  INV_X1 U7275 ( .A(n13456), .ZN(n13453) );
  INV_X1 U7276 ( .A(n13453), .ZN(n13454) );
  INV_X1 U7277 ( .A(n66020), .ZN(n13455) );
  INV_X1 U7278 ( .A(n13455), .ZN(n13456) );
  BUF_X1 U7279 ( .A(n13459), .Z(n13457) );
  INV_X1 U7280 ( .A(n13461), .ZN(n13458) );
  INV_X1 U7281 ( .A(n13458), .ZN(n13459) );
  INV_X1 U7282 ( .A(n66010), .ZN(n13460) );
  INV_X1 U7283 ( .A(n13460), .ZN(n13461) );
  BUF_X1 U7284 ( .A(n13464), .Z(n13462) );
  INV_X1 U7285 ( .A(n13466), .ZN(n13463) );
  INV_X1 U7286 ( .A(n13463), .ZN(n13464) );
  INV_X1 U7287 ( .A(n66000), .ZN(n13465) );
  INV_X1 U7288 ( .A(n13465), .ZN(n13466) );
  BUF_X1 U7289 ( .A(n13469), .Z(n13467) );
  INV_X1 U7290 ( .A(n13471), .ZN(n13468) );
  INV_X1 U7291 ( .A(n13468), .ZN(n13469) );
  INV_X1 U7292 ( .A(n6599), .ZN(n13470) );
  INV_X1 U7293 ( .A(n13470), .ZN(n13471) );
  BUF_X1 U7294 ( .A(n13474), .Z(n13472) );
  INV_X1 U7295 ( .A(n13476), .ZN(n13473) );
  INV_X1 U7296 ( .A(n13473), .ZN(n13474) );
  INV_X1 U7297 ( .A(n6598), .ZN(n13475) );
  INV_X1 U7298 ( .A(n13475), .ZN(n13476) );
  BUF_X1 U7299 ( .A(n13479), .Z(n13477) );
  INV_X1 U7300 ( .A(n13481), .ZN(n13478) );
  INV_X1 U7301 ( .A(n13478), .ZN(n13479) );
  INV_X1 U7302 ( .A(n6597), .ZN(n13480) );
  INV_X1 U7303 ( .A(n13480), .ZN(n13481) );
  BUF_X1 U7304 ( .A(n13484), .Z(n13482) );
  INV_X1 U7305 ( .A(n13486), .ZN(n13483) );
  INV_X1 U7306 ( .A(n13483), .ZN(n13484) );
  INV_X1 U7307 ( .A(n6596), .ZN(n13485) );
  INV_X1 U7308 ( .A(n13485), .ZN(n13486) );
  BUF_X1 U7309 ( .A(n13489), .Z(n13487) );
  INV_X1 U7310 ( .A(n13491), .ZN(n13488) );
  INV_X1 U7311 ( .A(n13488), .ZN(n13489) );
  INV_X1 U7312 ( .A(n6595), .ZN(n13490) );
  INV_X1 U7313 ( .A(n13490), .ZN(n13491) );
  BUF_X1 U7314 ( .A(n13494), .Z(n13492) );
  INV_X1 U7315 ( .A(n13496), .ZN(n13493) );
  INV_X1 U7316 ( .A(n13493), .ZN(n13494) );
  INV_X1 U7317 ( .A(n6594), .ZN(n13495) );
  INV_X1 U7318 ( .A(n13495), .ZN(n13496) );
  BUF_X1 U7319 ( .A(n13499), .Z(n13497) );
  INV_X1 U7320 ( .A(n13501), .ZN(n13498) );
  INV_X1 U7321 ( .A(n13498), .ZN(n13499) );
  INV_X1 U7322 ( .A(n6593), .ZN(n13500) );
  INV_X1 U7323 ( .A(n13500), .ZN(n13501) );
  BUF_X1 U7324 ( .A(n13504), .Z(n13502) );
  INV_X1 U7325 ( .A(n13506), .ZN(n13503) );
  INV_X1 U7326 ( .A(n13503), .ZN(n13504) );
  INV_X1 U7327 ( .A(n6592), .ZN(n13505) );
  INV_X1 U7328 ( .A(n13505), .ZN(n13506) );
  BUF_X1 U7329 ( .A(n13509), .Z(n13507) );
  INV_X1 U7330 ( .A(n13511), .ZN(n13508) );
  INV_X1 U7331 ( .A(n13508), .ZN(n13509) );
  INV_X1 U7332 ( .A(n6591), .ZN(n13510) );
  INV_X1 U7333 ( .A(n13510), .ZN(n13511) );
  BUF_X1 U7334 ( .A(n13514), .Z(n13512) );
  INV_X1 U7335 ( .A(n13516), .ZN(n13513) );
  INV_X1 U7336 ( .A(n13513), .ZN(n13514) );
  INV_X1 U7337 ( .A(n6590), .ZN(n13515) );
  INV_X1 U7338 ( .A(n13515), .ZN(n13516) );
  BUF_X1 U7339 ( .A(n13519), .Z(n13517) );
  INV_X1 U7340 ( .A(n13521), .ZN(n13518) );
  INV_X1 U7341 ( .A(n13518), .ZN(n13519) );
  INV_X1 U7342 ( .A(n6589), .ZN(n13520) );
  INV_X1 U7343 ( .A(n13520), .ZN(n13521) );
  BUF_X1 U7344 ( .A(n13524), .Z(n13522) );
  INV_X1 U7345 ( .A(n13526), .ZN(n13523) );
  INV_X1 U7346 ( .A(n13523), .ZN(n13524) );
  INV_X1 U7347 ( .A(n6588), .ZN(n13525) );
  INV_X1 U7348 ( .A(n13525), .ZN(n13526) );
  BUF_X1 U7349 ( .A(n13529), .Z(n13527) );
  INV_X1 U7350 ( .A(n13531), .ZN(n13528) );
  INV_X1 U7351 ( .A(n13528), .ZN(n13529) );
  INV_X1 U7352 ( .A(n6587), .ZN(n13530) );
  INV_X1 U7353 ( .A(n13530), .ZN(n13531) );
  BUF_X1 U7354 ( .A(n13534), .Z(n13532) );
  INV_X1 U7355 ( .A(n13536), .ZN(n13533) );
  INV_X1 U7356 ( .A(n13533), .ZN(n13534) );
  INV_X1 U7357 ( .A(n6586), .ZN(n13535) );
  INV_X1 U7358 ( .A(n13535), .ZN(n13536) );
  BUF_X1 U7359 ( .A(n13539), .Z(n13537) );
  INV_X1 U7360 ( .A(n13541), .ZN(n13538) );
  INV_X1 U7361 ( .A(n13538), .ZN(n13539) );
  INV_X1 U7362 ( .A(n6585), .ZN(n13540) );
  INV_X1 U7363 ( .A(n13540), .ZN(n13541) );
  BUF_X1 U7364 ( .A(n13544), .Z(n13542) );
  INV_X1 U7365 ( .A(n13546), .ZN(n13543) );
  INV_X1 U7366 ( .A(n13543), .ZN(n13544) );
  INV_X1 U7367 ( .A(n6584), .ZN(n13545) );
  INV_X1 U7368 ( .A(n13545), .ZN(n13546) );
  BUF_X1 U7369 ( .A(n13549), .Z(n13547) );
  INV_X1 U7370 ( .A(n13551), .ZN(n13548) );
  INV_X1 U7371 ( .A(n13548), .ZN(n13549) );
  INV_X1 U7372 ( .A(n6583), .ZN(n13550) );
  INV_X1 U7373 ( .A(n13550), .ZN(n13551) );
  BUF_X1 U7374 ( .A(n13554), .Z(n13552) );
  INV_X1 U7375 ( .A(n13556), .ZN(n13553) );
  INV_X1 U7376 ( .A(n13553), .ZN(n13554) );
  INV_X1 U7377 ( .A(n65820), .ZN(n13555) );
  INV_X1 U7378 ( .A(n13555), .ZN(n13556) );
  BUF_X1 U7379 ( .A(n13559), .Z(n13557) );
  INV_X1 U7380 ( .A(n13561), .ZN(n13558) );
  INV_X1 U7381 ( .A(n13558), .ZN(n13559) );
  INV_X1 U7382 ( .A(n65810), .ZN(n13560) );
  INV_X1 U7383 ( .A(n13560), .ZN(n13561) );
  BUF_X1 U7384 ( .A(n13564), .Z(n13562) );
  INV_X1 U7385 ( .A(n13566), .ZN(n13563) );
  INV_X1 U7386 ( .A(n13563), .ZN(n13564) );
  INV_X1 U7387 ( .A(n65800), .ZN(n13565) );
  INV_X1 U7388 ( .A(n13565), .ZN(n13566) );
  BUF_X1 U7389 ( .A(n13569), .Z(n13567) );
  INV_X1 U7390 ( .A(n13571), .ZN(n13568) );
  INV_X1 U7391 ( .A(n13568), .ZN(n13569) );
  INV_X1 U7392 ( .A(n65790), .ZN(n13570) );
  INV_X1 U7393 ( .A(n13570), .ZN(n13571) );
  BUF_X1 U7394 ( .A(n13574), .Z(n13572) );
  INV_X1 U7395 ( .A(n13576), .ZN(n13573) );
  INV_X1 U7396 ( .A(n13573), .ZN(n13574) );
  INV_X1 U7397 ( .A(n65780), .ZN(n13575) );
  INV_X1 U7398 ( .A(n13575), .ZN(n13576) );
  BUF_X1 U7399 ( .A(n13579), .Z(n13577) );
  INV_X1 U7400 ( .A(n13581), .ZN(n13578) );
  INV_X1 U7401 ( .A(n13578), .ZN(n13579) );
  INV_X1 U7402 ( .A(n65770), .ZN(n13580) );
  INV_X1 U7403 ( .A(n13580), .ZN(n13581) );
  BUF_X1 U7404 ( .A(n13584), .Z(n13582) );
  INV_X1 U7405 ( .A(n13586), .ZN(n13583) );
  INV_X1 U7406 ( .A(n13583), .ZN(n13584) );
  INV_X1 U7407 ( .A(n65760), .ZN(n13585) );
  INV_X1 U7408 ( .A(n13585), .ZN(n13586) );
  BUF_X1 U7409 ( .A(n13589), .Z(n13587) );
  INV_X1 U7410 ( .A(n13591), .ZN(n13588) );
  INV_X1 U7411 ( .A(n13588), .ZN(n13589) );
  INV_X1 U7412 ( .A(n65750), .ZN(n13590) );
  INV_X1 U7413 ( .A(n13590), .ZN(n13591) );
  BUF_X1 U7414 ( .A(n13594), .Z(n13592) );
  INV_X1 U7415 ( .A(n13596), .ZN(n13593) );
  INV_X1 U7416 ( .A(n13593), .ZN(n13594) );
  INV_X1 U7417 ( .A(n65740), .ZN(n13595) );
  INV_X1 U7418 ( .A(n13595), .ZN(n13596) );
  BUF_X1 U7419 ( .A(n13599), .Z(n13597) );
  INV_X1 U7420 ( .A(n13601), .ZN(n13598) );
  INV_X1 U7421 ( .A(n13598), .ZN(n13599) );
  INV_X1 U7422 ( .A(n65730), .ZN(n13600) );
  INV_X1 U7423 ( .A(n13600), .ZN(n13601) );
  BUF_X1 U7424 ( .A(n13604), .Z(n13602) );
  INV_X1 U7425 ( .A(n13606), .ZN(n13603) );
  INV_X1 U7426 ( .A(n13603), .ZN(n13604) );
  INV_X1 U7427 ( .A(n65720), .ZN(n13605) );
  INV_X1 U7428 ( .A(n13605), .ZN(n13606) );
  BUF_X1 U7429 ( .A(n13609), .Z(n13607) );
  INV_X1 U7430 ( .A(n13611), .ZN(n13608) );
  INV_X1 U7431 ( .A(n13608), .ZN(n13609) );
  INV_X1 U7432 ( .A(n65710), .ZN(n13610) );
  INV_X1 U7433 ( .A(n13610), .ZN(n13611) );
  BUF_X1 U7434 ( .A(n13614), .Z(n13612) );
  INV_X1 U7435 ( .A(n13616), .ZN(n13613) );
  INV_X1 U7436 ( .A(n13613), .ZN(n13614) );
  INV_X1 U7437 ( .A(n65700), .ZN(n13615) );
  INV_X1 U7438 ( .A(n13615), .ZN(n13616) );
  BUF_X1 U7439 ( .A(n13619), .Z(n13617) );
  INV_X1 U7440 ( .A(n13621), .ZN(n13618) );
  INV_X1 U7441 ( .A(n13618), .ZN(n13619) );
  INV_X1 U7442 ( .A(n65690), .ZN(n13620) );
  INV_X1 U7443 ( .A(n13620), .ZN(n13621) );
  BUF_X1 U7444 ( .A(n13624), .Z(n13622) );
  INV_X1 U7445 ( .A(n13626), .ZN(n13623) );
  INV_X1 U7446 ( .A(n13623), .ZN(n13624) );
  INV_X1 U7447 ( .A(n65680), .ZN(n13625) );
  INV_X1 U7448 ( .A(n13625), .ZN(n13626) );
  BUF_X1 U7449 ( .A(n13629), .Z(n13627) );
  INV_X1 U7450 ( .A(n13631), .ZN(n13628) );
  INV_X1 U7451 ( .A(n13628), .ZN(n13629) );
  INV_X1 U7452 ( .A(n65670), .ZN(n13630) );
  INV_X1 U7453 ( .A(n13630), .ZN(n13631) );
  BUF_X1 U7454 ( .A(n13634), .Z(n13632) );
  INV_X1 U7455 ( .A(n13636), .ZN(n13633) );
  INV_X1 U7456 ( .A(n13633), .ZN(n13634) );
  INV_X1 U7457 ( .A(n6566), .ZN(n13635) );
  INV_X1 U7458 ( .A(n13635), .ZN(n13636) );
  BUF_X1 U7459 ( .A(n13639), .Z(n13637) );
  INV_X1 U7460 ( .A(n13641), .ZN(n13638) );
  INV_X1 U7461 ( .A(n13638), .ZN(n13639) );
  INV_X1 U7462 ( .A(n6565), .ZN(n13640) );
  INV_X1 U7463 ( .A(n13640), .ZN(n13641) );
  BUF_X1 U7464 ( .A(n13644), .Z(n13642) );
  INV_X1 U7465 ( .A(n13646), .ZN(n13643) );
  INV_X1 U7466 ( .A(n13643), .ZN(n13644) );
  INV_X1 U7467 ( .A(n6564), .ZN(n13645) );
  INV_X1 U7468 ( .A(n13645), .ZN(n13646) );
  BUF_X1 U7469 ( .A(n13649), .Z(n13647) );
  INV_X1 U7470 ( .A(n13651), .ZN(n13648) );
  INV_X1 U7471 ( .A(n13648), .ZN(n13649) );
  INV_X1 U7472 ( .A(n65630), .ZN(n13650) );
  INV_X1 U7473 ( .A(n13650), .ZN(n13651) );
  BUF_X1 U7474 ( .A(n13654), .Z(n13652) );
  INV_X1 U7475 ( .A(n13656), .ZN(n13653) );
  INV_X1 U7476 ( .A(n13653), .ZN(n13654) );
  INV_X1 U7477 ( .A(n6562), .ZN(n13655) );
  INV_X1 U7478 ( .A(n13655), .ZN(n13656) );
  BUF_X1 U7479 ( .A(n13659), .Z(n13657) );
  INV_X1 U7480 ( .A(n13661), .ZN(n13658) );
  INV_X1 U7481 ( .A(n13658), .ZN(n13659) );
  INV_X1 U7482 ( .A(n6561), .ZN(n13660) );
  INV_X1 U7483 ( .A(n13660), .ZN(n13661) );
  BUF_X1 U7484 ( .A(n13664), .Z(n13662) );
  INV_X1 U7485 ( .A(n13666), .ZN(n13663) );
  INV_X1 U7486 ( .A(n13663), .ZN(n13664) );
  INV_X1 U7487 ( .A(n6560), .ZN(n13665) );
  INV_X1 U7488 ( .A(n13665), .ZN(n13666) );
  BUF_X1 U7489 ( .A(n13669), .Z(n13667) );
  INV_X1 U7490 ( .A(n13671), .ZN(n13668) );
  INV_X1 U7491 ( .A(n13668), .ZN(n13669) );
  INV_X1 U7492 ( .A(n6559), .ZN(n13670) );
  INV_X1 U7493 ( .A(n13670), .ZN(n13671) );
  BUF_X1 U7494 ( .A(n13674), .Z(n13672) );
  INV_X1 U7495 ( .A(n13676), .ZN(n13673) );
  INV_X1 U7496 ( .A(n13673), .ZN(n13674) );
  INV_X1 U7497 ( .A(n6558), .ZN(n13675) );
  INV_X1 U7498 ( .A(n13675), .ZN(n13676) );
  BUF_X1 U7499 ( .A(n13679), .Z(n13677) );
  INV_X1 U7500 ( .A(n13681), .ZN(n13678) );
  INV_X1 U7501 ( .A(n13678), .ZN(n13679) );
  INV_X1 U7502 ( .A(n6557), .ZN(n13680) );
  INV_X1 U7503 ( .A(n13680), .ZN(n13681) );
  BUF_X1 U7504 ( .A(n13684), .Z(n13682) );
  INV_X1 U7505 ( .A(n13686), .ZN(n13683) );
  INV_X1 U7506 ( .A(n13683), .ZN(n13684) );
  INV_X1 U7507 ( .A(n6556), .ZN(n13685) );
  INV_X1 U7508 ( .A(n13685), .ZN(n13686) );
  BUF_X1 U7509 ( .A(n13689), .Z(n13687) );
  INV_X1 U7510 ( .A(n13691), .ZN(n13688) );
  INV_X1 U7511 ( .A(n13688), .ZN(n13689) );
  INV_X1 U7512 ( .A(n6555), .ZN(n13690) );
  INV_X1 U7513 ( .A(n13690), .ZN(n13691) );
  BUF_X1 U7514 ( .A(n13694), .Z(n13692) );
  INV_X1 U7515 ( .A(n13696), .ZN(n13693) );
  INV_X1 U7516 ( .A(n13693), .ZN(n13694) );
  INV_X1 U7517 ( .A(n6554), .ZN(n13695) );
  INV_X1 U7518 ( .A(n13695), .ZN(n13696) );
  BUF_X1 U7519 ( .A(n13699), .Z(n13697) );
  INV_X1 U7520 ( .A(n13701), .ZN(n13698) );
  INV_X1 U7521 ( .A(n13698), .ZN(n13699) );
  INV_X1 U7522 ( .A(n6553), .ZN(n13700) );
  INV_X1 U7523 ( .A(n13700), .ZN(n13701) );
  BUF_X1 U7524 ( .A(n13704), .Z(n13702) );
  INV_X1 U7525 ( .A(n13706), .ZN(n13703) );
  INV_X1 U7526 ( .A(n13703), .ZN(n13704) );
  INV_X1 U7527 ( .A(n6552), .ZN(n13705) );
  INV_X1 U7528 ( .A(n13705), .ZN(n13706) );
  BUF_X1 U7529 ( .A(n13709), .Z(n13707) );
  INV_X1 U7530 ( .A(n13711), .ZN(n13708) );
  INV_X1 U7531 ( .A(n13708), .ZN(n13709) );
  INV_X1 U7532 ( .A(n6551), .ZN(n13710) );
  INV_X1 U7533 ( .A(n13710), .ZN(n13711) );
  BUF_X1 U7534 ( .A(n13714), .Z(n13712) );
  INV_X1 U7535 ( .A(n13716), .ZN(n13713) );
  INV_X1 U7536 ( .A(n13713), .ZN(n13714) );
  INV_X1 U7537 ( .A(n6550), .ZN(n13715) );
  INV_X1 U7538 ( .A(n13715), .ZN(n13716) );
  BUF_X1 U7539 ( .A(n13719), .Z(n13717) );
  INV_X1 U7540 ( .A(n13721), .ZN(n13718) );
  INV_X1 U7541 ( .A(n13718), .ZN(n13719) );
  INV_X1 U7542 ( .A(n6549), .ZN(n13720) );
  INV_X1 U7543 ( .A(n13720), .ZN(n13721) );
  BUF_X1 U7544 ( .A(n13724), .Z(n13722) );
  INV_X1 U7545 ( .A(n13726), .ZN(n13723) );
  INV_X1 U7546 ( .A(n13723), .ZN(n13724) );
  INV_X1 U7547 ( .A(n6548), .ZN(n13725) );
  INV_X1 U7548 ( .A(n13725), .ZN(n13726) );
  BUF_X1 U7549 ( .A(n13729), .Z(n13727) );
  INV_X1 U7550 ( .A(n13731), .ZN(n13728) );
  INV_X1 U7551 ( .A(n13728), .ZN(n13729) );
  INV_X1 U7552 ( .A(n6547), .ZN(n13730) );
  INV_X1 U7553 ( .A(n13730), .ZN(n13731) );
  BUF_X1 U7554 ( .A(n13734), .Z(n13732) );
  INV_X1 U7555 ( .A(n13736), .ZN(n13733) );
  INV_X1 U7556 ( .A(n13733), .ZN(n13734) );
  INV_X1 U7557 ( .A(n6546), .ZN(n13735) );
  INV_X1 U7558 ( .A(n13735), .ZN(n13736) );
  BUF_X1 U7559 ( .A(n13739), .Z(n13737) );
  INV_X1 U7560 ( .A(n13741), .ZN(n13738) );
  INV_X1 U7561 ( .A(n13738), .ZN(n13739) );
  INV_X1 U7562 ( .A(n6545), .ZN(n13740) );
  INV_X1 U7563 ( .A(n13740), .ZN(n13741) );
  BUF_X1 U7564 ( .A(n13744), .Z(n13742) );
  INV_X1 U7565 ( .A(n13746), .ZN(n13743) );
  INV_X1 U7566 ( .A(n13743), .ZN(n13744) );
  INV_X1 U7567 ( .A(n6544), .ZN(n13745) );
  INV_X1 U7568 ( .A(n13745), .ZN(n13746) );
  BUF_X1 U7569 ( .A(n13749), .Z(n13747) );
  INV_X1 U7570 ( .A(n13751), .ZN(n13748) );
  INV_X1 U7571 ( .A(n13748), .ZN(n13749) );
  INV_X1 U7572 ( .A(n6543), .ZN(n13750) );
  INV_X1 U7573 ( .A(n13750), .ZN(n13751) );
  BUF_X1 U7574 ( .A(n13754), .Z(n13752) );
  INV_X1 U7575 ( .A(n13756), .ZN(n13753) );
  INV_X1 U7576 ( .A(n13753), .ZN(n13754) );
  INV_X1 U7577 ( .A(n6542), .ZN(n13755) );
  INV_X1 U7578 ( .A(n13755), .ZN(n13756) );
  BUF_X1 U7579 ( .A(n13759), .Z(n13757) );
  INV_X1 U7580 ( .A(n13761), .ZN(n13758) );
  INV_X1 U7581 ( .A(n13758), .ZN(n13759) );
  INV_X1 U7582 ( .A(n6541), .ZN(n13760) );
  INV_X1 U7583 ( .A(n13760), .ZN(n13761) );
  BUF_X1 U7584 ( .A(n13764), .Z(n13762) );
  INV_X1 U7585 ( .A(n13766), .ZN(n13763) );
  INV_X1 U7586 ( .A(n13763), .ZN(n13764) );
  INV_X1 U7587 ( .A(n6540), .ZN(n13765) );
  INV_X1 U7588 ( .A(n13765), .ZN(n13766) );
  BUF_X1 U7589 ( .A(n13769), .Z(n13767) );
  INV_X1 U7590 ( .A(n13771), .ZN(n13768) );
  INV_X1 U7591 ( .A(n13768), .ZN(n13769) );
  INV_X1 U7592 ( .A(n6539), .ZN(n13770) );
  INV_X1 U7593 ( .A(n13770), .ZN(n13771) );
  BUF_X1 U7594 ( .A(n13774), .Z(n13772) );
  INV_X1 U7595 ( .A(n13776), .ZN(n13773) );
  INV_X1 U7596 ( .A(n13773), .ZN(n13774) );
  INV_X1 U7597 ( .A(n65380), .ZN(n13775) );
  INV_X1 U7598 ( .A(n13775), .ZN(n13776) );
  BUF_X1 U7599 ( .A(n13779), .Z(n13777) );
  INV_X1 U7600 ( .A(n13781), .ZN(n13778) );
  INV_X1 U7601 ( .A(n13778), .ZN(n13779) );
  INV_X1 U7602 ( .A(n65370), .ZN(n13780) );
  INV_X1 U7603 ( .A(n13780), .ZN(n13781) );
  BUF_X1 U7604 ( .A(n13784), .Z(n13782) );
  INV_X1 U7605 ( .A(n13786), .ZN(n13783) );
  INV_X1 U7606 ( .A(n13783), .ZN(n13784) );
  INV_X1 U7607 ( .A(n65360), .ZN(n13785) );
  INV_X1 U7608 ( .A(n13785), .ZN(n13786) );
  BUF_X1 U7609 ( .A(n13789), .Z(n13787) );
  INV_X1 U7610 ( .A(n13791), .ZN(n13788) );
  INV_X1 U7611 ( .A(n13788), .ZN(n13789) );
  INV_X1 U7612 ( .A(n65350), .ZN(n13790) );
  INV_X1 U7613 ( .A(n13790), .ZN(n13791) );
  BUF_X1 U7614 ( .A(n13794), .Z(n13792) );
  INV_X1 U7615 ( .A(n13796), .ZN(n13793) );
  INV_X1 U7616 ( .A(n13793), .ZN(n13794) );
  INV_X1 U7617 ( .A(n65340), .ZN(n13795) );
  INV_X1 U7618 ( .A(n13795), .ZN(n13796) );
  BUF_X1 U7619 ( .A(n13799), .Z(n13797) );
  INV_X1 U7620 ( .A(n13801), .ZN(n13798) );
  INV_X1 U7621 ( .A(n13798), .ZN(n13799) );
  INV_X1 U7622 ( .A(n65330), .ZN(n13800) );
  INV_X1 U7623 ( .A(n13800), .ZN(n13801) );
  BUF_X1 U7624 ( .A(n13804), .Z(n13802) );
  INV_X1 U7625 ( .A(n13806), .ZN(n13803) );
  INV_X1 U7626 ( .A(n13803), .ZN(n13804) );
  INV_X1 U7627 ( .A(n65320), .ZN(n13805) );
  INV_X1 U7628 ( .A(n13805), .ZN(n13806) );
  BUF_X1 U7629 ( .A(n13809), .Z(n13807) );
  INV_X1 U7630 ( .A(n13811), .ZN(n13808) );
  INV_X1 U7631 ( .A(n13808), .ZN(n13809) );
  INV_X1 U7632 ( .A(n65310), .ZN(n13810) );
  INV_X1 U7633 ( .A(n13810), .ZN(n13811) );
  BUF_X1 U7634 ( .A(n13814), .Z(n13812) );
  INV_X1 U7635 ( .A(n13816), .ZN(n13813) );
  INV_X1 U7636 ( .A(n13813), .ZN(n13814) );
  INV_X1 U7637 ( .A(n65300), .ZN(n13815) );
  INV_X1 U7638 ( .A(n13815), .ZN(n13816) );
  BUF_X1 U7639 ( .A(n13819), .Z(n13817) );
  INV_X1 U7640 ( .A(n13821), .ZN(n13818) );
  INV_X1 U7641 ( .A(n13818), .ZN(n13819) );
  INV_X1 U7642 ( .A(n65290), .ZN(n13820) );
  INV_X1 U7643 ( .A(n13820), .ZN(n13821) );
  BUF_X1 U7644 ( .A(n13824), .Z(n13822) );
  INV_X1 U7645 ( .A(n13826), .ZN(n13823) );
  INV_X1 U7646 ( .A(n13823), .ZN(n13824) );
  INV_X1 U7647 ( .A(n65280), .ZN(n13825) );
  INV_X1 U7648 ( .A(n13825), .ZN(n13826) );
  BUF_X1 U7649 ( .A(n13829), .Z(n13827) );
  INV_X1 U7650 ( .A(n13831), .ZN(n13828) );
  INV_X1 U7651 ( .A(n13828), .ZN(n13829) );
  INV_X1 U7652 ( .A(n65270), .ZN(n13830) );
  INV_X1 U7653 ( .A(n13830), .ZN(n13831) );
  BUF_X1 U7654 ( .A(n13834), .Z(n13832) );
  INV_X1 U7655 ( .A(n13836), .ZN(n13833) );
  INV_X1 U7656 ( .A(n13833), .ZN(n13834) );
  INV_X1 U7657 ( .A(n65260), .ZN(n13835) );
  INV_X1 U7658 ( .A(n13835), .ZN(n13836) );
  BUF_X1 U7659 ( .A(n13839), .Z(n13837) );
  INV_X1 U7660 ( .A(n13841), .ZN(n13838) );
  INV_X1 U7661 ( .A(n13838), .ZN(n13839) );
  INV_X1 U7662 ( .A(n65250), .ZN(n13840) );
  INV_X1 U7663 ( .A(n13840), .ZN(n13841) );
  BUF_X1 U7664 ( .A(n13844), .Z(n13842) );
  INV_X1 U7665 ( .A(n13846), .ZN(n13843) );
  INV_X1 U7666 ( .A(n13843), .ZN(n13844) );
  INV_X1 U7667 ( .A(n65240), .ZN(n13845) );
  INV_X1 U7668 ( .A(n13845), .ZN(n13846) );
  BUF_X1 U7669 ( .A(n13849), .Z(n13847) );
  INV_X1 U7670 ( .A(n13851), .ZN(n13848) );
  INV_X1 U7671 ( .A(n13848), .ZN(n13849) );
  INV_X1 U7672 ( .A(n65230), .ZN(n13850) );
  INV_X1 U7673 ( .A(n13850), .ZN(n13851) );
  BUF_X1 U7674 ( .A(n13854), .Z(n13852) );
  INV_X1 U7675 ( .A(n13856), .ZN(n13853) );
  INV_X1 U7676 ( .A(n13853), .ZN(n13854) );
  INV_X1 U7677 ( .A(n65220), .ZN(n13855) );
  INV_X1 U7678 ( .A(n13855), .ZN(n13856) );
  BUF_X1 U7679 ( .A(n13859), .Z(n13857) );
  INV_X1 U7680 ( .A(n13861), .ZN(n13858) );
  INV_X1 U7681 ( .A(n13858), .ZN(n13859) );
  INV_X1 U7682 ( .A(n65210), .ZN(n13860) );
  INV_X1 U7683 ( .A(n13860), .ZN(n13861) );
  BUF_X1 U7684 ( .A(n13864), .Z(n13862) );
  INV_X1 U7685 ( .A(n13866), .ZN(n13863) );
  INV_X1 U7686 ( .A(n13863), .ZN(n13864) );
  INV_X1 U7687 ( .A(n65200), .ZN(n13865) );
  INV_X1 U7688 ( .A(n13865), .ZN(n13866) );
  BUF_X1 U7689 ( .A(n13869), .Z(n13867) );
  INV_X1 U7690 ( .A(n13871), .ZN(n13868) );
  INV_X1 U7691 ( .A(n13868), .ZN(n13869) );
  INV_X1 U7692 ( .A(n65190), .ZN(n13870) );
  INV_X1 U7693 ( .A(n13870), .ZN(n13871) );
  BUF_X1 U7694 ( .A(n13874), .Z(n13872) );
  INV_X1 U7695 ( .A(n13876), .ZN(n13873) );
  INV_X1 U7696 ( .A(n13873), .ZN(n13874) );
  INV_X1 U7697 ( .A(n65180), .ZN(n13875) );
  INV_X1 U7698 ( .A(n13875), .ZN(n13876) );
  BUF_X1 U7699 ( .A(n13879), .Z(n13877) );
  INV_X1 U7700 ( .A(n13881), .ZN(n13878) );
  INV_X1 U7701 ( .A(n13878), .ZN(n13879) );
  INV_X1 U7702 ( .A(n6517), .ZN(n13880) );
  INV_X1 U7703 ( .A(n13880), .ZN(n13881) );
  BUF_X1 U7704 ( .A(n13884), .Z(n13882) );
  INV_X1 U7705 ( .A(n13886), .ZN(n13883) );
  INV_X1 U7706 ( .A(n13883), .ZN(n13884) );
  INV_X1 U7707 ( .A(n6516), .ZN(n13885) );
  INV_X1 U7708 ( .A(n13885), .ZN(n13886) );
  BUF_X1 U7709 ( .A(n13889), .Z(n13887) );
  INV_X1 U7710 ( .A(n13891), .ZN(n13888) );
  INV_X1 U7711 ( .A(n13888), .ZN(n13889) );
  INV_X1 U7712 ( .A(n6515), .ZN(n13890) );
  INV_X1 U7713 ( .A(n13890), .ZN(n13891) );
  BUF_X1 U7714 ( .A(n13894), .Z(n13892) );
  INV_X1 U7715 ( .A(n13896), .ZN(n13893) );
  INV_X1 U7716 ( .A(n13893), .ZN(n13894) );
  INV_X1 U7717 ( .A(n6514), .ZN(n13895) );
  INV_X1 U7718 ( .A(n13895), .ZN(n13896) );
  BUF_X1 U7719 ( .A(n13899), .Z(n13897) );
  INV_X1 U7720 ( .A(n13901), .ZN(n13898) );
  INV_X1 U7721 ( .A(n13898), .ZN(n13899) );
  INV_X1 U7722 ( .A(n6513), .ZN(n13900) );
  INV_X1 U7723 ( .A(n13900), .ZN(n13901) );
  BUF_X1 U7724 ( .A(n13904), .Z(n13902) );
  INV_X1 U7725 ( .A(n13906), .ZN(n13903) );
  INV_X1 U7726 ( .A(n13903), .ZN(n13904) );
  INV_X1 U7727 ( .A(n6512), .ZN(n13905) );
  INV_X1 U7728 ( .A(n13905), .ZN(n13906) );
  BUF_X1 U7729 ( .A(n13909), .Z(n13907) );
  INV_X1 U7730 ( .A(n13911), .ZN(n13908) );
  INV_X1 U7731 ( .A(n13908), .ZN(n13909) );
  INV_X1 U7732 ( .A(n6511), .ZN(n13910) );
  INV_X1 U7733 ( .A(n13910), .ZN(n13911) );
  BUF_X1 U7734 ( .A(n13914), .Z(n13912) );
  INV_X1 U7735 ( .A(n13916), .ZN(n13913) );
  INV_X1 U7736 ( .A(n13913), .ZN(n13914) );
  INV_X1 U7737 ( .A(n6510), .ZN(n13915) );
  INV_X1 U7738 ( .A(n13915), .ZN(n13916) );
  BUF_X1 U7739 ( .A(n13919), .Z(n13917) );
  INV_X1 U7740 ( .A(n13921), .ZN(n13918) );
  INV_X1 U7741 ( .A(n13918), .ZN(n13919) );
  INV_X1 U7742 ( .A(n6509), .ZN(n13920) );
  INV_X1 U7743 ( .A(n13920), .ZN(n13921) );
  BUF_X1 U7744 ( .A(n13924), .Z(n13922) );
  INV_X1 U7745 ( .A(n13926), .ZN(n13923) );
  INV_X1 U7746 ( .A(n13923), .ZN(n13924) );
  INV_X1 U7747 ( .A(n6508), .ZN(n13925) );
  INV_X1 U7748 ( .A(n13925), .ZN(n13926) );
  BUF_X1 U7749 ( .A(n13929), .Z(n13927) );
  INV_X1 U7750 ( .A(n13931), .ZN(n13928) );
  INV_X1 U7751 ( .A(n13928), .ZN(n13929) );
  INV_X1 U7752 ( .A(n6507), .ZN(n13930) );
  INV_X1 U7753 ( .A(n13930), .ZN(n13931) );
  BUF_X1 U7754 ( .A(n13934), .Z(n13932) );
  INV_X1 U7755 ( .A(n13936), .ZN(n13933) );
  INV_X1 U7756 ( .A(n13933), .ZN(n13934) );
  INV_X1 U7757 ( .A(n6506), .ZN(n13935) );
  INV_X1 U7758 ( .A(n13935), .ZN(n13936) );
  BUF_X1 U7759 ( .A(n13939), .Z(n13937) );
  INV_X1 U7760 ( .A(n13941), .ZN(n13938) );
  INV_X1 U7761 ( .A(n13938), .ZN(n13939) );
  INV_X1 U7762 ( .A(n6505), .ZN(n13940) );
  INV_X1 U7763 ( .A(n13940), .ZN(n13941) );
  BUF_X1 U7764 ( .A(n13944), .Z(n13942) );
  INV_X1 U7765 ( .A(n13946), .ZN(n13943) );
  INV_X1 U7766 ( .A(n13943), .ZN(n13944) );
  INV_X1 U7767 ( .A(n6504), .ZN(n13945) );
  INV_X1 U7768 ( .A(n13945), .ZN(n13946) );
  BUF_X1 U7769 ( .A(n13949), .Z(n13947) );
  INV_X1 U7770 ( .A(n13951), .ZN(n13948) );
  INV_X1 U7771 ( .A(n13948), .ZN(n13949) );
  INV_X1 U7772 ( .A(n6503), .ZN(n13950) );
  INV_X1 U7773 ( .A(n13950), .ZN(n13951) );
  BUF_X1 U7774 ( .A(n13954), .Z(n13952) );
  INV_X1 U7775 ( .A(n13956), .ZN(n13953) );
  INV_X1 U7776 ( .A(n13953), .ZN(n13954) );
  INV_X1 U7777 ( .A(n6502), .ZN(n13955) );
  INV_X1 U7778 ( .A(n13955), .ZN(n13956) );
  BUF_X1 U7779 ( .A(n13959), .Z(n13957) );
  INV_X1 U7780 ( .A(n13961), .ZN(n13958) );
  INV_X1 U7781 ( .A(n13958), .ZN(n13959) );
  INV_X1 U7782 ( .A(n6501), .ZN(n13960) );
  INV_X1 U7783 ( .A(n13960), .ZN(n13961) );
  BUF_X1 U7784 ( .A(n13964), .Z(n13962) );
  INV_X1 U7785 ( .A(n13966), .ZN(n13963) );
  INV_X1 U7786 ( .A(n13963), .ZN(n13964) );
  INV_X1 U7787 ( .A(n65000), .ZN(n13965) );
  INV_X1 U7788 ( .A(n13965), .ZN(n13966) );
  BUF_X1 U7789 ( .A(n13969), .Z(n13967) );
  INV_X1 U7790 ( .A(n13971), .ZN(n13968) );
  INV_X1 U7791 ( .A(n13968), .ZN(n13969) );
  INV_X1 U7792 ( .A(n64990), .ZN(n13970) );
  INV_X1 U7793 ( .A(n13970), .ZN(n13971) );
  BUF_X1 U7794 ( .A(n13974), .Z(n13972) );
  INV_X1 U7795 ( .A(n13976), .ZN(n13973) );
  INV_X1 U7796 ( .A(n13973), .ZN(n13974) );
  INV_X1 U7797 ( .A(n64980), .ZN(n13975) );
  INV_X1 U7798 ( .A(n13975), .ZN(n13976) );
  BUF_X1 U7799 ( .A(n13979), .Z(n13977) );
  INV_X1 U7800 ( .A(n13981), .ZN(n13978) );
  INV_X1 U7801 ( .A(n13978), .ZN(n13979) );
  INV_X1 U7802 ( .A(n64970), .ZN(n13980) );
  INV_X1 U7803 ( .A(n13980), .ZN(n13981) );
  BUF_X1 U7804 ( .A(n13984), .Z(n13982) );
  INV_X1 U7805 ( .A(n13986), .ZN(n13983) );
  INV_X1 U7806 ( .A(n13983), .ZN(n13984) );
  INV_X1 U7807 ( .A(n64960), .ZN(n13985) );
  INV_X1 U7808 ( .A(n13985), .ZN(n13986) );
  BUF_X1 U7809 ( .A(n13989), .Z(n13987) );
  INV_X1 U7810 ( .A(n13991), .ZN(n13988) );
  INV_X1 U7811 ( .A(n13988), .ZN(n13989) );
  INV_X1 U7812 ( .A(n64950), .ZN(n13990) );
  INV_X1 U7813 ( .A(n13990), .ZN(n13991) );
  BUF_X1 U7814 ( .A(n13994), .Z(n13992) );
  INV_X1 U7815 ( .A(n13996), .ZN(n13993) );
  INV_X1 U7816 ( .A(n13993), .ZN(n13994) );
  INV_X1 U7817 ( .A(n64940), .ZN(n13995) );
  INV_X1 U7818 ( .A(n13995), .ZN(n13996) );
  BUF_X1 U7819 ( .A(n13999), .Z(n13997) );
  INV_X1 U7820 ( .A(n14001), .ZN(n13998) );
  INV_X1 U7821 ( .A(n13998), .ZN(n13999) );
  INV_X1 U7822 ( .A(n64930), .ZN(n14000) );
  INV_X1 U7823 ( .A(n14000), .ZN(n14001) );
  BUF_X1 U7824 ( .A(n14004), .Z(n14002) );
  INV_X1 U7825 ( .A(n14006), .ZN(n14003) );
  INV_X1 U7826 ( .A(n14003), .ZN(n14004) );
  INV_X1 U7827 ( .A(n64920), .ZN(n14005) );
  INV_X1 U7828 ( .A(n14005), .ZN(n14006) );
  BUF_X1 U7829 ( .A(n14009), .Z(n14007) );
  INV_X1 U7830 ( .A(n14011), .ZN(n14008) );
  INV_X1 U7831 ( .A(n14008), .ZN(n14009) );
  INV_X1 U7832 ( .A(n64910), .ZN(n14010) );
  INV_X1 U7833 ( .A(n14010), .ZN(n14011) );
  BUF_X1 U7834 ( .A(n14014), .Z(n14012) );
  INV_X1 U7835 ( .A(n14016), .ZN(n14013) );
  INV_X1 U7836 ( .A(n14013), .ZN(n14014) );
  INV_X1 U7837 ( .A(n64900), .ZN(n14015) );
  INV_X1 U7838 ( .A(n14015), .ZN(n14016) );
  BUF_X1 U7839 ( .A(n14019), .Z(n14017) );
  INV_X1 U7840 ( .A(n14021), .ZN(n14018) );
  INV_X1 U7841 ( .A(n14018), .ZN(n14019) );
  INV_X1 U7842 ( .A(n64890), .ZN(n14020) );
  INV_X1 U7843 ( .A(n14020), .ZN(n14021) );
  BUF_X1 U7844 ( .A(n14024), .Z(n14022) );
  INV_X1 U7845 ( .A(n14026), .ZN(n14023) );
  INV_X1 U7846 ( .A(n14023), .ZN(n14024) );
  INV_X1 U7847 ( .A(n64880), .ZN(n14025) );
  INV_X1 U7848 ( .A(n14025), .ZN(n14026) );
  BUF_X1 U7849 ( .A(n14029), .Z(n14027) );
  INV_X1 U7850 ( .A(n14031), .ZN(n14028) );
  INV_X1 U7851 ( .A(n14028), .ZN(n14029) );
  INV_X1 U7852 ( .A(n64870), .ZN(n14030) );
  INV_X1 U7853 ( .A(n14030), .ZN(n14031) );
  BUF_X1 U7854 ( .A(n14034), .Z(n14032) );
  INV_X1 U7855 ( .A(n14036), .ZN(n14033) );
  INV_X1 U7856 ( .A(n14033), .ZN(n14034) );
  INV_X1 U7857 ( .A(n64860), .ZN(n14035) );
  INV_X1 U7858 ( .A(n14035), .ZN(n14036) );
  BUF_X1 U7859 ( .A(n14039), .Z(n14037) );
  INV_X1 U7860 ( .A(n14041), .ZN(n14038) );
  INV_X1 U7861 ( .A(n14038), .ZN(n14039) );
  INV_X1 U7862 ( .A(n64850), .ZN(n14040) );
  INV_X1 U7863 ( .A(n14040), .ZN(n14041) );
  BUF_X1 U7864 ( .A(n14044), .Z(n14042) );
  INV_X1 U7865 ( .A(n14046), .ZN(n14043) );
  INV_X1 U7866 ( .A(n14043), .ZN(n14044) );
  INV_X1 U7867 ( .A(n6484), .ZN(n14045) );
  INV_X1 U7868 ( .A(n14045), .ZN(n14046) );
  BUF_X1 U7869 ( .A(n14049), .Z(n14047) );
  INV_X1 U7870 ( .A(n14051), .ZN(n14048) );
  INV_X1 U7871 ( .A(n14048), .ZN(n14049) );
  INV_X1 U7872 ( .A(n6483), .ZN(n14050) );
  INV_X1 U7873 ( .A(n14050), .ZN(n14051) );
  BUF_X1 U7874 ( .A(n14054), .Z(n14052) );
  INV_X1 U7875 ( .A(n14056), .ZN(n14053) );
  INV_X1 U7876 ( .A(n14053), .ZN(n14054) );
  INV_X1 U7877 ( .A(n6482), .ZN(n14055) );
  INV_X1 U7878 ( .A(n14055), .ZN(n14056) );
  BUF_X1 U7879 ( .A(n14059), .Z(n14057) );
  INV_X1 U7880 ( .A(n14061), .ZN(n14058) );
  INV_X1 U7881 ( .A(n14058), .ZN(n14059) );
  INV_X1 U7882 ( .A(n6481), .ZN(n14060) );
  INV_X1 U7883 ( .A(n14060), .ZN(n14061) );
  BUF_X1 U7884 ( .A(n14064), .Z(n14062) );
  INV_X1 U7885 ( .A(n14066), .ZN(n14063) );
  INV_X1 U7886 ( .A(n14063), .ZN(n14064) );
  INV_X1 U7887 ( .A(n6480), .ZN(n14065) );
  INV_X1 U7888 ( .A(n14065), .ZN(n14066) );
  BUF_X1 U7889 ( .A(n14069), .Z(n14067) );
  INV_X1 U7890 ( .A(n14071), .ZN(n14068) );
  INV_X1 U7891 ( .A(n14068), .ZN(n14069) );
  INV_X1 U7892 ( .A(n6479), .ZN(n14070) );
  INV_X1 U7893 ( .A(n14070), .ZN(n14071) );
  BUF_X1 U7894 ( .A(n14074), .Z(n14072) );
  INV_X1 U7895 ( .A(n14076), .ZN(n14073) );
  INV_X1 U7896 ( .A(n14073), .ZN(n14074) );
  INV_X1 U7897 ( .A(n6478), .ZN(n14075) );
  INV_X1 U7898 ( .A(n14075), .ZN(n14076) );
  BUF_X1 U7899 ( .A(n14079), .Z(n14077) );
  INV_X1 U7900 ( .A(n14081), .ZN(n14078) );
  INV_X1 U7901 ( .A(n14078), .ZN(n14079) );
  INV_X1 U7902 ( .A(n6477), .ZN(n14080) );
  INV_X1 U7903 ( .A(n14080), .ZN(n14081) );
  BUF_X1 U7904 ( .A(n14084), .Z(n14082) );
  INV_X1 U7905 ( .A(n14086), .ZN(n14083) );
  INV_X1 U7906 ( .A(n14083), .ZN(n14084) );
  INV_X1 U7907 ( .A(n6476), .ZN(n14085) );
  INV_X1 U7908 ( .A(n14085), .ZN(n14086) );
  BUF_X1 U7909 ( .A(n14089), .Z(n14087) );
  INV_X1 U7910 ( .A(n14091), .ZN(n14088) );
  INV_X1 U7911 ( .A(n14088), .ZN(n14089) );
  INV_X1 U7912 ( .A(n6475), .ZN(n14090) );
  INV_X1 U7913 ( .A(n14090), .ZN(n14091) );
  BUF_X1 U7914 ( .A(n14094), .Z(n14092) );
  INV_X1 U7915 ( .A(n14096), .ZN(n14093) );
  INV_X1 U7916 ( .A(n14093), .ZN(n14094) );
  INV_X1 U7917 ( .A(n6474), .ZN(n14095) );
  INV_X1 U7918 ( .A(n14095), .ZN(n14096) );
  BUF_X1 U7919 ( .A(n14099), .Z(n14097) );
  INV_X1 U7920 ( .A(n14101), .ZN(n14098) );
  INV_X1 U7921 ( .A(n14098), .ZN(n14099) );
  INV_X1 U7922 ( .A(n6473), .ZN(n14100) );
  INV_X1 U7923 ( .A(n14100), .ZN(n14101) );
  BUF_X1 U7924 ( .A(n14104), .Z(n14102) );
  INV_X1 U7925 ( .A(n14106), .ZN(n14103) );
  INV_X1 U7926 ( .A(n14103), .ZN(n14104) );
  INV_X1 U7927 ( .A(n6472), .ZN(n14105) );
  INV_X1 U7928 ( .A(n14105), .ZN(n14106) );
  BUF_X1 U7929 ( .A(n14109), .Z(n14107) );
  INV_X1 U7930 ( .A(n14111), .ZN(n14108) );
  INV_X1 U7931 ( .A(n14108), .ZN(n14109) );
  INV_X1 U7932 ( .A(n6471), .ZN(n14110) );
  INV_X1 U7933 ( .A(n14110), .ZN(n14111) );
  BUF_X1 U7934 ( .A(n14114), .Z(n14112) );
  INV_X1 U7935 ( .A(n14116), .ZN(n14113) );
  INV_X1 U7936 ( .A(n14113), .ZN(n14114) );
  INV_X1 U7937 ( .A(n6470), .ZN(n14115) );
  INV_X1 U7938 ( .A(n14115), .ZN(n14116) );
  BUF_X1 U7939 ( .A(n14119), .Z(n14117) );
  INV_X1 U7940 ( .A(n14121), .ZN(n14118) );
  INV_X1 U7941 ( .A(n14118), .ZN(n14119) );
  INV_X1 U7942 ( .A(n6469), .ZN(n14120) );
  INV_X1 U7943 ( .A(n14120), .ZN(n14121) );
  BUF_X1 U7944 ( .A(n14124), .Z(n14122) );
  INV_X1 U7945 ( .A(n14126), .ZN(n14123) );
  INV_X1 U7946 ( .A(n14123), .ZN(n14124) );
  INV_X1 U7947 ( .A(n6468), .ZN(n14125) );
  INV_X1 U7948 ( .A(n14125), .ZN(n14126) );
  BUF_X1 U7949 ( .A(n14129), .Z(n14127) );
  INV_X1 U7950 ( .A(n14131), .ZN(n14128) );
  INV_X1 U7951 ( .A(n14128), .ZN(n14129) );
  INV_X1 U7952 ( .A(n6467), .ZN(n14130) );
  INV_X1 U7953 ( .A(n14130), .ZN(n14131) );
  BUF_X1 U7954 ( .A(n14134), .Z(n14132) );
  INV_X1 U7955 ( .A(n14136), .ZN(n14133) );
  INV_X1 U7956 ( .A(n14133), .ZN(n14134) );
  INV_X1 U7957 ( .A(n6466), .ZN(n14135) );
  INV_X1 U7958 ( .A(n14135), .ZN(n14136) );
  BUF_X1 U7959 ( .A(n14139), .Z(n14137) );
  INV_X1 U7960 ( .A(n14141), .ZN(n14138) );
  INV_X1 U7961 ( .A(n14138), .ZN(n14139) );
  INV_X1 U7962 ( .A(n6465), .ZN(n14140) );
  INV_X1 U7963 ( .A(n14140), .ZN(n14141) );
  BUF_X1 U7964 ( .A(n14144), .Z(n14142) );
  INV_X1 U7965 ( .A(n14146), .ZN(n14143) );
  INV_X1 U7966 ( .A(n14143), .ZN(n14144) );
  INV_X1 U7967 ( .A(n6464), .ZN(n14145) );
  INV_X1 U7968 ( .A(n14145), .ZN(n14146) );
  BUF_X1 U7969 ( .A(n14149), .Z(n14147) );
  INV_X1 U7970 ( .A(n14151), .ZN(n14148) );
  INV_X1 U7971 ( .A(n14148), .ZN(n14149) );
  INV_X1 U7972 ( .A(n6463), .ZN(n14150) );
  INV_X1 U7973 ( .A(n14150), .ZN(n14151) );
  BUF_X1 U7974 ( .A(n14154), .Z(n14152) );
  INV_X1 U7975 ( .A(n14156), .ZN(n14153) );
  INV_X1 U7976 ( .A(n14153), .ZN(n14154) );
  INV_X1 U7977 ( .A(n6462), .ZN(n14155) );
  INV_X1 U7978 ( .A(n14155), .ZN(n14156) );
  BUF_X1 U7979 ( .A(n14159), .Z(n14157) );
  INV_X1 U7980 ( .A(n14161), .ZN(n14158) );
  INV_X1 U7981 ( .A(n14158), .ZN(n14159) );
  INV_X1 U7982 ( .A(n6461), .ZN(n14160) );
  INV_X1 U7983 ( .A(n14160), .ZN(n14161) );
  BUF_X1 U7984 ( .A(n14164), .Z(n14162) );
  INV_X1 U7985 ( .A(n14166), .ZN(n14163) );
  INV_X1 U7986 ( .A(n14163), .ZN(n14164) );
  INV_X1 U7987 ( .A(n6460), .ZN(n14165) );
  INV_X1 U7988 ( .A(n14165), .ZN(n14166) );
  BUF_X1 U7989 ( .A(n14169), .Z(n14167) );
  INV_X1 U7990 ( .A(n14171), .ZN(n14168) );
  INV_X1 U7991 ( .A(n14168), .ZN(n14169) );
  INV_X1 U7992 ( .A(n6459), .ZN(n14170) );
  INV_X1 U7993 ( .A(n14170), .ZN(n14171) );
  BUF_X1 U7994 ( .A(n14174), .Z(n14172) );
  INV_X1 U7995 ( .A(n14176), .ZN(n14173) );
  INV_X1 U7996 ( .A(n14173), .ZN(n14174) );
  INV_X1 U7997 ( .A(n6458), .ZN(n14175) );
  INV_X1 U7998 ( .A(n14175), .ZN(n14176) );
  BUF_X1 U7999 ( .A(n14179), .Z(n14177) );
  INV_X1 U8000 ( .A(n14181), .ZN(n14178) );
  INV_X1 U8001 ( .A(n14178), .ZN(n14179) );
  INV_X1 U8002 ( .A(n6457), .ZN(n14180) );
  INV_X1 U8003 ( .A(n14180), .ZN(n14181) );
  BUF_X1 U8004 ( .A(n14184), .Z(n14182) );
  INV_X1 U8005 ( .A(n14186), .ZN(n14183) );
  INV_X1 U8006 ( .A(n14183), .ZN(n14184) );
  INV_X1 U8007 ( .A(n6456), .ZN(n14185) );
  INV_X1 U8008 ( .A(n14185), .ZN(n14186) );
  BUF_X1 U8009 ( .A(n14189), .Z(n14187) );
  INV_X1 U8010 ( .A(n14191), .ZN(n14188) );
  INV_X1 U8011 ( .A(n14188), .ZN(n14189) );
  INV_X1 U8012 ( .A(n6455), .ZN(n14190) );
  INV_X1 U8013 ( .A(n14190), .ZN(n14191) );
  BUF_X1 U8014 ( .A(n14194), .Z(n14192) );
  INV_X1 U8015 ( .A(n14196), .ZN(n14193) );
  INV_X1 U8016 ( .A(n14193), .ZN(n14194) );
  INV_X1 U8017 ( .A(n6454), .ZN(n14195) );
  INV_X1 U8018 ( .A(n14195), .ZN(n14196) );
  BUF_X1 U8019 ( .A(n14199), .Z(n14197) );
  INV_X1 U8020 ( .A(n14201), .ZN(n14198) );
  INV_X1 U8021 ( .A(n14198), .ZN(n14199) );
  INV_X1 U8022 ( .A(n6453), .ZN(n14200) );
  INV_X1 U8023 ( .A(n14200), .ZN(n14201) );
  BUF_X1 U8024 ( .A(n14204), .Z(n14202) );
  INV_X1 U8025 ( .A(n14206), .ZN(n14203) );
  INV_X1 U8026 ( .A(n14203), .ZN(n14204) );
  INV_X1 U8027 ( .A(n6452), .ZN(n14205) );
  INV_X1 U8028 ( .A(n14205), .ZN(n14206) );
  BUF_X1 U8029 ( .A(n14209), .Z(n14207) );
  INV_X1 U8030 ( .A(n14211), .ZN(n14208) );
  INV_X1 U8031 ( .A(n14208), .ZN(n14209) );
  INV_X1 U8032 ( .A(n6451), .ZN(n14210) );
  INV_X1 U8033 ( .A(n14210), .ZN(n14211) );
  BUF_X1 U8034 ( .A(n14214), .Z(n14212) );
  INV_X1 U8035 ( .A(n14216), .ZN(n14213) );
  INV_X1 U8036 ( .A(n14213), .ZN(n14214) );
  INV_X1 U8037 ( .A(n6450), .ZN(n14215) );
  INV_X1 U8038 ( .A(n14215), .ZN(n14216) );
  INV_X1 U8039 ( .A(n1396), .ZN(n14246) );
  BUF_X1 U8040 ( .A(n14247), .Z(n14217) );
  INV_X1 U8041 ( .A(n6898), .ZN(n14218) );
  INV_X1 U8042 ( .A(n14218), .ZN(n14219) );
  INV_X1 U8043 ( .A(n1395), .ZN(n14253) );
  BUF_X1 U8044 ( .A(n14254), .Z(n14220) );
  INV_X1 U8045 ( .A(n6899), .ZN(n14221) );
  INV_X1 U8046 ( .A(n14221), .ZN(n14222) );
  INV_X1 U8047 ( .A(n1394), .ZN(n14260) );
  BUF_X1 U8048 ( .A(n14261), .Z(n14223) );
  INV_X1 U8049 ( .A(n6900), .ZN(n14224) );
  INV_X1 U8050 ( .A(n14224), .ZN(n14225) );
  INV_X1 U8051 ( .A(n1393), .ZN(n14267) );
  BUF_X1 U8052 ( .A(n14268), .Z(n14226) );
  INV_X1 U8053 ( .A(n6901), .ZN(n14227) );
  INV_X1 U8054 ( .A(n14227), .ZN(n14228) );
  INV_X1 U8055 ( .A(n1392), .ZN(n14274) );
  BUF_X1 U8056 ( .A(n14275), .Z(n14229) );
  INV_X1 U8057 ( .A(n6902), .ZN(n14230) );
  INV_X1 U8058 ( .A(n14230), .ZN(n14231) );
  INV_X1 U8059 ( .A(n1391), .ZN(n14281) );
  BUF_X1 U8060 ( .A(n14282), .Z(n14232) );
  INV_X1 U8061 ( .A(n6903), .ZN(n14233) );
  INV_X1 U8062 ( .A(n14233), .ZN(n14234) );
  INV_X1 U8063 ( .A(n1390), .ZN(n14288) );
  BUF_X1 U8064 ( .A(n14289), .Z(n14235) );
  INV_X1 U8065 ( .A(n6904), .ZN(n14236) );
  INV_X1 U8066 ( .A(n14236), .ZN(n14237) );
  INV_X1 U8067 ( .A(n1389), .ZN(n14295) );
  BUF_X1 U8068 ( .A(n14296), .Z(n14238) );
  INV_X1 U8069 ( .A(n6905), .ZN(n14239) );
  INV_X1 U8070 ( .A(n14239), .ZN(n14240) );
  BUF_X1 U8071 ( .A(n14243), .Z(n14241) );
  INV_X1 U8072 ( .A(n14245), .ZN(n14242) );
  INV_X1 U8073 ( .A(n14242), .ZN(n14243) );
  INV_X1 U8074 ( .A(n74090), .ZN(n14244) );
  INV_X1 U8075 ( .A(n14244), .ZN(n14245) );
  INV_X1 U8076 ( .A(n14246), .ZN(n14247) );
  BUF_X1 U8077 ( .A(n14250), .Z(n14248) );
  INV_X1 U8078 ( .A(n14252), .ZN(n14249) );
  INV_X1 U8079 ( .A(n14249), .ZN(n14250) );
  INV_X1 U8080 ( .A(n74080), .ZN(n14251) );
  INV_X1 U8081 ( .A(n14251), .ZN(n14252) );
  INV_X1 U8082 ( .A(n14253), .ZN(n14254) );
  BUF_X1 U8083 ( .A(n14257), .Z(n14255) );
  INV_X1 U8084 ( .A(n14259), .ZN(n14256) );
  INV_X1 U8085 ( .A(n14256), .ZN(n14257) );
  INV_X1 U8086 ( .A(n74070), .ZN(n14258) );
  INV_X1 U8087 ( .A(n14258), .ZN(n14259) );
  INV_X1 U8088 ( .A(n14260), .ZN(n14261) );
  BUF_X1 U8089 ( .A(n14264), .Z(n14262) );
  INV_X1 U8090 ( .A(n14266), .ZN(n14263) );
  INV_X1 U8091 ( .A(n14263), .ZN(n14264) );
  INV_X1 U8092 ( .A(n74060), .ZN(n14265) );
  INV_X1 U8093 ( .A(n14265), .ZN(n14266) );
  INV_X1 U8094 ( .A(n14267), .ZN(n14268) );
  BUF_X1 U8095 ( .A(n14271), .Z(n14269) );
  INV_X1 U8096 ( .A(n14273), .ZN(n14270) );
  INV_X1 U8097 ( .A(n14270), .ZN(n14271) );
  INV_X1 U8098 ( .A(n74050), .ZN(n14272) );
  INV_X1 U8099 ( .A(n14272), .ZN(n14273) );
  INV_X1 U8100 ( .A(n14274), .ZN(n14275) );
  BUF_X1 U8101 ( .A(n14278), .Z(n14276) );
  INV_X1 U8102 ( .A(n14280), .ZN(n14277) );
  INV_X1 U8103 ( .A(n14277), .ZN(n14278) );
  INV_X1 U8104 ( .A(n74040), .ZN(n14279) );
  INV_X1 U8105 ( .A(n14279), .ZN(n14280) );
  INV_X1 U8106 ( .A(n14281), .ZN(n14282) );
  BUF_X1 U8107 ( .A(n14285), .Z(n14283) );
  INV_X1 U8108 ( .A(n14287), .ZN(n14284) );
  INV_X1 U8109 ( .A(n14284), .ZN(n14285) );
  INV_X1 U8110 ( .A(n74030), .ZN(n14286) );
  INV_X1 U8111 ( .A(n14286), .ZN(n14287) );
  INV_X1 U8112 ( .A(n14288), .ZN(n14289) );
  BUF_X1 U8113 ( .A(n14292), .Z(n14290) );
  INV_X1 U8114 ( .A(n14294), .ZN(n14291) );
  INV_X1 U8115 ( .A(n14291), .ZN(n14292) );
  INV_X1 U8116 ( .A(n74020), .ZN(n14293) );
  INV_X1 U8117 ( .A(n14293), .ZN(n14294) );
  INV_X1 U8118 ( .A(n14295), .ZN(n14296) );
  BUF_X1 U8119 ( .A(n14299), .Z(n14297) );
  INV_X1 U8120 ( .A(n14301), .ZN(n14298) );
  INV_X1 U8121 ( .A(n14298), .ZN(n14299) );
  INV_X1 U8122 ( .A(n74010), .ZN(n14300) );
  INV_X1 U8123 ( .A(n14300), .ZN(n14301) );
  BUF_X1 U8124 ( .A(n14304), .Z(n14302) );
  INV_X1 U8125 ( .A(n14306), .ZN(n14303) );
  INV_X1 U8126 ( .A(n14303), .ZN(n14304) );
  INV_X1 U8127 ( .A(n74000), .ZN(n14305) );
  INV_X1 U8128 ( .A(n14305), .ZN(n14306) );
  BUF_X1 U8129 ( .A(n14309), .Z(n14307) );
  INV_X1 U8130 ( .A(n14311), .ZN(n14308) );
  INV_X1 U8131 ( .A(n14308), .ZN(n14309) );
  INV_X1 U8132 ( .A(n73990), .ZN(n14310) );
  INV_X1 U8133 ( .A(n14310), .ZN(n14311) );
  BUF_X1 U8134 ( .A(n14314), .Z(n14312) );
  INV_X1 U8135 ( .A(n14316), .ZN(n14313) );
  INV_X1 U8136 ( .A(n14313), .ZN(n14314) );
  INV_X1 U8137 ( .A(n73980), .ZN(n14315) );
  INV_X1 U8138 ( .A(n14315), .ZN(n14316) );
  BUF_X1 U8139 ( .A(n14319), .Z(n14317) );
  INV_X1 U8140 ( .A(n14321), .ZN(n14318) );
  INV_X1 U8141 ( .A(n14318), .ZN(n14319) );
  INV_X1 U8142 ( .A(n73970), .ZN(n14320) );
  INV_X1 U8143 ( .A(n14320), .ZN(n14321) );
  BUF_X1 U8144 ( .A(n14324), .Z(n14322) );
  INV_X1 U8145 ( .A(n14326), .ZN(n14323) );
  INV_X1 U8146 ( .A(n14323), .ZN(n14324) );
  INV_X1 U8147 ( .A(n73960), .ZN(n14325) );
  INV_X1 U8148 ( .A(n14325), .ZN(n14326) );
  BUF_X1 U8149 ( .A(n14329), .Z(n14327) );
  INV_X1 U8150 ( .A(n14331), .ZN(n14328) );
  INV_X1 U8151 ( .A(n14328), .ZN(n14329) );
  INV_X1 U8152 ( .A(n73950), .ZN(n14330) );
  INV_X1 U8153 ( .A(n14330), .ZN(n14331) );
  BUF_X1 U8154 ( .A(n14334), .Z(n14332) );
  INV_X1 U8155 ( .A(n14336), .ZN(n14333) );
  INV_X1 U8156 ( .A(n14333), .ZN(n14334) );
  INV_X1 U8157 ( .A(n73940), .ZN(n14335) );
  INV_X1 U8158 ( .A(n14335), .ZN(n14336) );
  BUF_X1 U8159 ( .A(n14339), .Z(n14337) );
  INV_X1 U8160 ( .A(n14341), .ZN(n14338) );
  INV_X1 U8161 ( .A(n14338), .ZN(n14339) );
  INV_X1 U8162 ( .A(n73930), .ZN(n14340) );
  INV_X1 U8163 ( .A(n14340), .ZN(n14341) );
  BUF_X1 U8164 ( .A(n14344), .Z(n14342) );
  INV_X1 U8165 ( .A(n14346), .ZN(n14343) );
  INV_X1 U8166 ( .A(n14343), .ZN(n14344) );
  INV_X1 U8167 ( .A(n7392), .ZN(n14345) );
  INV_X1 U8168 ( .A(n14345), .ZN(n14346) );
  BUF_X1 U8169 ( .A(n14349), .Z(n14347) );
  INV_X1 U8170 ( .A(n14351), .ZN(n14348) );
  INV_X1 U8171 ( .A(n14348), .ZN(n14349) );
  INV_X1 U8172 ( .A(n7391), .ZN(n14350) );
  INV_X1 U8173 ( .A(n14350), .ZN(n14351) );
  BUF_X1 U8174 ( .A(n14354), .Z(n14352) );
  INV_X1 U8175 ( .A(n14356), .ZN(n14353) );
  INV_X1 U8176 ( .A(n14353), .ZN(n14354) );
  INV_X1 U8177 ( .A(n7390), .ZN(n14355) );
  INV_X1 U8178 ( .A(n14355), .ZN(n14356) );
  BUF_X1 U8179 ( .A(n14359), .Z(n14357) );
  INV_X1 U8180 ( .A(n14361), .ZN(n14358) );
  INV_X1 U8181 ( .A(n14358), .ZN(n14359) );
  INV_X1 U8182 ( .A(n7389), .ZN(n14360) );
  INV_X1 U8183 ( .A(n14360), .ZN(n14361) );
  BUF_X1 U8184 ( .A(n14364), .Z(n14362) );
  INV_X1 U8185 ( .A(n14366), .ZN(n14363) );
  INV_X1 U8186 ( .A(n14363), .ZN(n14364) );
  INV_X1 U8187 ( .A(n7388), .ZN(n14365) );
  INV_X1 U8188 ( .A(n14365), .ZN(n14366) );
  BUF_X1 U8189 ( .A(n14369), .Z(n14367) );
  INV_X1 U8190 ( .A(n14371), .ZN(n14368) );
  INV_X1 U8191 ( .A(n14368), .ZN(n14369) );
  INV_X1 U8192 ( .A(n7387), .ZN(n14370) );
  INV_X1 U8193 ( .A(n14370), .ZN(n14371) );
  BUF_X1 U8194 ( .A(n14374), .Z(n14372) );
  INV_X1 U8195 ( .A(n14376), .ZN(n14373) );
  INV_X1 U8196 ( .A(n14373), .ZN(n14374) );
  INV_X1 U8197 ( .A(n7386), .ZN(n14375) );
  INV_X1 U8198 ( .A(n14375), .ZN(n14376) );
  BUF_X1 U8199 ( .A(n14379), .Z(n14377) );
  INV_X1 U8200 ( .A(n14381), .ZN(n14378) );
  INV_X1 U8201 ( .A(n14378), .ZN(n14379) );
  INV_X1 U8202 ( .A(n7385), .ZN(n14380) );
  INV_X1 U8203 ( .A(n14380), .ZN(n14381) );
  BUF_X1 U8204 ( .A(n14384), .Z(n14382) );
  INV_X1 U8205 ( .A(n14386), .ZN(n14383) );
  INV_X1 U8206 ( .A(n14383), .ZN(n14384) );
  INV_X1 U8207 ( .A(n7384), .ZN(n14385) );
  INV_X1 U8208 ( .A(n14385), .ZN(n14386) );
  BUF_X1 U8209 ( .A(n14389), .Z(n14387) );
  INV_X1 U8210 ( .A(n14391), .ZN(n14388) );
  INV_X1 U8211 ( .A(n14388), .ZN(n14389) );
  INV_X1 U8212 ( .A(n7383), .ZN(n14390) );
  INV_X1 U8213 ( .A(n14390), .ZN(n14391) );
  BUF_X1 U8214 ( .A(n14394), .Z(n14392) );
  INV_X1 U8215 ( .A(n14396), .ZN(n14393) );
  INV_X1 U8216 ( .A(n14393), .ZN(n14394) );
  INV_X1 U8217 ( .A(n7382), .ZN(n14395) );
  INV_X1 U8218 ( .A(n14395), .ZN(n14396) );
  BUF_X1 U8219 ( .A(n14399), .Z(n14397) );
  INV_X1 U8220 ( .A(n14401), .ZN(n14398) );
  INV_X1 U8221 ( .A(n14398), .ZN(n14399) );
  INV_X1 U8222 ( .A(n7381), .ZN(n14400) );
  INV_X1 U8223 ( .A(n14400), .ZN(n14401) );
  BUF_X1 U8224 ( .A(n14404), .Z(n14402) );
  INV_X1 U8225 ( .A(n14406), .ZN(n14403) );
  INV_X1 U8226 ( .A(n14403), .ZN(n14404) );
  INV_X1 U8227 ( .A(n7380), .ZN(n14405) );
  INV_X1 U8228 ( .A(n14405), .ZN(n14406) );
  BUF_X1 U8229 ( .A(n14409), .Z(n14407) );
  INV_X1 U8230 ( .A(n14411), .ZN(n14408) );
  INV_X1 U8231 ( .A(n14408), .ZN(n14409) );
  INV_X1 U8232 ( .A(n7379), .ZN(n14410) );
  INV_X1 U8233 ( .A(n14410), .ZN(n14411) );
  BUF_X1 U8234 ( .A(n14414), .Z(n14412) );
  INV_X1 U8235 ( .A(n14416), .ZN(n14413) );
  INV_X1 U8236 ( .A(n14413), .ZN(n14414) );
  INV_X1 U8237 ( .A(n7378), .ZN(n14415) );
  INV_X1 U8238 ( .A(n14415), .ZN(n14416) );
  BUF_X1 U8239 ( .A(n14419), .Z(n14417) );
  INV_X1 U8240 ( .A(n14421), .ZN(n14418) );
  INV_X1 U8241 ( .A(n14418), .ZN(n14419) );
  INV_X1 U8242 ( .A(n7377), .ZN(n14420) );
  INV_X1 U8243 ( .A(n14420), .ZN(n14421) );
  BUF_X1 U8244 ( .A(n14424), .Z(n14422) );
  INV_X1 U8245 ( .A(n14426), .ZN(n14423) );
  INV_X1 U8246 ( .A(n14423), .ZN(n14424) );
  INV_X1 U8247 ( .A(n7376), .ZN(n14425) );
  INV_X1 U8248 ( .A(n14425), .ZN(n14426) );
  BUF_X1 U8249 ( .A(n14429), .Z(n14427) );
  INV_X1 U8250 ( .A(n14431), .ZN(n14428) );
  INV_X1 U8251 ( .A(n14428), .ZN(n14429) );
  INV_X1 U8252 ( .A(n73750), .ZN(n14430) );
  INV_X1 U8253 ( .A(n14430), .ZN(n14431) );
  BUF_X1 U8254 ( .A(n14434), .Z(n14432) );
  INV_X1 U8255 ( .A(n14436), .ZN(n14433) );
  INV_X1 U8256 ( .A(n14433), .ZN(n14434) );
  INV_X1 U8257 ( .A(n73740), .ZN(n14435) );
  INV_X1 U8258 ( .A(n14435), .ZN(n14436) );
  BUF_X1 U8259 ( .A(n14439), .Z(n14437) );
  INV_X1 U8260 ( .A(n14441), .ZN(n14438) );
  INV_X1 U8261 ( .A(n14438), .ZN(n14439) );
  INV_X1 U8262 ( .A(n73730), .ZN(n14440) );
  INV_X1 U8263 ( .A(n14440), .ZN(n14441) );
  BUF_X1 U8264 ( .A(n14444), .Z(n14442) );
  INV_X1 U8265 ( .A(n14446), .ZN(n14443) );
  INV_X1 U8266 ( .A(n14443), .ZN(n14444) );
  INV_X1 U8267 ( .A(n73720), .ZN(n14445) );
  INV_X1 U8268 ( .A(n14445), .ZN(n14446) );
  BUF_X1 U8269 ( .A(n14449), .Z(n14447) );
  INV_X1 U8270 ( .A(n14451), .ZN(n14448) );
  INV_X1 U8271 ( .A(n14448), .ZN(n14449) );
  INV_X1 U8272 ( .A(n73710), .ZN(n14450) );
  INV_X1 U8273 ( .A(n14450), .ZN(n14451) );
  BUF_X1 U8274 ( .A(n14454), .Z(n14452) );
  INV_X1 U8275 ( .A(n14456), .ZN(n14453) );
  INV_X1 U8276 ( .A(n14453), .ZN(n14454) );
  INV_X1 U8277 ( .A(n73700), .ZN(n14455) );
  INV_X1 U8278 ( .A(n14455), .ZN(n14456) );
  BUF_X1 U8279 ( .A(n14459), .Z(n14457) );
  INV_X1 U8280 ( .A(n14461), .ZN(n14458) );
  INV_X1 U8281 ( .A(n14458), .ZN(n14459) );
  INV_X1 U8282 ( .A(n73690), .ZN(n14460) );
  INV_X1 U8283 ( .A(n14460), .ZN(n14461) );
  BUF_X1 U8284 ( .A(n14464), .Z(n14462) );
  INV_X1 U8285 ( .A(n14466), .ZN(n14463) );
  INV_X1 U8286 ( .A(n14463), .ZN(n14464) );
  INV_X1 U8287 ( .A(n73680), .ZN(n14465) );
  INV_X1 U8288 ( .A(n14465), .ZN(n14466) );
  BUF_X1 U8289 ( .A(n14469), .Z(n14467) );
  INV_X1 U8290 ( .A(n14471), .ZN(n14468) );
  INV_X1 U8291 ( .A(n14468), .ZN(n14469) );
  INV_X1 U8292 ( .A(n73670), .ZN(n14470) );
  INV_X1 U8293 ( .A(n14470), .ZN(n14471) );
  BUF_X1 U8294 ( .A(n14474), .Z(n14472) );
  INV_X1 U8295 ( .A(n14476), .ZN(n14473) );
  INV_X1 U8296 ( .A(n14473), .ZN(n14474) );
  INV_X1 U8297 ( .A(n73660), .ZN(n14475) );
  INV_X1 U8298 ( .A(n14475), .ZN(n14476) );
  BUF_X1 U8299 ( .A(n14479), .Z(n14477) );
  INV_X1 U8300 ( .A(n14481), .ZN(n14478) );
  INV_X1 U8301 ( .A(n14478), .ZN(n14479) );
  INV_X1 U8302 ( .A(n73650), .ZN(n14480) );
  INV_X1 U8303 ( .A(n14480), .ZN(n14481) );
  BUF_X1 U8304 ( .A(n14484), .Z(n14482) );
  INV_X1 U8305 ( .A(n14486), .ZN(n14483) );
  INV_X1 U8306 ( .A(n14483), .ZN(n14484) );
  INV_X1 U8307 ( .A(n73640), .ZN(n14485) );
  INV_X1 U8308 ( .A(n14485), .ZN(n14486) );
  BUF_X1 U8309 ( .A(n14489), .Z(n14487) );
  INV_X1 U8310 ( .A(n14491), .ZN(n14488) );
  INV_X1 U8311 ( .A(n14488), .ZN(n14489) );
  INV_X1 U8312 ( .A(n73630), .ZN(n14490) );
  INV_X1 U8313 ( .A(n14490), .ZN(n14491) );
  BUF_X1 U8314 ( .A(n14494), .Z(n14492) );
  INV_X1 U8315 ( .A(n14496), .ZN(n14493) );
  INV_X1 U8316 ( .A(n14493), .ZN(n14494) );
  INV_X1 U8317 ( .A(n73620), .ZN(n14495) );
  INV_X1 U8318 ( .A(n14495), .ZN(n14496) );
  BUF_X1 U8319 ( .A(n14499), .Z(n14497) );
  INV_X1 U8320 ( .A(n14501), .ZN(n14498) );
  INV_X1 U8321 ( .A(n14498), .ZN(n14499) );
  INV_X1 U8322 ( .A(n73610), .ZN(n14500) );
  INV_X1 U8323 ( .A(n14500), .ZN(n14501) );
  BUF_X1 U8324 ( .A(n14504), .Z(n14502) );
  INV_X1 U8325 ( .A(n14506), .ZN(n14503) );
  INV_X1 U8326 ( .A(n14503), .ZN(n14504) );
  INV_X1 U8327 ( .A(n73600), .ZN(n14505) );
  INV_X1 U8328 ( .A(n14505), .ZN(n14506) );
  BUF_X1 U8329 ( .A(n14509), .Z(n14507) );
  INV_X1 U8330 ( .A(n14511), .ZN(n14508) );
  INV_X1 U8331 ( .A(n14508), .ZN(n14509) );
  INV_X1 U8332 ( .A(n7359), .ZN(n14510) );
  INV_X1 U8333 ( .A(n14510), .ZN(n14511) );
  BUF_X1 U8334 ( .A(n14514), .Z(n14512) );
  INV_X1 U8335 ( .A(n14516), .ZN(n14513) );
  INV_X1 U8336 ( .A(n14513), .ZN(n14514) );
  INV_X1 U8337 ( .A(n7358), .ZN(n14515) );
  INV_X1 U8338 ( .A(n14515), .ZN(n14516) );
  BUF_X1 U8339 ( .A(n14519), .Z(n14517) );
  INV_X1 U8340 ( .A(n14521), .ZN(n14518) );
  INV_X1 U8341 ( .A(n14518), .ZN(n14519) );
  INV_X1 U8342 ( .A(n7357), .ZN(n14520) );
  INV_X1 U8343 ( .A(n14520), .ZN(n14521) );
  BUF_X1 U8344 ( .A(n14524), .Z(n14522) );
  INV_X1 U8345 ( .A(n14526), .ZN(n14523) );
  INV_X1 U8346 ( .A(n14523), .ZN(n14524) );
  INV_X1 U8347 ( .A(n7356), .ZN(n14525) );
  INV_X1 U8348 ( .A(n14525), .ZN(n14526) );
  BUF_X1 U8349 ( .A(n14529), .Z(n14527) );
  INV_X1 U8350 ( .A(n14531), .ZN(n14528) );
  INV_X1 U8351 ( .A(n14528), .ZN(n14529) );
  INV_X1 U8352 ( .A(n7355), .ZN(n14530) );
  INV_X1 U8353 ( .A(n14530), .ZN(n14531) );
  BUF_X1 U8354 ( .A(n14534), .Z(n14532) );
  INV_X1 U8355 ( .A(n14536), .ZN(n14533) );
  INV_X1 U8356 ( .A(n14533), .ZN(n14534) );
  INV_X1 U8357 ( .A(n7354), .ZN(n14535) );
  INV_X1 U8358 ( .A(n14535), .ZN(n14536) );
  INV_X1 U8359 ( .A(n1340), .ZN(n14566) );
  BUF_X1 U8360 ( .A(n14567), .Z(n14537) );
  INV_X1 U8361 ( .A(n7353), .ZN(n14538) );
  INV_X1 U8362 ( .A(n14538), .ZN(n14539) );
  INV_X1 U8363 ( .A(n1339), .ZN(n14573) );
  BUF_X1 U8364 ( .A(n14574), .Z(n14540) );
  INV_X1 U8365 ( .A(n7352), .ZN(n14541) );
  INV_X1 U8366 ( .A(n14541), .ZN(n14542) );
  INV_X1 U8367 ( .A(n1338), .ZN(n14580) );
  BUF_X1 U8368 ( .A(n14581), .Z(n14543) );
  INV_X1 U8369 ( .A(n7351), .ZN(n14544) );
  INV_X1 U8370 ( .A(n14544), .ZN(n14545) );
  INV_X1 U8371 ( .A(n1337), .ZN(n14587) );
  BUF_X1 U8372 ( .A(n14588), .Z(n14546) );
  INV_X1 U8373 ( .A(n7350), .ZN(n14547) );
  INV_X1 U8374 ( .A(n14547), .ZN(n14548) );
  INV_X1 U8375 ( .A(n1336), .ZN(n14594) );
  BUF_X1 U8376 ( .A(n14595), .Z(n14549) );
  INV_X1 U8377 ( .A(n7349), .ZN(n14550) );
  INV_X1 U8378 ( .A(n14550), .ZN(n14551) );
  INV_X1 U8379 ( .A(n1335), .ZN(n14601) );
  BUF_X1 U8380 ( .A(n14602), .Z(n14552) );
  INV_X1 U8381 ( .A(n7348), .ZN(n14553) );
  INV_X1 U8382 ( .A(n14553), .ZN(n14554) );
  INV_X1 U8383 ( .A(n1334), .ZN(n14608) );
  BUF_X1 U8384 ( .A(n14609), .Z(n14555) );
  INV_X1 U8385 ( .A(n7347), .ZN(n14556) );
  INV_X1 U8386 ( .A(n14556), .ZN(n14557) );
  INV_X1 U8387 ( .A(n1333), .ZN(n14615) );
  BUF_X1 U8388 ( .A(n14616), .Z(n14558) );
  INV_X1 U8389 ( .A(n7346), .ZN(n14559) );
  INV_X1 U8390 ( .A(n14559), .ZN(n14560) );
  BUF_X1 U8391 ( .A(n14563), .Z(n14561) );
  INV_X1 U8392 ( .A(n14565), .ZN(n14562) );
  INV_X1 U8393 ( .A(n14562), .ZN(n14563) );
  INV_X1 U8394 ( .A(n7345), .ZN(n14564) );
  INV_X1 U8395 ( .A(n14564), .ZN(n14565) );
  INV_X1 U8396 ( .A(n14566), .ZN(n14567) );
  BUF_X1 U8397 ( .A(n14570), .Z(n14568) );
  INV_X1 U8398 ( .A(n14572), .ZN(n14569) );
  INV_X1 U8399 ( .A(n14569), .ZN(n14570) );
  INV_X1 U8400 ( .A(n7344), .ZN(n14571) );
  INV_X1 U8401 ( .A(n14571), .ZN(n14572) );
  INV_X1 U8402 ( .A(n14573), .ZN(n14574) );
  BUF_X1 U8403 ( .A(n14577), .Z(n14575) );
  INV_X1 U8404 ( .A(n14579), .ZN(n14576) );
  INV_X1 U8405 ( .A(n14576), .ZN(n14577) );
  INV_X1 U8406 ( .A(n7343), .ZN(n14578) );
  INV_X1 U8407 ( .A(n14578), .ZN(n14579) );
  INV_X1 U8408 ( .A(n14580), .ZN(n14581) );
  BUF_X1 U8409 ( .A(n14584), .Z(n14582) );
  INV_X1 U8410 ( .A(n14586), .ZN(n14583) );
  INV_X1 U8411 ( .A(n14583), .ZN(n14584) );
  INV_X1 U8412 ( .A(n7342), .ZN(n14585) );
  INV_X1 U8413 ( .A(n14585), .ZN(n14586) );
  INV_X1 U8414 ( .A(n14587), .ZN(n14588) );
  BUF_X1 U8415 ( .A(n14591), .Z(n14589) );
  INV_X1 U8416 ( .A(n14593), .ZN(n14590) );
  INV_X1 U8417 ( .A(n14590), .ZN(n14591) );
  INV_X1 U8418 ( .A(n7341), .ZN(n14592) );
  INV_X1 U8419 ( .A(n14592), .ZN(n14593) );
  INV_X1 U8420 ( .A(n14594), .ZN(n14595) );
  BUF_X1 U8421 ( .A(n14598), .Z(n14596) );
  INV_X1 U8422 ( .A(n14600), .ZN(n14597) );
  INV_X1 U8423 ( .A(n14597), .ZN(n14598) );
  INV_X1 U8424 ( .A(n7340), .ZN(n14599) );
  INV_X1 U8425 ( .A(n14599), .ZN(n14600) );
  INV_X1 U8426 ( .A(n14601), .ZN(n14602) );
  BUF_X1 U8427 ( .A(n14605), .Z(n14603) );
  INV_X1 U8428 ( .A(n14607), .ZN(n14604) );
  INV_X1 U8429 ( .A(n14604), .ZN(n14605) );
  INV_X1 U8430 ( .A(n7339), .ZN(n14606) );
  INV_X1 U8431 ( .A(n14606), .ZN(n14607) );
  INV_X1 U8432 ( .A(n14608), .ZN(n14609) );
  BUF_X1 U8433 ( .A(n14612), .Z(n14610) );
  INV_X1 U8434 ( .A(n14614), .ZN(n14611) );
  INV_X1 U8435 ( .A(n14611), .ZN(n14612) );
  INV_X1 U8436 ( .A(n7338), .ZN(n14613) );
  INV_X1 U8437 ( .A(n14613), .ZN(n14614) );
  INV_X1 U8438 ( .A(n14615), .ZN(n14616) );
  BUF_X1 U8439 ( .A(n14619), .Z(n14617) );
  INV_X1 U8440 ( .A(n14621), .ZN(n14618) );
  INV_X1 U8441 ( .A(n14618), .ZN(n14619) );
  INV_X1 U8442 ( .A(n7337), .ZN(n14620) );
  INV_X1 U8443 ( .A(n14620), .ZN(n14621) );
  BUF_X1 U8444 ( .A(n14624), .Z(n14622) );
  INV_X1 U8445 ( .A(n14626), .ZN(n14623) );
  INV_X1 U8446 ( .A(n14623), .ZN(n14624) );
  INV_X1 U8447 ( .A(n7336), .ZN(n14625) );
  INV_X1 U8448 ( .A(n14625), .ZN(n14626) );
  BUF_X1 U8449 ( .A(n14629), .Z(n14627) );
  INV_X1 U8450 ( .A(n14631), .ZN(n14628) );
  INV_X1 U8451 ( .A(n14628), .ZN(n14629) );
  INV_X1 U8452 ( .A(n7335), .ZN(n14630) );
  INV_X1 U8453 ( .A(n14630), .ZN(n14631) );
  BUF_X1 U8454 ( .A(n14634), .Z(n14632) );
  INV_X1 U8455 ( .A(n14636), .ZN(n14633) );
  INV_X1 U8456 ( .A(n14633), .ZN(n14634) );
  INV_X1 U8457 ( .A(n7334), .ZN(n14635) );
  INV_X1 U8458 ( .A(n14635), .ZN(n14636) );
  BUF_X1 U8459 ( .A(n14639), .Z(n14637) );
  INV_X1 U8460 ( .A(n14641), .ZN(n14638) );
  INV_X1 U8461 ( .A(n14638), .ZN(n14639) );
  INV_X1 U8462 ( .A(n7333), .ZN(n14640) );
  INV_X1 U8463 ( .A(n14640), .ZN(n14641) );
  BUF_X1 U8464 ( .A(n14644), .Z(n14642) );
  INV_X1 U8465 ( .A(n14646), .ZN(n14643) );
  INV_X1 U8466 ( .A(n14643), .ZN(n14644) );
  INV_X1 U8467 ( .A(n7332), .ZN(n14645) );
  INV_X1 U8468 ( .A(n14645), .ZN(n14646) );
  BUF_X1 U8469 ( .A(n14649), .Z(n14647) );
  INV_X1 U8470 ( .A(n14651), .ZN(n14648) );
  INV_X1 U8471 ( .A(n14648), .ZN(n14649) );
  INV_X1 U8472 ( .A(n7331), .ZN(n14650) );
  INV_X1 U8473 ( .A(n14650), .ZN(n14651) );
  BUF_X1 U8474 ( .A(n14654), .Z(n14652) );
  INV_X1 U8475 ( .A(n14656), .ZN(n14653) );
  INV_X1 U8476 ( .A(n14653), .ZN(n14654) );
  INV_X1 U8477 ( .A(n7330), .ZN(n14655) );
  INV_X1 U8478 ( .A(n14655), .ZN(n14656) );
  BUF_X1 U8479 ( .A(n14659), .Z(n14657) );
  INV_X1 U8480 ( .A(n14661), .ZN(n14658) );
  INV_X1 U8481 ( .A(n14658), .ZN(n14659) );
  INV_X1 U8482 ( .A(n7329), .ZN(n14660) );
  INV_X1 U8483 ( .A(n14660), .ZN(n14661) );
  BUF_X1 U8484 ( .A(n14664), .Z(n14662) );
  INV_X1 U8485 ( .A(n14666), .ZN(n14663) );
  INV_X1 U8486 ( .A(n14663), .ZN(n14664) );
  INV_X1 U8487 ( .A(n7328), .ZN(n14665) );
  INV_X1 U8488 ( .A(n14665), .ZN(n14666) );
  BUF_X1 U8489 ( .A(n14669), .Z(n14667) );
  INV_X1 U8490 ( .A(n14671), .ZN(n14668) );
  INV_X1 U8491 ( .A(n14668), .ZN(n14669) );
  INV_X1 U8492 ( .A(n7327), .ZN(n14670) );
  INV_X1 U8493 ( .A(n14670), .ZN(n14671) );
  BUF_X1 U8494 ( .A(n14674), .Z(n14672) );
  INV_X1 U8495 ( .A(n14676), .ZN(n14673) );
  INV_X1 U8496 ( .A(n14673), .ZN(n14674) );
  INV_X1 U8497 ( .A(n7326), .ZN(n14675) );
  INV_X1 U8498 ( .A(n14675), .ZN(n14676) );
  BUF_X1 U8499 ( .A(n14679), .Z(n14677) );
  INV_X1 U8500 ( .A(n14681), .ZN(n14678) );
  INV_X1 U8501 ( .A(n14678), .ZN(n14679) );
  INV_X1 U8502 ( .A(n7325), .ZN(n14680) );
  INV_X1 U8503 ( .A(n14680), .ZN(n14681) );
  BUF_X1 U8504 ( .A(n14684), .Z(n14682) );
  INV_X1 U8505 ( .A(n14686), .ZN(n14683) );
  INV_X1 U8506 ( .A(n14683), .ZN(n14684) );
  INV_X1 U8507 ( .A(n73240), .ZN(n14685) );
  INV_X1 U8508 ( .A(n14685), .ZN(n14686) );
  BUF_X1 U8509 ( .A(n14689), .Z(n14687) );
  INV_X1 U8510 ( .A(n14691), .ZN(n14688) );
  INV_X1 U8511 ( .A(n14688), .ZN(n14689) );
  INV_X1 U8512 ( .A(n73230), .ZN(n14690) );
  INV_X1 U8513 ( .A(n14690), .ZN(n14691) );
  BUF_X1 U8514 ( .A(n14694), .Z(n14692) );
  INV_X1 U8515 ( .A(n14696), .ZN(n14693) );
  INV_X1 U8516 ( .A(n14693), .ZN(n14694) );
  INV_X1 U8517 ( .A(n73220), .ZN(n14695) );
  INV_X1 U8518 ( .A(n14695), .ZN(n14696) );
  BUF_X1 U8519 ( .A(n14699), .Z(n14697) );
  INV_X1 U8520 ( .A(n14701), .ZN(n14698) );
  INV_X1 U8521 ( .A(n14698), .ZN(n14699) );
  INV_X1 U8522 ( .A(n73210), .ZN(n14700) );
  INV_X1 U8523 ( .A(n14700), .ZN(n14701) );
  BUF_X1 U8524 ( .A(n14704), .Z(n14702) );
  INV_X1 U8525 ( .A(n14706), .ZN(n14703) );
  INV_X1 U8526 ( .A(n14703), .ZN(n14704) );
  INV_X1 U8527 ( .A(n73200), .ZN(n14705) );
  INV_X1 U8528 ( .A(n14705), .ZN(n14706) );
  BUF_X1 U8529 ( .A(n14709), .Z(n14707) );
  INV_X1 U8530 ( .A(n14711), .ZN(n14708) );
  INV_X1 U8531 ( .A(n14708), .ZN(n14709) );
  INV_X1 U8532 ( .A(n73190), .ZN(n14710) );
  INV_X1 U8533 ( .A(n14710), .ZN(n14711) );
  BUF_X1 U8534 ( .A(n14714), .Z(n14712) );
  INV_X1 U8535 ( .A(n14716), .ZN(n14713) );
  INV_X1 U8536 ( .A(n14713), .ZN(n14714) );
  INV_X1 U8537 ( .A(n73180), .ZN(n14715) );
  INV_X1 U8538 ( .A(n14715), .ZN(n14716) );
  BUF_X1 U8539 ( .A(n14719), .Z(n14717) );
  INV_X1 U8540 ( .A(n14721), .ZN(n14718) );
  INV_X1 U8541 ( .A(n14718), .ZN(n14719) );
  INV_X1 U8542 ( .A(n73170), .ZN(n14720) );
  INV_X1 U8543 ( .A(n14720), .ZN(n14721) );
  BUF_X1 U8544 ( .A(n14724), .Z(n14722) );
  INV_X1 U8545 ( .A(n14726), .ZN(n14723) );
  INV_X1 U8546 ( .A(n14723), .ZN(n14724) );
  INV_X1 U8547 ( .A(n73160), .ZN(n14725) );
  INV_X1 U8548 ( .A(n14725), .ZN(n14726) );
  BUF_X1 U8549 ( .A(n14729), .Z(n14727) );
  INV_X1 U8550 ( .A(n14731), .ZN(n14728) );
  INV_X1 U8551 ( .A(n14728), .ZN(n14729) );
  INV_X1 U8552 ( .A(n73150), .ZN(n14730) );
  INV_X1 U8553 ( .A(n14730), .ZN(n14731) );
  BUF_X1 U8554 ( .A(n14734), .Z(n14732) );
  INV_X1 U8555 ( .A(n14736), .ZN(n14733) );
  INV_X1 U8556 ( .A(n14733), .ZN(n14734) );
  INV_X1 U8557 ( .A(n73140), .ZN(n14735) );
  INV_X1 U8558 ( .A(n14735), .ZN(n14736) );
  BUF_X1 U8559 ( .A(n14739), .Z(n14737) );
  INV_X1 U8560 ( .A(n14741), .ZN(n14738) );
  INV_X1 U8561 ( .A(n14738), .ZN(n14739) );
  INV_X1 U8562 ( .A(n73130), .ZN(n14740) );
  INV_X1 U8563 ( .A(n14740), .ZN(n14741) );
  BUF_X1 U8564 ( .A(n14744), .Z(n14742) );
  INV_X1 U8565 ( .A(n14746), .ZN(n14743) );
  INV_X1 U8566 ( .A(n14743), .ZN(n14744) );
  INV_X1 U8567 ( .A(n73120), .ZN(n14745) );
  INV_X1 U8568 ( .A(n14745), .ZN(n14746) );
  BUF_X1 U8569 ( .A(n14749), .Z(n14747) );
  INV_X1 U8570 ( .A(n14751), .ZN(n14748) );
  INV_X1 U8571 ( .A(n14748), .ZN(n14749) );
  INV_X1 U8572 ( .A(n73110), .ZN(n14750) );
  INV_X1 U8573 ( .A(n14750), .ZN(n14751) );
  BUF_X1 U8574 ( .A(n14754), .Z(n14752) );
  INV_X1 U8575 ( .A(n14756), .ZN(n14753) );
  INV_X1 U8576 ( .A(n14753), .ZN(n14754) );
  INV_X1 U8577 ( .A(n73100), .ZN(n14755) );
  INV_X1 U8578 ( .A(n14755), .ZN(n14756) );
  BUF_X1 U8579 ( .A(n14759), .Z(n14757) );
  INV_X1 U8580 ( .A(n14761), .ZN(n14758) );
  INV_X1 U8581 ( .A(n14758), .ZN(n14759) );
  INV_X1 U8582 ( .A(n73090), .ZN(n14760) );
  INV_X1 U8583 ( .A(n14760), .ZN(n14761) );
  BUF_X1 U8584 ( .A(n14764), .Z(n14762) );
  INV_X1 U8585 ( .A(n14766), .ZN(n14763) );
  INV_X1 U8586 ( .A(n14763), .ZN(n14764) );
  INV_X1 U8587 ( .A(n73080), .ZN(n14765) );
  INV_X1 U8588 ( .A(n14765), .ZN(n14766) );
  BUF_X1 U8589 ( .A(n14769), .Z(n14767) );
  INV_X1 U8590 ( .A(n14771), .ZN(n14768) );
  INV_X1 U8591 ( .A(n14768), .ZN(n14769) );
  INV_X1 U8592 ( .A(n73070), .ZN(n14770) );
  INV_X1 U8593 ( .A(n14770), .ZN(n14771) );
  BUF_X1 U8594 ( .A(n14774), .Z(n14772) );
  INV_X1 U8595 ( .A(n14776), .ZN(n14773) );
  INV_X1 U8596 ( .A(n14773), .ZN(n14774) );
  INV_X1 U8597 ( .A(n73060), .ZN(n14775) );
  INV_X1 U8598 ( .A(n14775), .ZN(n14776) );
  BUF_X1 U8599 ( .A(n14779), .Z(n14777) );
  INV_X1 U8600 ( .A(n14781), .ZN(n14778) );
  INV_X1 U8601 ( .A(n14778), .ZN(n14779) );
  INV_X1 U8602 ( .A(n73050), .ZN(n14780) );
  INV_X1 U8603 ( .A(n14780), .ZN(n14781) );
  BUF_X1 U8604 ( .A(n14784), .Z(n14782) );
  INV_X1 U8605 ( .A(n14786), .ZN(n14783) );
  INV_X1 U8606 ( .A(n14783), .ZN(n14784) );
  INV_X1 U8607 ( .A(n73040), .ZN(n14785) );
  INV_X1 U8608 ( .A(n14785), .ZN(n14786) );
  BUF_X1 U8609 ( .A(n14789), .Z(n14787) );
  INV_X1 U8610 ( .A(n14791), .ZN(n14788) );
  INV_X1 U8611 ( .A(n14788), .ZN(n14789) );
  INV_X1 U8612 ( .A(n7303), .ZN(n14790) );
  INV_X1 U8613 ( .A(n14790), .ZN(n14791) );
  BUF_X1 U8614 ( .A(n14794), .Z(n14792) );
  INV_X1 U8615 ( .A(n14796), .ZN(n14793) );
  INV_X1 U8616 ( .A(n14793), .ZN(n14794) );
  INV_X1 U8617 ( .A(n7302), .ZN(n14795) );
  INV_X1 U8618 ( .A(n14795), .ZN(n14796) );
  BUF_X1 U8619 ( .A(n14799), .Z(n14797) );
  INV_X1 U8620 ( .A(n14801), .ZN(n14798) );
  INV_X1 U8621 ( .A(n14798), .ZN(n14799) );
  INV_X1 U8622 ( .A(n7301), .ZN(n14800) );
  INV_X1 U8623 ( .A(n14800), .ZN(n14801) );
  BUF_X1 U8624 ( .A(n14804), .Z(n14802) );
  INV_X1 U8625 ( .A(n14806), .ZN(n14803) );
  INV_X1 U8626 ( .A(n14803), .ZN(n14804) );
  INV_X1 U8627 ( .A(n7300), .ZN(n14805) );
  INV_X1 U8628 ( .A(n14805), .ZN(n14806) );
  BUF_X1 U8629 ( .A(n14809), .Z(n14807) );
  INV_X1 U8630 ( .A(n14811), .ZN(n14808) );
  INV_X1 U8631 ( .A(n14808), .ZN(n14809) );
  INV_X1 U8632 ( .A(n7299), .ZN(n14810) );
  INV_X1 U8633 ( .A(n14810), .ZN(n14811) );
  BUF_X1 U8634 ( .A(n14814), .Z(n14812) );
  INV_X1 U8635 ( .A(n14816), .ZN(n14813) );
  INV_X1 U8636 ( .A(n14813), .ZN(n14814) );
  INV_X1 U8637 ( .A(n7298), .ZN(n14815) );
  INV_X1 U8638 ( .A(n14815), .ZN(n14816) );
  BUF_X1 U8639 ( .A(n14819), .Z(n14817) );
  INV_X1 U8640 ( .A(n14821), .ZN(n14818) );
  INV_X1 U8641 ( .A(n14818), .ZN(n14819) );
  INV_X1 U8642 ( .A(n7297), .ZN(n14820) );
  INV_X1 U8643 ( .A(n14820), .ZN(n14821) );
  BUF_X1 U8644 ( .A(n14824), .Z(n14822) );
  INV_X1 U8645 ( .A(n14826), .ZN(n14823) );
  INV_X1 U8646 ( .A(n14823), .ZN(n14824) );
  INV_X1 U8647 ( .A(n7296), .ZN(n14825) );
  INV_X1 U8648 ( .A(n14825), .ZN(n14826) );
  BUF_X1 U8649 ( .A(n14829), .Z(n14827) );
  INV_X1 U8650 ( .A(n14831), .ZN(n14828) );
  INV_X1 U8651 ( .A(n14828), .ZN(n14829) );
  INV_X1 U8652 ( .A(n7295), .ZN(n14830) );
  INV_X1 U8653 ( .A(n14830), .ZN(n14831) );
  BUF_X1 U8654 ( .A(n14834), .Z(n14832) );
  INV_X1 U8655 ( .A(n14836), .ZN(n14833) );
  INV_X1 U8656 ( .A(n14833), .ZN(n14834) );
  INV_X1 U8657 ( .A(n7294), .ZN(n14835) );
  INV_X1 U8658 ( .A(n14835), .ZN(n14836) );
  BUF_X1 U8659 ( .A(n14839), .Z(n14837) );
  INV_X1 U8660 ( .A(n14841), .ZN(n14838) );
  INV_X1 U8661 ( .A(n14838), .ZN(n14839) );
  INV_X1 U8662 ( .A(n7293), .ZN(n14840) );
  INV_X1 U8663 ( .A(n14840), .ZN(n14841) );
  BUF_X1 U8664 ( .A(n14844), .Z(n14842) );
  INV_X1 U8665 ( .A(n14846), .ZN(n14843) );
  INV_X1 U8666 ( .A(n14843), .ZN(n14844) );
  INV_X1 U8667 ( .A(n7292), .ZN(n14845) );
  INV_X1 U8668 ( .A(n14845), .ZN(n14846) );
  BUF_X1 U8669 ( .A(n14849), .Z(n14847) );
  INV_X1 U8670 ( .A(n14851), .ZN(n14848) );
  INV_X1 U8671 ( .A(n14848), .ZN(n14849) );
  INV_X1 U8672 ( .A(n7291), .ZN(n14850) );
  INV_X1 U8673 ( .A(n14850), .ZN(n14851) );
  BUF_X1 U8674 ( .A(n14854), .Z(n14852) );
  INV_X1 U8675 ( .A(n14856), .ZN(n14853) );
  INV_X1 U8676 ( .A(n14853), .ZN(n14854) );
  INV_X1 U8677 ( .A(n7290), .ZN(n14855) );
  INV_X1 U8678 ( .A(n14855), .ZN(n14856) );
  INV_X1 U8679 ( .A(n1284), .ZN(n14886) );
  BUF_X1 U8680 ( .A(n14887), .Z(n14857) );
  INV_X1 U8681 ( .A(n7289), .ZN(n14858) );
  INV_X1 U8682 ( .A(n14858), .ZN(n14859) );
  INV_X1 U8683 ( .A(n1283), .ZN(n14893) );
  BUF_X1 U8684 ( .A(n14894), .Z(n14860) );
  INV_X1 U8685 ( .A(n7288), .ZN(n14861) );
  INV_X1 U8686 ( .A(n14861), .ZN(n14862) );
  INV_X1 U8687 ( .A(n1282), .ZN(n14900) );
  BUF_X1 U8688 ( .A(n14901), .Z(n14863) );
  INV_X1 U8689 ( .A(n7287), .ZN(n14864) );
  INV_X1 U8690 ( .A(n14864), .ZN(n14865) );
  INV_X1 U8691 ( .A(n1281), .ZN(n14907) );
  BUF_X1 U8692 ( .A(n14908), .Z(n14866) );
  INV_X1 U8693 ( .A(n72860), .ZN(n14867) );
  INV_X1 U8694 ( .A(n14867), .ZN(n14868) );
  INV_X1 U8695 ( .A(n1280), .ZN(n14914) );
  BUF_X1 U8696 ( .A(n14915), .Z(n14869) );
  INV_X1 U8697 ( .A(n72850), .ZN(n14870) );
  INV_X1 U8698 ( .A(n14870), .ZN(n14871) );
  INV_X1 U8699 ( .A(n1279), .ZN(n14921) );
  BUF_X1 U8700 ( .A(n14922), .Z(n14872) );
  INV_X1 U8701 ( .A(n72840), .ZN(n14873) );
  INV_X1 U8702 ( .A(n14873), .ZN(n14874) );
  INV_X1 U8703 ( .A(n1278), .ZN(n14928) );
  BUF_X1 U8704 ( .A(n14929), .Z(n14875) );
  INV_X1 U8705 ( .A(n72830), .ZN(n14876) );
  INV_X1 U8706 ( .A(n14876), .ZN(n14877) );
  INV_X1 U8707 ( .A(n1277), .ZN(n14935) );
  BUF_X1 U8708 ( .A(n14936), .Z(n14878) );
  INV_X1 U8709 ( .A(n72820), .ZN(n14879) );
  INV_X1 U8710 ( .A(n14879), .ZN(n14880) );
  BUF_X1 U8711 ( .A(n14883), .Z(n14881) );
  INV_X1 U8712 ( .A(n14885), .ZN(n14882) );
  INV_X1 U8713 ( .A(n14882), .ZN(n14883) );
  INV_X1 U8714 ( .A(n72810), .ZN(n14884) );
  INV_X1 U8715 ( .A(n14884), .ZN(n14885) );
  INV_X1 U8716 ( .A(n14886), .ZN(n14887) );
  BUF_X1 U8717 ( .A(n14890), .Z(n14888) );
  INV_X1 U8718 ( .A(n14892), .ZN(n14889) );
  INV_X1 U8719 ( .A(n14889), .ZN(n14890) );
  INV_X1 U8720 ( .A(n72800), .ZN(n14891) );
  INV_X1 U8721 ( .A(n14891), .ZN(n14892) );
  INV_X1 U8722 ( .A(n14893), .ZN(n14894) );
  BUF_X1 U8723 ( .A(n14897), .Z(n14895) );
  INV_X1 U8724 ( .A(n14899), .ZN(n14896) );
  INV_X1 U8725 ( .A(n14896), .ZN(n14897) );
  INV_X1 U8726 ( .A(n72790), .ZN(n14898) );
  INV_X1 U8727 ( .A(n14898), .ZN(n14899) );
  INV_X1 U8728 ( .A(n14900), .ZN(n14901) );
  BUF_X1 U8729 ( .A(n14904), .Z(n14902) );
  INV_X1 U8730 ( .A(n14906), .ZN(n14903) );
  INV_X1 U8731 ( .A(n14903), .ZN(n14904) );
  INV_X1 U8732 ( .A(n72780), .ZN(n14905) );
  INV_X1 U8733 ( .A(n14905), .ZN(n14906) );
  INV_X1 U8734 ( .A(n14907), .ZN(n14908) );
  BUF_X1 U8735 ( .A(n14911), .Z(n14909) );
  INV_X1 U8736 ( .A(n14913), .ZN(n14910) );
  INV_X1 U8737 ( .A(n14910), .ZN(n14911) );
  INV_X1 U8738 ( .A(n72770), .ZN(n14912) );
  INV_X1 U8739 ( .A(n14912), .ZN(n14913) );
  INV_X1 U8740 ( .A(n14914), .ZN(n14915) );
  BUF_X1 U8741 ( .A(n14918), .Z(n14916) );
  INV_X1 U8742 ( .A(n14920), .ZN(n14917) );
  INV_X1 U8743 ( .A(n14917), .ZN(n14918) );
  INV_X1 U8744 ( .A(n72760), .ZN(n14919) );
  INV_X1 U8745 ( .A(n14919), .ZN(n14920) );
  INV_X1 U8746 ( .A(n14921), .ZN(n14922) );
  BUF_X1 U8747 ( .A(n14925), .Z(n14923) );
  INV_X1 U8748 ( .A(n14927), .ZN(n14924) );
  INV_X1 U8749 ( .A(n14924), .ZN(n14925) );
  INV_X1 U8750 ( .A(n72750), .ZN(n14926) );
  INV_X1 U8751 ( .A(n14926), .ZN(n14927) );
  INV_X1 U8752 ( .A(n14928), .ZN(n14929) );
  BUF_X1 U8753 ( .A(n14932), .Z(n14930) );
  INV_X1 U8754 ( .A(n14934), .ZN(n14931) );
  INV_X1 U8755 ( .A(n14931), .ZN(n14932) );
  INV_X1 U8756 ( .A(n72740), .ZN(n14933) );
  INV_X1 U8757 ( .A(n14933), .ZN(n14934) );
  INV_X1 U8758 ( .A(n14935), .ZN(n14936) );
  BUF_X1 U8759 ( .A(n14939), .Z(n14937) );
  INV_X1 U8760 ( .A(n14941), .ZN(n14938) );
  INV_X1 U8761 ( .A(n14938), .ZN(n14939) );
  INV_X1 U8762 ( .A(n72730), .ZN(n14940) );
  INV_X1 U8763 ( .A(n14940), .ZN(n14941) );
  BUF_X1 U8764 ( .A(n14944), .Z(n14942) );
  INV_X1 U8765 ( .A(n14946), .ZN(n14943) );
  INV_X1 U8766 ( .A(n14943), .ZN(n14944) );
  INV_X1 U8767 ( .A(n72720), .ZN(n14945) );
  INV_X1 U8768 ( .A(n14945), .ZN(n14946) );
  BUF_X1 U8769 ( .A(n14949), .Z(n14947) );
  INV_X1 U8770 ( .A(n14951), .ZN(n14948) );
  INV_X1 U8771 ( .A(n14948), .ZN(n14949) );
  INV_X1 U8772 ( .A(n72710), .ZN(n14950) );
  INV_X1 U8773 ( .A(n14950), .ZN(n14951) );
  BUF_X1 U8774 ( .A(n14954), .Z(n14952) );
  INV_X1 U8775 ( .A(n14956), .ZN(n14953) );
  INV_X1 U8776 ( .A(n14953), .ZN(n14954) );
  INV_X1 U8777 ( .A(n7270), .ZN(n14955) );
  INV_X1 U8778 ( .A(n14955), .ZN(n14956) );
  BUF_X1 U8779 ( .A(n14959), .Z(n14957) );
  INV_X1 U8780 ( .A(n14961), .ZN(n14958) );
  INV_X1 U8781 ( .A(n14958), .ZN(n14959) );
  INV_X1 U8782 ( .A(n7269), .ZN(n14960) );
  INV_X1 U8783 ( .A(n14960), .ZN(n14961) );
  BUF_X1 U8784 ( .A(n14964), .Z(n14962) );
  INV_X1 U8785 ( .A(n14966), .ZN(n14963) );
  INV_X1 U8786 ( .A(n14963), .ZN(n14964) );
  INV_X1 U8787 ( .A(n7268), .ZN(n14965) );
  INV_X1 U8788 ( .A(n14965), .ZN(n14966) );
  BUF_X1 U8789 ( .A(n14969), .Z(n14967) );
  INV_X1 U8790 ( .A(n14971), .ZN(n14968) );
  INV_X1 U8791 ( .A(n14968), .ZN(n14969) );
  INV_X1 U8792 ( .A(n72670), .ZN(n14970) );
  INV_X1 U8793 ( .A(n14970), .ZN(n14971) );
  BUF_X1 U8794 ( .A(n14974), .Z(n14972) );
  INV_X1 U8795 ( .A(n14976), .ZN(n14973) );
  INV_X1 U8796 ( .A(n14973), .ZN(n14974) );
  INV_X1 U8797 ( .A(n7266), .ZN(n14975) );
  INV_X1 U8798 ( .A(n14975), .ZN(n14976) );
  BUF_X1 U8799 ( .A(n14979), .Z(n14977) );
  INV_X1 U8800 ( .A(n14981), .ZN(n14978) );
  INV_X1 U8801 ( .A(n14978), .ZN(n14979) );
  INV_X1 U8802 ( .A(n7265), .ZN(n14980) );
  INV_X1 U8803 ( .A(n14980), .ZN(n14981) );
  BUF_X1 U8804 ( .A(n14984), .Z(n14982) );
  INV_X1 U8805 ( .A(n14986), .ZN(n14983) );
  INV_X1 U8806 ( .A(n14983), .ZN(n14984) );
  INV_X1 U8807 ( .A(n7264), .ZN(n14985) );
  INV_X1 U8808 ( .A(n14985), .ZN(n14986) );
  BUF_X1 U8809 ( .A(n14989), .Z(n14987) );
  INV_X1 U8810 ( .A(n14991), .ZN(n14988) );
  INV_X1 U8811 ( .A(n14988), .ZN(n14989) );
  INV_X1 U8812 ( .A(n7263), .ZN(n14990) );
  INV_X1 U8813 ( .A(n14990), .ZN(n14991) );
  BUF_X1 U8814 ( .A(n14994), .Z(n14992) );
  INV_X1 U8815 ( .A(n14996), .ZN(n14993) );
  INV_X1 U8816 ( .A(n14993), .ZN(n14994) );
  INV_X1 U8817 ( .A(n7262), .ZN(n14995) );
  INV_X1 U8818 ( .A(n14995), .ZN(n14996) );
  BUF_X1 U8819 ( .A(n14999), .Z(n14997) );
  INV_X1 U8820 ( .A(n15001), .ZN(n14998) );
  INV_X1 U8821 ( .A(n14998), .ZN(n14999) );
  INV_X1 U8822 ( .A(n7261), .ZN(n15000) );
  INV_X1 U8823 ( .A(n15000), .ZN(n15001) );
  BUF_X1 U8824 ( .A(n15004), .Z(n15002) );
  INV_X1 U8825 ( .A(n15006), .ZN(n15003) );
  INV_X1 U8826 ( .A(n15003), .ZN(n15004) );
  INV_X1 U8827 ( .A(n7260), .ZN(n15005) );
  INV_X1 U8828 ( .A(n15005), .ZN(n15006) );
  BUF_X1 U8829 ( .A(n15009), .Z(n15007) );
  INV_X1 U8830 ( .A(n15011), .ZN(n15008) );
  INV_X1 U8831 ( .A(n15008), .ZN(n15009) );
  INV_X1 U8832 ( .A(n7259), .ZN(n15010) );
  INV_X1 U8833 ( .A(n15010), .ZN(n15011) );
  BUF_X1 U8834 ( .A(n15014), .Z(n15012) );
  INV_X1 U8835 ( .A(n15016), .ZN(n15013) );
  INV_X1 U8836 ( .A(n15013), .ZN(n15014) );
  INV_X1 U8837 ( .A(n7258), .ZN(n15015) );
  INV_X1 U8838 ( .A(n15015), .ZN(n15016) );
  BUF_X1 U8839 ( .A(n15019), .Z(n15017) );
  INV_X1 U8840 ( .A(n15021), .ZN(n15018) );
  INV_X1 U8841 ( .A(n15018), .ZN(n15019) );
  INV_X1 U8842 ( .A(n7257), .ZN(n15020) );
  INV_X1 U8843 ( .A(n15020), .ZN(n15021) );
  BUF_X1 U8844 ( .A(n15024), .Z(n15022) );
  INV_X1 U8845 ( .A(n15026), .ZN(n15023) );
  INV_X1 U8846 ( .A(n15023), .ZN(n15024) );
  INV_X1 U8847 ( .A(n7256), .ZN(n15025) );
  INV_X1 U8848 ( .A(n15025), .ZN(n15026) );
  BUF_X1 U8849 ( .A(n15029), .Z(n15027) );
  INV_X1 U8850 ( .A(n15031), .ZN(n15028) );
  INV_X1 U8851 ( .A(n15028), .ZN(n15029) );
  INV_X1 U8852 ( .A(n7255), .ZN(n15030) );
  INV_X1 U8853 ( .A(n15030), .ZN(n15031) );
  BUF_X1 U8854 ( .A(n15034), .Z(n15032) );
  INV_X1 U8855 ( .A(n15036), .ZN(n15033) );
  INV_X1 U8856 ( .A(n15033), .ZN(n15034) );
  INV_X1 U8857 ( .A(n7254), .ZN(n15035) );
  INV_X1 U8858 ( .A(n15035), .ZN(n15036) );
  BUF_X1 U8859 ( .A(n15039), .Z(n15037) );
  INV_X1 U8860 ( .A(n15041), .ZN(n15038) );
  INV_X1 U8861 ( .A(n15038), .ZN(n15039) );
  INV_X1 U8862 ( .A(n7253), .ZN(n15040) );
  INV_X1 U8863 ( .A(n15040), .ZN(n15041) );
  BUF_X1 U8864 ( .A(n15044), .Z(n15042) );
  INV_X1 U8865 ( .A(n15046), .ZN(n15043) );
  INV_X1 U8866 ( .A(n15043), .ZN(n15044) );
  INV_X1 U8867 ( .A(n7252), .ZN(n15045) );
  INV_X1 U8868 ( .A(n15045), .ZN(n15046) );
  BUF_X1 U8869 ( .A(n15049), .Z(n15047) );
  INV_X1 U8870 ( .A(n15051), .ZN(n15048) );
  INV_X1 U8871 ( .A(n15048), .ZN(n15049) );
  INV_X1 U8872 ( .A(n7251), .ZN(n15050) );
  INV_X1 U8873 ( .A(n15050), .ZN(n15051) );
  BUF_X1 U8874 ( .A(n15054), .Z(n15052) );
  INV_X1 U8875 ( .A(n15056), .ZN(n15053) );
  INV_X1 U8876 ( .A(n15053), .ZN(n15054) );
  INV_X1 U8877 ( .A(n7250), .ZN(n15055) );
  INV_X1 U8878 ( .A(n15055), .ZN(n15056) );
  BUF_X1 U8879 ( .A(n15059), .Z(n15057) );
  INV_X1 U8880 ( .A(n15061), .ZN(n15058) );
  INV_X1 U8881 ( .A(n15058), .ZN(n15059) );
  INV_X1 U8882 ( .A(n7249), .ZN(n15060) );
  INV_X1 U8883 ( .A(n15060), .ZN(n15061) );
  BUF_X1 U8884 ( .A(n15064), .Z(n15062) );
  INV_X1 U8885 ( .A(n15066), .ZN(n15063) );
  INV_X1 U8886 ( .A(n15063), .ZN(n15064) );
  INV_X1 U8887 ( .A(n7248), .ZN(n15065) );
  INV_X1 U8888 ( .A(n15065), .ZN(n15066) );
  BUF_X1 U8889 ( .A(n15069), .Z(n15067) );
  INV_X1 U8890 ( .A(n15071), .ZN(n15068) );
  INV_X1 U8891 ( .A(n15068), .ZN(n15069) );
  INV_X1 U8892 ( .A(n7247), .ZN(n15070) );
  INV_X1 U8893 ( .A(n15070), .ZN(n15071) );
  BUF_X1 U8894 ( .A(n15074), .Z(n15072) );
  INV_X1 U8895 ( .A(n15076), .ZN(n15073) );
  INV_X1 U8896 ( .A(n15073), .ZN(n15074) );
  INV_X1 U8897 ( .A(n7246), .ZN(n15075) );
  INV_X1 U8898 ( .A(n15075), .ZN(n15076) );
  BUF_X1 U8899 ( .A(n15079), .Z(n15077) );
  INV_X1 U8900 ( .A(n15081), .ZN(n15078) );
  INV_X1 U8901 ( .A(n15078), .ZN(n15079) );
  INV_X1 U8902 ( .A(n7245), .ZN(n15080) );
  INV_X1 U8903 ( .A(n15080), .ZN(n15081) );
  BUF_X1 U8904 ( .A(n15084), .Z(n15082) );
  INV_X1 U8905 ( .A(n15086), .ZN(n15083) );
  INV_X1 U8906 ( .A(n15083), .ZN(n15084) );
  INV_X1 U8907 ( .A(n7244), .ZN(n15085) );
  INV_X1 U8908 ( .A(n15085), .ZN(n15086) );
  BUF_X1 U8909 ( .A(n15089), .Z(n15087) );
  INV_X1 U8910 ( .A(n15091), .ZN(n15088) );
  INV_X1 U8911 ( .A(n15088), .ZN(n15089) );
  INV_X1 U8912 ( .A(n7243), .ZN(n15090) );
  INV_X1 U8913 ( .A(n15090), .ZN(n15091) );
  BUF_X1 U8914 ( .A(n15094), .Z(n15092) );
  INV_X1 U8915 ( .A(n15096), .ZN(n15093) );
  INV_X1 U8916 ( .A(n15093), .ZN(n15094) );
  INV_X1 U8917 ( .A(n72420), .ZN(n15095) );
  INV_X1 U8918 ( .A(n15095), .ZN(n15096) );
  BUF_X1 U8919 ( .A(n15099), .Z(n15097) );
  INV_X1 U8920 ( .A(n15101), .ZN(n15098) );
  INV_X1 U8921 ( .A(n15098), .ZN(n15099) );
  INV_X1 U8922 ( .A(n72410), .ZN(n15100) );
  INV_X1 U8923 ( .A(n15100), .ZN(n15101) );
  BUF_X1 U8924 ( .A(n15104), .Z(n15102) );
  INV_X1 U8925 ( .A(n15106), .ZN(n15103) );
  INV_X1 U8926 ( .A(n15103), .ZN(n15104) );
  INV_X1 U8927 ( .A(n72400), .ZN(n15105) );
  INV_X1 U8928 ( .A(n15105), .ZN(n15106) );
  BUF_X1 U8929 ( .A(n15109), .Z(n15107) );
  INV_X1 U8930 ( .A(n15111), .ZN(n15108) );
  INV_X1 U8931 ( .A(n15108), .ZN(n15109) );
  INV_X1 U8932 ( .A(n72390), .ZN(n15110) );
  INV_X1 U8933 ( .A(n15110), .ZN(n15111) );
  BUF_X1 U8934 ( .A(n15114), .Z(n15112) );
  INV_X1 U8935 ( .A(n15116), .ZN(n15113) );
  INV_X1 U8936 ( .A(n15113), .ZN(n15114) );
  INV_X1 U8937 ( .A(n72380), .ZN(n15115) );
  INV_X1 U8938 ( .A(n15115), .ZN(n15116) );
  BUF_X1 U8939 ( .A(n15119), .Z(n15117) );
  INV_X1 U8940 ( .A(n15121), .ZN(n15118) );
  INV_X1 U8941 ( .A(n15118), .ZN(n15119) );
  INV_X1 U8942 ( .A(n72370), .ZN(n15120) );
  INV_X1 U8943 ( .A(n15120), .ZN(n15121) );
  BUF_X1 U8944 ( .A(n15124), .Z(n15122) );
  INV_X1 U8945 ( .A(n15126), .ZN(n15123) );
  INV_X1 U8946 ( .A(n15123), .ZN(n15124) );
  INV_X1 U8947 ( .A(n72360), .ZN(n15125) );
  INV_X1 U8948 ( .A(n15125), .ZN(n15126) );
  BUF_X1 U8949 ( .A(n15129), .Z(n15127) );
  INV_X1 U8950 ( .A(n15131), .ZN(n15128) );
  INV_X1 U8951 ( .A(n15128), .ZN(n15129) );
  INV_X1 U8952 ( .A(n72350), .ZN(n15130) );
  INV_X1 U8953 ( .A(n15130), .ZN(n15131) );
  BUF_X1 U8954 ( .A(n15134), .Z(n15132) );
  INV_X1 U8955 ( .A(n15136), .ZN(n15133) );
  INV_X1 U8956 ( .A(n15133), .ZN(n15134) );
  INV_X1 U8957 ( .A(n72340), .ZN(n15135) );
  INV_X1 U8958 ( .A(n15135), .ZN(n15136) );
  BUF_X1 U8959 ( .A(n15139), .Z(n15137) );
  INV_X1 U8960 ( .A(n15141), .ZN(n15138) );
  INV_X1 U8961 ( .A(n15138), .ZN(n15139) );
  INV_X1 U8962 ( .A(n72330), .ZN(n15140) );
  INV_X1 U8963 ( .A(n15140), .ZN(n15141) );
  BUF_X1 U8964 ( .A(n15144), .Z(n15142) );
  INV_X1 U8965 ( .A(n15146), .ZN(n15143) );
  INV_X1 U8966 ( .A(n15143), .ZN(n15144) );
  INV_X1 U8967 ( .A(n72320), .ZN(n15145) );
  INV_X1 U8968 ( .A(n15145), .ZN(n15146) );
  BUF_X1 U8969 ( .A(n15149), .Z(n15147) );
  INV_X1 U8970 ( .A(n15151), .ZN(n15148) );
  INV_X1 U8971 ( .A(n15148), .ZN(n15149) );
  INV_X1 U8972 ( .A(n72310), .ZN(n15150) );
  INV_X1 U8973 ( .A(n15150), .ZN(n15151) );
  BUF_X1 U8974 ( .A(n15154), .Z(n15152) );
  INV_X1 U8975 ( .A(n15156), .ZN(n15153) );
  INV_X1 U8976 ( .A(n15153), .ZN(n15154) );
  INV_X1 U8977 ( .A(n72300), .ZN(n15155) );
  INV_X1 U8978 ( .A(n15155), .ZN(n15156) );
  BUF_X1 U8979 ( .A(n15159), .Z(n15157) );
  INV_X1 U8980 ( .A(n15161), .ZN(n15158) );
  INV_X1 U8981 ( .A(n15158), .ZN(n15159) );
  INV_X1 U8982 ( .A(n72290), .ZN(n15160) );
  INV_X1 U8983 ( .A(n15160), .ZN(n15161) );
  BUF_X1 U8984 ( .A(n15164), .Z(n15162) );
  INV_X1 U8985 ( .A(n15166), .ZN(n15163) );
  INV_X1 U8986 ( .A(n15163), .ZN(n15164) );
  INV_X1 U8987 ( .A(n72280), .ZN(n15165) );
  INV_X1 U8988 ( .A(n15165), .ZN(n15166) );
  BUF_X1 U8989 ( .A(n15169), .Z(n15167) );
  INV_X1 U8990 ( .A(n15171), .ZN(n15168) );
  INV_X1 U8991 ( .A(n15168), .ZN(n15169) );
  INV_X1 U8992 ( .A(n72270), .ZN(n15170) );
  INV_X1 U8993 ( .A(n15170), .ZN(n15171) );
  BUF_X1 U8994 ( .A(n15174), .Z(n15172) );
  INV_X1 U8995 ( .A(n15176), .ZN(n15173) );
  INV_X1 U8996 ( .A(n15173), .ZN(n15174) );
  INV_X1 U8997 ( .A(n72260), .ZN(n15175) );
  INV_X1 U8998 ( .A(n15175), .ZN(n15176) );
  INV_X1 U8999 ( .A(n1228), .ZN(n15206) );
  BUF_X1 U9000 ( .A(n15207), .Z(n15177) );
  INV_X1 U9001 ( .A(n72250), .ZN(n15178) );
  INV_X1 U9002 ( .A(n15178), .ZN(n15179) );
  INV_X1 U9003 ( .A(n1227), .ZN(n15213) );
  BUF_X1 U9004 ( .A(n15214), .Z(n15180) );
  INV_X1 U9005 ( .A(n72240), .ZN(n15181) );
  INV_X1 U9006 ( .A(n15181), .ZN(n15182) );
  INV_X1 U9007 ( .A(n1226), .ZN(n15220) );
  BUF_X1 U9008 ( .A(n15221), .Z(n15183) );
  INV_X1 U9009 ( .A(n72230), .ZN(n15184) );
  INV_X1 U9010 ( .A(n15184), .ZN(n15185) );
  INV_X1 U9011 ( .A(n1225), .ZN(n15227) );
  BUF_X1 U9012 ( .A(n15228), .Z(n15186) );
  INV_X1 U9013 ( .A(n72220), .ZN(n15187) );
  INV_X1 U9014 ( .A(n15187), .ZN(n15188) );
  INV_X1 U9015 ( .A(n1224), .ZN(n15234) );
  BUF_X1 U9016 ( .A(n15235), .Z(n15189) );
  INV_X1 U9017 ( .A(n7221), .ZN(n15190) );
  INV_X1 U9018 ( .A(n15190), .ZN(n15191) );
  INV_X1 U9019 ( .A(n1223), .ZN(n15241) );
  BUF_X1 U9020 ( .A(n15242), .Z(n15192) );
  INV_X1 U9021 ( .A(n7220), .ZN(n15193) );
  INV_X1 U9022 ( .A(n15193), .ZN(n15194) );
  INV_X1 U9023 ( .A(n1222), .ZN(n15248) );
  BUF_X1 U9024 ( .A(n15249), .Z(n15195) );
  INV_X1 U9025 ( .A(n7219), .ZN(n15196) );
  INV_X1 U9026 ( .A(n15196), .ZN(n15197) );
  INV_X1 U9027 ( .A(n1221), .ZN(n15255) );
  BUF_X1 U9028 ( .A(n15256), .Z(n15198) );
  INV_X1 U9029 ( .A(n7218), .ZN(n15199) );
  INV_X1 U9030 ( .A(n15199), .ZN(n15200) );
  BUF_X1 U9031 ( .A(n15203), .Z(n15201) );
  INV_X1 U9032 ( .A(n15205), .ZN(n15202) );
  INV_X1 U9033 ( .A(n15202), .ZN(n15203) );
  INV_X1 U9034 ( .A(n7217), .ZN(n15204) );
  INV_X1 U9035 ( .A(n15204), .ZN(n15205) );
  INV_X1 U9036 ( .A(n15206), .ZN(n15207) );
  BUF_X1 U9037 ( .A(n15210), .Z(n15208) );
  INV_X1 U9038 ( .A(n15212), .ZN(n15209) );
  INV_X1 U9039 ( .A(n15209), .ZN(n15210) );
  INV_X1 U9040 ( .A(n7216), .ZN(n15211) );
  INV_X1 U9041 ( .A(n15211), .ZN(n15212) );
  INV_X1 U9042 ( .A(n15213), .ZN(n15214) );
  BUF_X1 U9043 ( .A(n15217), .Z(n15215) );
  INV_X1 U9044 ( .A(n15219), .ZN(n15216) );
  INV_X1 U9045 ( .A(n15216), .ZN(n15217) );
  INV_X1 U9046 ( .A(n7215), .ZN(n15218) );
  INV_X1 U9047 ( .A(n15218), .ZN(n15219) );
  INV_X1 U9048 ( .A(n15220), .ZN(n15221) );
  BUF_X1 U9049 ( .A(n15224), .Z(n15222) );
  INV_X1 U9050 ( .A(n15226), .ZN(n15223) );
  INV_X1 U9051 ( .A(n15223), .ZN(n15224) );
  INV_X1 U9052 ( .A(n7214), .ZN(n15225) );
  INV_X1 U9053 ( .A(n15225), .ZN(n15226) );
  INV_X1 U9054 ( .A(n15227), .ZN(n15228) );
  BUF_X1 U9055 ( .A(n15231), .Z(n15229) );
  INV_X1 U9056 ( .A(n15233), .ZN(n15230) );
  INV_X1 U9057 ( .A(n15230), .ZN(n15231) );
  INV_X1 U9058 ( .A(n7213), .ZN(n15232) );
  INV_X1 U9059 ( .A(n15232), .ZN(n15233) );
  INV_X1 U9060 ( .A(n15234), .ZN(n15235) );
  BUF_X1 U9061 ( .A(n15238), .Z(n15236) );
  INV_X1 U9062 ( .A(n15240), .ZN(n15237) );
  INV_X1 U9063 ( .A(n15237), .ZN(n15238) );
  INV_X1 U9064 ( .A(n7212), .ZN(n15239) );
  INV_X1 U9065 ( .A(n15239), .ZN(n15240) );
  INV_X1 U9066 ( .A(n15241), .ZN(n15242) );
  BUF_X1 U9067 ( .A(n15245), .Z(n15243) );
  INV_X1 U9068 ( .A(n15247), .ZN(n15244) );
  INV_X1 U9069 ( .A(n15244), .ZN(n15245) );
  INV_X1 U9070 ( .A(n7211), .ZN(n15246) );
  INV_X1 U9071 ( .A(n15246), .ZN(n15247) );
  INV_X1 U9072 ( .A(n15248), .ZN(n15249) );
  BUF_X1 U9073 ( .A(n15252), .Z(n15250) );
  INV_X1 U9074 ( .A(n15254), .ZN(n15251) );
  INV_X1 U9075 ( .A(n15251), .ZN(n15252) );
  INV_X1 U9076 ( .A(n7210), .ZN(n15253) );
  INV_X1 U9077 ( .A(n15253), .ZN(n15254) );
  INV_X1 U9078 ( .A(n15255), .ZN(n15256) );
  BUF_X1 U9079 ( .A(n15259), .Z(n15257) );
  INV_X1 U9080 ( .A(n15261), .ZN(n15258) );
  INV_X1 U9081 ( .A(n15258), .ZN(n15259) );
  INV_X1 U9082 ( .A(n7209), .ZN(n15260) );
  INV_X1 U9083 ( .A(n15260), .ZN(n15261) );
  BUF_X1 U9084 ( .A(n15264), .Z(n15262) );
  INV_X1 U9085 ( .A(n15266), .ZN(n15263) );
  INV_X1 U9086 ( .A(n15263), .ZN(n15264) );
  INV_X1 U9087 ( .A(n7208), .ZN(n15265) );
  INV_X1 U9088 ( .A(n15265), .ZN(n15266) );
  BUF_X1 U9089 ( .A(n15269), .Z(n15267) );
  INV_X1 U9090 ( .A(n15271), .ZN(n15268) );
  INV_X1 U9091 ( .A(n15268), .ZN(n15269) );
  INV_X1 U9092 ( .A(n7207), .ZN(n15270) );
  INV_X1 U9093 ( .A(n15270), .ZN(n15271) );
  BUF_X1 U9094 ( .A(n15274), .Z(n15272) );
  INV_X1 U9095 ( .A(n15276), .ZN(n15273) );
  INV_X1 U9096 ( .A(n15273), .ZN(n15274) );
  INV_X1 U9097 ( .A(n7206), .ZN(n15275) );
  INV_X1 U9098 ( .A(n15275), .ZN(n15276) );
  BUF_X1 U9099 ( .A(n15279), .Z(n15277) );
  INV_X1 U9100 ( .A(n15281), .ZN(n15278) );
  INV_X1 U9101 ( .A(n15278), .ZN(n15279) );
  INV_X1 U9102 ( .A(n7205), .ZN(n15280) );
  INV_X1 U9103 ( .A(n15280), .ZN(n15281) );
  BUF_X1 U9104 ( .A(n15284), .Z(n15282) );
  INV_X1 U9105 ( .A(n15286), .ZN(n15283) );
  INV_X1 U9106 ( .A(n15283), .ZN(n15284) );
  INV_X1 U9107 ( .A(n72040), .ZN(n15285) );
  INV_X1 U9108 ( .A(n15285), .ZN(n15286) );
  BUF_X1 U9109 ( .A(n15289), .Z(n15287) );
  INV_X1 U9110 ( .A(n15291), .ZN(n15288) );
  INV_X1 U9111 ( .A(n15288), .ZN(n15289) );
  INV_X1 U9112 ( .A(n72030), .ZN(n15290) );
  INV_X1 U9113 ( .A(n15290), .ZN(n15291) );
  BUF_X1 U9114 ( .A(n15294), .Z(n15292) );
  INV_X1 U9115 ( .A(n15296), .ZN(n15293) );
  INV_X1 U9116 ( .A(n15293), .ZN(n15294) );
  INV_X1 U9117 ( .A(n72020), .ZN(n15295) );
  INV_X1 U9118 ( .A(n15295), .ZN(n15296) );
  BUF_X1 U9119 ( .A(n15299), .Z(n15297) );
  INV_X1 U9120 ( .A(n15301), .ZN(n15298) );
  INV_X1 U9121 ( .A(n15298), .ZN(n15299) );
  INV_X1 U9122 ( .A(n72010), .ZN(n15300) );
  INV_X1 U9123 ( .A(n15300), .ZN(n15301) );
  BUF_X1 U9124 ( .A(n15304), .Z(n15302) );
  INV_X1 U9125 ( .A(n15306), .ZN(n15303) );
  INV_X1 U9126 ( .A(n15303), .ZN(n15304) );
  INV_X1 U9127 ( .A(n72000), .ZN(n15305) );
  INV_X1 U9128 ( .A(n15305), .ZN(n15306) );
  BUF_X1 U9129 ( .A(n15309), .Z(n15307) );
  INV_X1 U9130 ( .A(n15311), .ZN(n15308) );
  INV_X1 U9131 ( .A(n15308), .ZN(n15309) );
  INV_X1 U9132 ( .A(n71990), .ZN(n15310) );
  INV_X1 U9133 ( .A(n15310), .ZN(n15311) );
  BUF_X1 U9134 ( .A(n15314), .Z(n15312) );
  INV_X1 U9135 ( .A(n15316), .ZN(n15313) );
  INV_X1 U9136 ( .A(n15313), .ZN(n15314) );
  INV_X1 U9137 ( .A(n71980), .ZN(n15315) );
  INV_X1 U9138 ( .A(n15315), .ZN(n15316) );
  BUF_X1 U9139 ( .A(n15319), .Z(n15317) );
  INV_X1 U9140 ( .A(n15321), .ZN(n15318) );
  INV_X1 U9141 ( .A(n15318), .ZN(n15319) );
  INV_X1 U9142 ( .A(n71970), .ZN(n15320) );
  INV_X1 U9143 ( .A(n15320), .ZN(n15321) );
  BUF_X1 U9144 ( .A(n15324), .Z(n15322) );
  INV_X1 U9145 ( .A(n15326), .ZN(n15323) );
  INV_X1 U9146 ( .A(n15323), .ZN(n15324) );
  INV_X1 U9147 ( .A(n71960), .ZN(n15325) );
  INV_X1 U9148 ( .A(n15325), .ZN(n15326) );
  BUF_X1 U9149 ( .A(n15329), .Z(n15327) );
  INV_X1 U9150 ( .A(n15331), .ZN(n15328) );
  INV_X1 U9151 ( .A(n15328), .ZN(n15329) );
  INV_X1 U9152 ( .A(n71950), .ZN(n15330) );
  INV_X1 U9153 ( .A(n15330), .ZN(n15331) );
  BUF_X1 U9154 ( .A(n15334), .Z(n15332) );
  INV_X1 U9155 ( .A(n15336), .ZN(n15333) );
  INV_X1 U9156 ( .A(n15333), .ZN(n15334) );
  INV_X1 U9157 ( .A(n71940), .ZN(n15335) );
  INV_X1 U9158 ( .A(n15335), .ZN(n15336) );
  BUF_X1 U9159 ( .A(n15339), .Z(n15337) );
  INV_X1 U9160 ( .A(n15341), .ZN(n15338) );
  INV_X1 U9161 ( .A(n15338), .ZN(n15339) );
  INV_X1 U9162 ( .A(n71930), .ZN(n15340) );
  INV_X1 U9163 ( .A(n15340), .ZN(n15341) );
  BUF_X1 U9164 ( .A(n15344), .Z(n15342) );
  INV_X1 U9165 ( .A(n15346), .ZN(n15343) );
  INV_X1 U9166 ( .A(n15343), .ZN(n15344) );
  INV_X1 U9167 ( .A(n71920), .ZN(n15345) );
  INV_X1 U9168 ( .A(n15345), .ZN(n15346) );
  BUF_X1 U9169 ( .A(n15349), .Z(n15347) );
  INV_X1 U9170 ( .A(n15351), .ZN(n15348) );
  INV_X1 U9171 ( .A(n15348), .ZN(n15349) );
  INV_X1 U9172 ( .A(n71910), .ZN(n15350) );
  INV_X1 U9173 ( .A(n15350), .ZN(n15351) );
  BUF_X1 U9174 ( .A(n15354), .Z(n15352) );
  INV_X1 U9175 ( .A(n15356), .ZN(n15353) );
  INV_X1 U9176 ( .A(n15353), .ZN(n15354) );
  INV_X1 U9177 ( .A(n71900), .ZN(n15355) );
  INV_X1 U9178 ( .A(n15355), .ZN(n15356) );
  BUF_X1 U9179 ( .A(n15359), .Z(n15357) );
  INV_X1 U9180 ( .A(n15361), .ZN(n15358) );
  INV_X1 U9181 ( .A(n15358), .ZN(n15359) );
  INV_X1 U9182 ( .A(n71890), .ZN(n15360) );
  INV_X1 U9183 ( .A(n15360), .ZN(n15361) );
  BUF_X1 U9184 ( .A(n15364), .Z(n15362) );
  INV_X1 U9185 ( .A(n15366), .ZN(n15363) );
  INV_X1 U9186 ( .A(n15363), .ZN(n15364) );
  INV_X1 U9187 ( .A(n7188), .ZN(n15365) );
  INV_X1 U9188 ( .A(n15365), .ZN(n15366) );
  BUF_X1 U9189 ( .A(n15369), .Z(n15367) );
  INV_X1 U9190 ( .A(n15371), .ZN(n15368) );
  INV_X1 U9191 ( .A(n15368), .ZN(n15369) );
  INV_X1 U9192 ( .A(n7187), .ZN(n15370) );
  INV_X1 U9193 ( .A(n15370), .ZN(n15371) );
  BUF_X1 U9194 ( .A(n15374), .Z(n15372) );
  INV_X1 U9195 ( .A(n15376), .ZN(n15373) );
  INV_X1 U9196 ( .A(n15373), .ZN(n15374) );
  INV_X1 U9197 ( .A(n7186), .ZN(n15375) );
  INV_X1 U9198 ( .A(n15375), .ZN(n15376) );
  BUF_X1 U9199 ( .A(n15379), .Z(n15377) );
  INV_X1 U9200 ( .A(n15381), .ZN(n15378) );
  INV_X1 U9201 ( .A(n15378), .ZN(n15379) );
  INV_X1 U9202 ( .A(n7185), .ZN(n15380) );
  INV_X1 U9203 ( .A(n15380), .ZN(n15381) );
  BUF_X1 U9204 ( .A(n15384), .Z(n15382) );
  INV_X1 U9205 ( .A(n15386), .ZN(n15383) );
  INV_X1 U9206 ( .A(n15383), .ZN(n15384) );
  INV_X1 U9207 ( .A(n7184), .ZN(n15385) );
  INV_X1 U9208 ( .A(n15385), .ZN(n15386) );
  BUF_X1 U9209 ( .A(n15389), .Z(n15387) );
  INV_X1 U9210 ( .A(n15391), .ZN(n15388) );
  INV_X1 U9211 ( .A(n15388), .ZN(n15389) );
  INV_X1 U9212 ( .A(n7183), .ZN(n15390) );
  INV_X1 U9213 ( .A(n15390), .ZN(n15391) );
  BUF_X1 U9214 ( .A(n15394), .Z(n15392) );
  INV_X1 U9215 ( .A(n15396), .ZN(n15393) );
  INV_X1 U9216 ( .A(n15393), .ZN(n15394) );
  INV_X1 U9217 ( .A(n7182), .ZN(n15395) );
  INV_X1 U9218 ( .A(n15395), .ZN(n15396) );
  BUF_X1 U9219 ( .A(n15399), .Z(n15397) );
  INV_X1 U9220 ( .A(n15401), .ZN(n15398) );
  INV_X1 U9221 ( .A(n15398), .ZN(n15399) );
  INV_X1 U9222 ( .A(n7181), .ZN(n15400) );
  INV_X1 U9223 ( .A(n15400), .ZN(n15401) );
  BUF_X1 U9224 ( .A(n15404), .Z(n15402) );
  INV_X1 U9225 ( .A(n15406), .ZN(n15403) );
  INV_X1 U9226 ( .A(n15403), .ZN(n15404) );
  INV_X1 U9227 ( .A(n7180), .ZN(n15405) );
  INV_X1 U9228 ( .A(n15405), .ZN(n15406) );
  BUF_X1 U9229 ( .A(n15409), .Z(n15407) );
  INV_X1 U9230 ( .A(n15411), .ZN(n15408) );
  INV_X1 U9231 ( .A(n15408), .ZN(n15409) );
  INV_X1 U9232 ( .A(n7179), .ZN(n15410) );
  INV_X1 U9233 ( .A(n15410), .ZN(n15411) );
  BUF_X1 U9234 ( .A(n15414), .Z(n15412) );
  INV_X1 U9235 ( .A(n15416), .ZN(n15413) );
  INV_X1 U9236 ( .A(n15413), .ZN(n15414) );
  INV_X1 U9237 ( .A(n7178), .ZN(n15415) );
  INV_X1 U9238 ( .A(n15415), .ZN(n15416) );
  BUF_X1 U9239 ( .A(n15419), .Z(n15417) );
  INV_X1 U9240 ( .A(n15421), .ZN(n15418) );
  INV_X1 U9241 ( .A(n15418), .ZN(n15419) );
  INV_X1 U9242 ( .A(n7177), .ZN(n15420) );
  INV_X1 U9243 ( .A(n15420), .ZN(n15421) );
  BUF_X1 U9244 ( .A(n15424), .Z(n15422) );
  INV_X1 U9245 ( .A(n15426), .ZN(n15423) );
  INV_X1 U9246 ( .A(n15423), .ZN(n15424) );
  INV_X1 U9247 ( .A(n7176), .ZN(n15425) );
  INV_X1 U9248 ( .A(n15425), .ZN(n15426) );
  BUF_X1 U9249 ( .A(n15429), .Z(n15427) );
  INV_X1 U9250 ( .A(n15431), .ZN(n15428) );
  INV_X1 U9251 ( .A(n15428), .ZN(n15429) );
  INV_X1 U9252 ( .A(n7175), .ZN(n15430) );
  INV_X1 U9253 ( .A(n15430), .ZN(n15431) );
  BUF_X1 U9254 ( .A(n15434), .Z(n15432) );
  INV_X1 U9255 ( .A(n15436), .ZN(n15433) );
  INV_X1 U9256 ( .A(n15433), .ZN(n15434) );
  INV_X1 U9257 ( .A(n7174), .ZN(n15435) );
  INV_X1 U9258 ( .A(n15435), .ZN(n15436) );
  BUF_X1 U9259 ( .A(n15439), .Z(n15437) );
  INV_X1 U9260 ( .A(n15441), .ZN(n15438) );
  INV_X1 U9261 ( .A(n15438), .ZN(n15439) );
  INV_X1 U9262 ( .A(n7173), .ZN(n15440) );
  INV_X1 U9263 ( .A(n15440), .ZN(n15441) );
  BUF_X1 U9264 ( .A(n15444), .Z(n15442) );
  INV_X1 U9265 ( .A(n15446), .ZN(n15443) );
  INV_X1 U9266 ( .A(n15443), .ZN(n15444) );
  INV_X1 U9267 ( .A(n7172), .ZN(n15445) );
  INV_X1 U9268 ( .A(n15445), .ZN(n15446) );
  BUF_X1 U9269 ( .A(n15449), .Z(n15447) );
  INV_X1 U9270 ( .A(n15451), .ZN(n15448) );
  INV_X1 U9271 ( .A(n15448), .ZN(n15449) );
  INV_X1 U9272 ( .A(n7171), .ZN(n15450) );
  INV_X1 U9273 ( .A(n15450), .ZN(n15451) );
  BUF_X1 U9274 ( .A(n15454), .Z(n15452) );
  INV_X1 U9275 ( .A(n15456), .ZN(n15453) );
  INV_X1 U9276 ( .A(n15453), .ZN(n15454) );
  INV_X1 U9277 ( .A(n7170), .ZN(n15455) );
  INV_X1 U9278 ( .A(n15455), .ZN(n15456) );
  BUF_X1 U9279 ( .A(n15459), .Z(n15457) );
  INV_X1 U9280 ( .A(n15461), .ZN(n15458) );
  INV_X1 U9281 ( .A(n15458), .ZN(n15459) );
  INV_X1 U9282 ( .A(n7169), .ZN(n15460) );
  INV_X1 U9283 ( .A(n15460), .ZN(n15461) );
  BUF_X1 U9284 ( .A(n15464), .Z(n15462) );
  INV_X1 U9285 ( .A(n15466), .ZN(n15463) );
  INV_X1 U9286 ( .A(n15463), .ZN(n15464) );
  INV_X1 U9287 ( .A(n7168), .ZN(n15465) );
  INV_X1 U9288 ( .A(n15465), .ZN(n15466) );
  BUF_X1 U9289 ( .A(n15469), .Z(n15467) );
  INV_X1 U9290 ( .A(n15471), .ZN(n15468) );
  INV_X1 U9291 ( .A(n15468), .ZN(n15469) );
  INV_X1 U9292 ( .A(n7167), .ZN(n15470) );
  INV_X1 U9293 ( .A(n15470), .ZN(n15471) );
  BUF_X1 U9294 ( .A(n15474), .Z(n15472) );
  INV_X1 U9295 ( .A(n15476), .ZN(n15473) );
  INV_X1 U9296 ( .A(n15473), .ZN(n15474) );
  INV_X1 U9297 ( .A(n7166), .ZN(n15475) );
  INV_X1 U9298 ( .A(n15475), .ZN(n15476) );
  BUF_X1 U9299 ( .A(n15479), .Z(n15477) );
  INV_X1 U9300 ( .A(n15481), .ZN(n15478) );
  INV_X1 U9301 ( .A(n15478), .ZN(n15479) );
  INV_X1 U9302 ( .A(n7165), .ZN(n15480) );
  INV_X1 U9303 ( .A(n15480), .ZN(n15481) );
  BUF_X1 U9304 ( .A(n15484), .Z(n15482) );
  INV_X1 U9305 ( .A(n15486), .ZN(n15483) );
  INV_X1 U9306 ( .A(n15483), .ZN(n15484) );
  INV_X1 U9307 ( .A(n7164), .ZN(n15485) );
  INV_X1 U9308 ( .A(n15485), .ZN(n15486) );
  BUF_X1 U9309 ( .A(n15489), .Z(n15487) );
  INV_X1 U9310 ( .A(n15491), .ZN(n15488) );
  INV_X1 U9311 ( .A(n15488), .ZN(n15489) );
  INV_X1 U9312 ( .A(n7163), .ZN(n15490) );
  INV_X1 U9313 ( .A(n15490), .ZN(n15491) );
  BUF_X1 U9314 ( .A(n15494), .Z(n15492) );
  INV_X1 U9315 ( .A(n15496), .ZN(n15493) );
  INV_X1 U9316 ( .A(n15493), .ZN(n15494) );
  INV_X1 U9317 ( .A(n7162), .ZN(n15495) );
  INV_X1 U9318 ( .A(n15495), .ZN(n15496) );
  INV_X1 U9319 ( .A(n1172), .ZN(n15526) );
  BUF_X1 U9320 ( .A(n15527), .Z(n15497) );
  INV_X1 U9321 ( .A(n7161), .ZN(n15498) );
  INV_X1 U9322 ( .A(n15498), .ZN(n15499) );
  INV_X1 U9323 ( .A(n1171), .ZN(n15533) );
  BUF_X1 U9324 ( .A(n15534), .Z(n15500) );
  INV_X1 U9325 ( .A(n7160), .ZN(n15501) );
  INV_X1 U9326 ( .A(n15501), .ZN(n15502) );
  INV_X1 U9327 ( .A(n1170), .ZN(n15540) );
  BUF_X1 U9328 ( .A(n15541), .Z(n15503) );
  INV_X1 U9329 ( .A(n7159), .ZN(n15504) );
  INV_X1 U9330 ( .A(n15504), .ZN(n15505) );
  INV_X1 U9331 ( .A(n1169), .ZN(n15547) );
  BUF_X1 U9332 ( .A(n15548), .Z(n15506) );
  INV_X1 U9333 ( .A(n7158), .ZN(n15507) );
  INV_X1 U9334 ( .A(n15507), .ZN(n15508) );
  INV_X1 U9335 ( .A(n1168), .ZN(n15554) );
  BUF_X1 U9336 ( .A(n15555), .Z(n15509) );
  INV_X1 U9337 ( .A(n7157), .ZN(n15510) );
  INV_X1 U9338 ( .A(n15510), .ZN(n15511) );
  INV_X1 U9339 ( .A(n1167), .ZN(n15561) );
  BUF_X1 U9340 ( .A(n15562), .Z(n15512) );
  INV_X1 U9341 ( .A(n7156), .ZN(n15513) );
  INV_X1 U9342 ( .A(n15513), .ZN(n15514) );
  INV_X1 U9343 ( .A(n1166), .ZN(n15568) );
  BUF_X1 U9344 ( .A(n15569), .Z(n15515) );
  INV_X1 U9345 ( .A(n7155), .ZN(n15516) );
  INV_X1 U9346 ( .A(n15516), .ZN(n15517) );
  INV_X1 U9347 ( .A(n1165), .ZN(n15575) );
  BUF_X1 U9348 ( .A(n15576), .Z(n15518) );
  INV_X1 U9349 ( .A(n7154), .ZN(n15519) );
  INV_X1 U9350 ( .A(n15519), .ZN(n15520) );
  BUF_X1 U9351 ( .A(n15523), .Z(n15521) );
  INV_X1 U9352 ( .A(n15525), .ZN(n15522) );
  INV_X1 U9353 ( .A(n15522), .ZN(n15523) );
  INV_X1 U9354 ( .A(n7153), .ZN(n15524) );
  INV_X1 U9355 ( .A(n15524), .ZN(n15525) );
  INV_X1 U9356 ( .A(n15526), .ZN(n15527) );
  BUF_X1 U9357 ( .A(n15530), .Z(n15528) );
  INV_X1 U9358 ( .A(n15532), .ZN(n15529) );
  INV_X1 U9359 ( .A(n15529), .ZN(n15530) );
  INV_X1 U9360 ( .A(n7152), .ZN(n15531) );
  INV_X1 U9361 ( .A(n15531), .ZN(n15532) );
  INV_X1 U9362 ( .A(n15533), .ZN(n15534) );
  BUF_X1 U9363 ( .A(n15537), .Z(n15535) );
  INV_X1 U9364 ( .A(n15539), .ZN(n15536) );
  INV_X1 U9365 ( .A(n15536), .ZN(n15537) );
  INV_X1 U9366 ( .A(n7151), .ZN(n15538) );
  INV_X1 U9367 ( .A(n15538), .ZN(n15539) );
  INV_X1 U9368 ( .A(n15540), .ZN(n15541) );
  BUF_X1 U9369 ( .A(n15544), .Z(n15542) );
  INV_X1 U9370 ( .A(n15546), .ZN(n15543) );
  INV_X1 U9371 ( .A(n15543), .ZN(n15544) );
  INV_X1 U9372 ( .A(n71500), .ZN(n15545) );
  INV_X1 U9373 ( .A(n15545), .ZN(n15546) );
  INV_X1 U9374 ( .A(n15547), .ZN(n15548) );
  BUF_X1 U9375 ( .A(n15551), .Z(n15549) );
  INV_X1 U9376 ( .A(n15553), .ZN(n15550) );
  INV_X1 U9377 ( .A(n15550), .ZN(n15551) );
  INV_X1 U9378 ( .A(n71490), .ZN(n15552) );
  INV_X1 U9379 ( .A(n15552), .ZN(n15553) );
  INV_X1 U9380 ( .A(n15554), .ZN(n15555) );
  BUF_X1 U9381 ( .A(n15558), .Z(n15556) );
  INV_X1 U9382 ( .A(n15560), .ZN(n15557) );
  INV_X1 U9383 ( .A(n15557), .ZN(n15558) );
  INV_X1 U9384 ( .A(n71480), .ZN(n15559) );
  INV_X1 U9385 ( .A(n15559), .ZN(n15560) );
  INV_X1 U9386 ( .A(n15561), .ZN(n15562) );
  BUF_X1 U9387 ( .A(n15565), .Z(n15563) );
  INV_X1 U9388 ( .A(n15567), .ZN(n15564) );
  INV_X1 U9389 ( .A(n15564), .ZN(n15565) );
  INV_X1 U9390 ( .A(n71470), .ZN(n15566) );
  INV_X1 U9391 ( .A(n15566), .ZN(n15567) );
  INV_X1 U9392 ( .A(n15568), .ZN(n15569) );
  BUF_X1 U9393 ( .A(n15572), .Z(n15570) );
  INV_X1 U9394 ( .A(n15574), .ZN(n15571) );
  INV_X1 U9395 ( .A(n15571), .ZN(n15572) );
  INV_X1 U9396 ( .A(n71460), .ZN(n15573) );
  INV_X1 U9397 ( .A(n15573), .ZN(n15574) );
  INV_X1 U9398 ( .A(n15575), .ZN(n15576) );
  BUF_X1 U9399 ( .A(n15579), .Z(n15577) );
  INV_X1 U9400 ( .A(n15581), .ZN(n15578) );
  INV_X1 U9401 ( .A(n15578), .ZN(n15579) );
  INV_X1 U9402 ( .A(n71450), .ZN(n15580) );
  INV_X1 U9403 ( .A(n15580), .ZN(n15581) );
  BUF_X1 U9404 ( .A(n15584), .Z(n15582) );
  INV_X1 U9405 ( .A(n15586), .ZN(n15583) );
  INV_X1 U9406 ( .A(n15583), .ZN(n15584) );
  INV_X1 U9407 ( .A(n71440), .ZN(n15585) );
  INV_X1 U9408 ( .A(n15585), .ZN(n15586) );
  BUF_X1 U9409 ( .A(n15589), .Z(n15587) );
  INV_X1 U9410 ( .A(n15591), .ZN(n15588) );
  INV_X1 U9411 ( .A(n15588), .ZN(n15589) );
  INV_X1 U9412 ( .A(n71430), .ZN(n15590) );
  INV_X1 U9413 ( .A(n15590), .ZN(n15591) );
  BUF_X1 U9414 ( .A(n15594), .Z(n15592) );
  INV_X1 U9415 ( .A(n15596), .ZN(n15593) );
  INV_X1 U9416 ( .A(n15593), .ZN(n15594) );
  INV_X1 U9417 ( .A(n71420), .ZN(n15595) );
  INV_X1 U9418 ( .A(n15595), .ZN(n15596) );
  BUF_X1 U9419 ( .A(n15599), .Z(n15597) );
  INV_X1 U9420 ( .A(n15601), .ZN(n15598) );
  INV_X1 U9421 ( .A(n15598), .ZN(n15599) );
  INV_X1 U9422 ( .A(n71410), .ZN(n15600) );
  INV_X1 U9423 ( .A(n15600), .ZN(n15601) );
  BUF_X1 U9424 ( .A(n15604), .Z(n15602) );
  INV_X1 U9425 ( .A(n15606), .ZN(n15603) );
  INV_X1 U9426 ( .A(n15603), .ZN(n15604) );
  INV_X1 U9427 ( .A(n71400), .ZN(n15605) );
  INV_X1 U9428 ( .A(n15605), .ZN(n15606) );
  BUF_X1 U9429 ( .A(n15609), .Z(n15607) );
  INV_X1 U9430 ( .A(n15611), .ZN(n15608) );
  INV_X1 U9431 ( .A(n15608), .ZN(n15609) );
  INV_X1 U9432 ( .A(n71390), .ZN(n15610) );
  INV_X1 U9433 ( .A(n15610), .ZN(n15611) );
  BUF_X1 U9434 ( .A(n15614), .Z(n15612) );
  INV_X1 U9435 ( .A(n15616), .ZN(n15613) );
  INV_X1 U9436 ( .A(n15613), .ZN(n15614) );
  INV_X1 U9437 ( .A(n71380), .ZN(n15615) );
  INV_X1 U9438 ( .A(n15615), .ZN(n15616) );
  BUF_X1 U9439 ( .A(n15619), .Z(n15617) );
  INV_X1 U9440 ( .A(n15621), .ZN(n15618) );
  INV_X1 U9441 ( .A(n15618), .ZN(n15619) );
  INV_X1 U9442 ( .A(n71370), .ZN(n15620) );
  INV_X1 U9443 ( .A(n15620), .ZN(n15621) );
  BUF_X1 U9444 ( .A(n15624), .Z(n15622) );
  INV_X1 U9445 ( .A(n15626), .ZN(n15623) );
  INV_X1 U9446 ( .A(n15623), .ZN(n15624) );
  INV_X1 U9447 ( .A(n71360), .ZN(n15625) );
  INV_X1 U9448 ( .A(n15625), .ZN(n15626) );
  BUF_X1 U9449 ( .A(n15629), .Z(n15627) );
  INV_X1 U9450 ( .A(n15631), .ZN(n15628) );
  INV_X1 U9451 ( .A(n15628), .ZN(n15629) );
  INV_X1 U9452 ( .A(n71350), .ZN(n15630) );
  INV_X1 U9453 ( .A(n15630), .ZN(n15631) );
  BUF_X1 U9454 ( .A(n15634), .Z(n15632) );
  INV_X1 U9455 ( .A(n15636), .ZN(n15633) );
  INV_X1 U9456 ( .A(n15633), .ZN(n15634) );
  INV_X1 U9457 ( .A(n71340), .ZN(n15635) );
  INV_X1 U9458 ( .A(n15635), .ZN(n15636) );
  BUF_X1 U9459 ( .A(n15639), .Z(n15637) );
  INV_X1 U9460 ( .A(n15641), .ZN(n15638) );
  INV_X1 U9461 ( .A(n15638), .ZN(n15639) );
  INV_X1 U9462 ( .A(n71330), .ZN(n15640) );
  INV_X1 U9463 ( .A(n15640), .ZN(n15641) );
  BUF_X1 U9464 ( .A(n15644), .Z(n15642) );
  INV_X1 U9465 ( .A(n15646), .ZN(n15643) );
  INV_X1 U9466 ( .A(n15643), .ZN(n15644) );
  INV_X1 U9467 ( .A(n71320), .ZN(n15645) );
  INV_X1 U9468 ( .A(n15645), .ZN(n15646) );
  BUF_X1 U9469 ( .A(n15649), .Z(n15647) );
  INV_X1 U9470 ( .A(n15651), .ZN(n15648) );
  INV_X1 U9471 ( .A(n15648), .ZN(n15649) );
  INV_X1 U9472 ( .A(n71310), .ZN(n15650) );
  INV_X1 U9473 ( .A(n15650), .ZN(n15651) );
  BUF_X1 U9474 ( .A(n15654), .Z(n15652) );
  INV_X1 U9475 ( .A(n15656), .ZN(n15653) );
  INV_X1 U9476 ( .A(n15653), .ZN(n15654) );
  INV_X1 U9477 ( .A(n71300), .ZN(n15655) );
  INV_X1 U9478 ( .A(n15655), .ZN(n15656) );
  BUF_X1 U9479 ( .A(n15659), .Z(n15657) );
  INV_X1 U9480 ( .A(n15661), .ZN(n15658) );
  INV_X1 U9481 ( .A(n15658), .ZN(n15659) );
  INV_X1 U9482 ( .A(n7129), .ZN(n15660) );
  INV_X1 U9483 ( .A(n15660), .ZN(n15661) );
  BUF_X1 U9484 ( .A(n15664), .Z(n15662) );
  INV_X1 U9485 ( .A(n15666), .ZN(n15663) );
  INV_X1 U9486 ( .A(n15663), .ZN(n15664) );
  INV_X1 U9487 ( .A(n7128), .ZN(n15665) );
  INV_X1 U9488 ( .A(n15665), .ZN(n15666) );
  BUF_X1 U9489 ( .A(n15669), .Z(n15667) );
  INV_X1 U9490 ( .A(n15671), .ZN(n15668) );
  INV_X1 U9491 ( .A(n15668), .ZN(n15669) );
  INV_X1 U9492 ( .A(n7127), .ZN(n15670) );
  INV_X1 U9493 ( .A(n15670), .ZN(n15671) );
  BUF_X1 U9494 ( .A(n15674), .Z(n15672) );
  INV_X1 U9495 ( .A(n15676), .ZN(n15673) );
  INV_X1 U9496 ( .A(n15673), .ZN(n15674) );
  INV_X1 U9497 ( .A(n7126), .ZN(n15675) );
  INV_X1 U9498 ( .A(n15675), .ZN(n15676) );
  BUF_X1 U9499 ( .A(n15679), .Z(n15677) );
  INV_X1 U9500 ( .A(n15681), .ZN(n15678) );
  INV_X1 U9501 ( .A(n15678), .ZN(n15679) );
  INV_X1 U9502 ( .A(n7125), .ZN(n15680) );
  INV_X1 U9503 ( .A(n15680), .ZN(n15681) );
  BUF_X1 U9504 ( .A(n15684), .Z(n15682) );
  INV_X1 U9505 ( .A(n15686), .ZN(n15683) );
  INV_X1 U9506 ( .A(n15683), .ZN(n15684) );
  INV_X1 U9507 ( .A(n7124), .ZN(n15685) );
  INV_X1 U9508 ( .A(n15685), .ZN(n15686) );
  BUF_X1 U9509 ( .A(n15689), .Z(n15687) );
  INV_X1 U9510 ( .A(n15691), .ZN(n15688) );
  INV_X1 U9511 ( .A(n15688), .ZN(n15689) );
  INV_X1 U9512 ( .A(n7123), .ZN(n15690) );
  INV_X1 U9513 ( .A(n15690), .ZN(n15691) );
  BUF_X1 U9514 ( .A(n15694), .Z(n15692) );
  INV_X1 U9515 ( .A(n15696), .ZN(n15693) );
  INV_X1 U9516 ( .A(n15693), .ZN(n15694) );
  INV_X1 U9517 ( .A(n7122), .ZN(n15695) );
  INV_X1 U9518 ( .A(n15695), .ZN(n15696) );
  BUF_X1 U9519 ( .A(n15699), .Z(n15697) );
  INV_X1 U9520 ( .A(n15701), .ZN(n15698) );
  INV_X1 U9521 ( .A(n15698), .ZN(n15699) );
  INV_X1 U9522 ( .A(n7121), .ZN(n15700) );
  INV_X1 U9523 ( .A(n15700), .ZN(n15701) );
  BUF_X1 U9524 ( .A(n15704), .Z(n15702) );
  INV_X1 U9525 ( .A(n15706), .ZN(n15703) );
  INV_X1 U9526 ( .A(n15703), .ZN(n15704) );
  INV_X1 U9527 ( .A(n7120), .ZN(n15705) );
  INV_X1 U9528 ( .A(n15705), .ZN(n15706) );
  BUF_X1 U9529 ( .A(n15709), .Z(n15707) );
  INV_X1 U9530 ( .A(n15711), .ZN(n15708) );
  INV_X1 U9531 ( .A(n15708), .ZN(n15709) );
  INV_X1 U9532 ( .A(n7119), .ZN(n15710) );
  INV_X1 U9533 ( .A(n15710), .ZN(n15711) );
  BUF_X1 U9534 ( .A(n15714), .Z(n15712) );
  INV_X1 U9535 ( .A(n15716), .ZN(n15713) );
  INV_X1 U9536 ( .A(n15713), .ZN(n15714) );
  INV_X1 U9537 ( .A(n7118), .ZN(n15715) );
  INV_X1 U9538 ( .A(n15715), .ZN(n15716) );
  BUF_X1 U9539 ( .A(n15719), .Z(n15717) );
  INV_X1 U9540 ( .A(n15721), .ZN(n15718) );
  INV_X1 U9541 ( .A(n15718), .ZN(n15719) );
  INV_X1 U9542 ( .A(n7117), .ZN(n15720) );
  INV_X1 U9543 ( .A(n15720), .ZN(n15721) );
  BUF_X1 U9544 ( .A(n15724), .Z(n15722) );
  INV_X1 U9545 ( .A(n15726), .ZN(n15723) );
  INV_X1 U9546 ( .A(n15723), .ZN(n15724) );
  INV_X1 U9547 ( .A(n7116), .ZN(n15725) );
  INV_X1 U9548 ( .A(n15725), .ZN(n15726) );
  BUF_X1 U9549 ( .A(n15729), .Z(n15727) );
  INV_X1 U9550 ( .A(n15731), .ZN(n15728) );
  INV_X1 U9551 ( .A(n15728), .ZN(n15729) );
  INV_X1 U9552 ( .A(n7115), .ZN(n15730) );
  INV_X1 U9553 ( .A(n15730), .ZN(n15731) );
  BUF_X1 U9554 ( .A(n15734), .Z(n15732) );
  INV_X1 U9555 ( .A(n15736), .ZN(n15733) );
  INV_X1 U9556 ( .A(n15733), .ZN(n15734) );
  INV_X1 U9557 ( .A(n7114), .ZN(n15735) );
  INV_X1 U9558 ( .A(n15735), .ZN(n15736) );
  BUF_X1 U9559 ( .A(n15739), .Z(n15737) );
  INV_X1 U9560 ( .A(n15741), .ZN(n15738) );
  INV_X1 U9561 ( .A(n15738), .ZN(n15739) );
  INV_X1 U9562 ( .A(n7113), .ZN(n15740) );
  INV_X1 U9563 ( .A(n15740), .ZN(n15741) );
  BUF_X1 U9564 ( .A(n15744), .Z(n15742) );
  INV_X1 U9565 ( .A(n15746), .ZN(n15743) );
  INV_X1 U9566 ( .A(n15743), .ZN(n15744) );
  INV_X1 U9567 ( .A(n71120), .ZN(n15745) );
  INV_X1 U9568 ( .A(n15745), .ZN(n15746) );
  BUF_X1 U9569 ( .A(n15749), .Z(n15747) );
  INV_X1 U9570 ( .A(n15751), .ZN(n15748) );
  INV_X1 U9571 ( .A(n15748), .ZN(n15749) );
  INV_X1 U9572 ( .A(n71110), .ZN(n15750) );
  INV_X1 U9573 ( .A(n15750), .ZN(n15751) );
  BUF_X1 U9574 ( .A(n15754), .Z(n15752) );
  INV_X1 U9575 ( .A(n15756), .ZN(n15753) );
  INV_X1 U9576 ( .A(n15753), .ZN(n15754) );
  INV_X1 U9577 ( .A(n71100), .ZN(n15755) );
  INV_X1 U9578 ( .A(n15755), .ZN(n15756) );
  BUF_X1 U9579 ( .A(n15759), .Z(n15757) );
  INV_X1 U9580 ( .A(n15761), .ZN(n15758) );
  INV_X1 U9581 ( .A(n15758), .ZN(n15759) );
  INV_X1 U9582 ( .A(n71090), .ZN(n15760) );
  INV_X1 U9583 ( .A(n15760), .ZN(n15761) );
  BUF_X1 U9584 ( .A(n15764), .Z(n15762) );
  INV_X1 U9585 ( .A(n15766), .ZN(n15763) );
  INV_X1 U9586 ( .A(n15763), .ZN(n15764) );
  INV_X1 U9587 ( .A(n71080), .ZN(n15765) );
  INV_X1 U9588 ( .A(n15765), .ZN(n15766) );
  BUF_X1 U9589 ( .A(n15769), .Z(n15767) );
  INV_X1 U9590 ( .A(n15771), .ZN(n15768) );
  INV_X1 U9591 ( .A(n15768), .ZN(n15769) );
  INV_X1 U9592 ( .A(n71070), .ZN(n15770) );
  INV_X1 U9593 ( .A(n15770), .ZN(n15771) );
  BUF_X1 U9594 ( .A(n15774), .Z(n15772) );
  INV_X1 U9595 ( .A(n15776), .ZN(n15773) );
  INV_X1 U9596 ( .A(n15773), .ZN(n15774) );
  INV_X1 U9597 ( .A(n71060), .ZN(n15775) );
  INV_X1 U9598 ( .A(n15775), .ZN(n15776) );
  BUF_X1 U9599 ( .A(n15779), .Z(n15777) );
  INV_X1 U9600 ( .A(n15781), .ZN(n15778) );
  INV_X1 U9601 ( .A(n15778), .ZN(n15779) );
  INV_X1 U9602 ( .A(n71050), .ZN(n15780) );
  INV_X1 U9603 ( .A(n15780), .ZN(n15781) );
  BUF_X1 U9604 ( .A(n15784), .Z(n15782) );
  INV_X1 U9605 ( .A(n15786), .ZN(n15783) );
  INV_X1 U9606 ( .A(n15783), .ZN(n15784) );
  INV_X1 U9607 ( .A(n71040), .ZN(n15785) );
  INV_X1 U9608 ( .A(n15785), .ZN(n15786) );
  BUF_X1 U9609 ( .A(n15789), .Z(n15787) );
  INV_X1 U9610 ( .A(n15791), .ZN(n15788) );
  INV_X1 U9611 ( .A(n15788), .ZN(n15789) );
  INV_X1 U9612 ( .A(n71030), .ZN(n15790) );
  INV_X1 U9613 ( .A(n15790), .ZN(n15791) );
  BUF_X1 U9614 ( .A(n15794), .Z(n15792) );
  INV_X1 U9615 ( .A(n15796), .ZN(n15793) );
  INV_X1 U9616 ( .A(n15793), .ZN(n15794) );
  INV_X1 U9617 ( .A(n71020), .ZN(n15795) );
  INV_X1 U9618 ( .A(n15795), .ZN(n15796) );
  BUF_X1 U9619 ( .A(n15799), .Z(n15797) );
  INV_X1 U9620 ( .A(n15801), .ZN(n15798) );
  INV_X1 U9621 ( .A(n15798), .ZN(n15799) );
  INV_X1 U9622 ( .A(n71010), .ZN(n15800) );
  INV_X1 U9623 ( .A(n15800), .ZN(n15801) );
  BUF_X1 U9624 ( .A(n15804), .Z(n15802) );
  INV_X1 U9625 ( .A(n15806), .ZN(n15803) );
  INV_X1 U9626 ( .A(n15803), .ZN(n15804) );
  INV_X1 U9627 ( .A(n71000), .ZN(n15805) );
  INV_X1 U9628 ( .A(n15805), .ZN(n15806) );
  BUF_X1 U9629 ( .A(n15809), .Z(n15807) );
  INV_X1 U9630 ( .A(n15811), .ZN(n15808) );
  INV_X1 U9631 ( .A(n15808), .ZN(n15809) );
  INV_X1 U9632 ( .A(n70990), .ZN(n15810) );
  INV_X1 U9633 ( .A(n15810), .ZN(n15811) );
  BUF_X1 U9634 ( .A(n15814), .Z(n15812) );
  INV_X1 U9635 ( .A(n15816), .ZN(n15813) );
  INV_X1 U9636 ( .A(n15813), .ZN(n15814) );
  INV_X1 U9637 ( .A(n70980), .ZN(n15815) );
  INV_X1 U9638 ( .A(n15815), .ZN(n15816) );
  INV_X1 U9639 ( .A(n1116), .ZN(n15846) );
  BUF_X1 U9640 ( .A(n15847), .Z(n15817) );
  INV_X1 U9641 ( .A(n70970), .ZN(n15818) );
  INV_X1 U9642 ( .A(n15818), .ZN(n15819) );
  INV_X1 U9643 ( .A(n1115), .ZN(n15853) );
  BUF_X1 U9644 ( .A(n15854), .Z(n15820) );
  INV_X1 U9645 ( .A(n7096), .ZN(n15821) );
  INV_X1 U9646 ( .A(n15821), .ZN(n15822) );
  INV_X1 U9647 ( .A(n1114), .ZN(n15860) );
  BUF_X1 U9648 ( .A(n15861), .Z(n15823) );
  INV_X1 U9649 ( .A(n7095), .ZN(n15824) );
  INV_X1 U9650 ( .A(n15824), .ZN(n15825) );
  INV_X1 U9651 ( .A(n1113), .ZN(n15867) );
  BUF_X1 U9652 ( .A(n15868), .Z(n15826) );
  INV_X1 U9653 ( .A(n7094), .ZN(n15827) );
  INV_X1 U9654 ( .A(n15827), .ZN(n15828) );
  INV_X1 U9655 ( .A(n1112), .ZN(n15874) );
  BUF_X1 U9656 ( .A(n15875), .Z(n15829) );
  INV_X1 U9657 ( .A(n7093), .ZN(n15830) );
  INV_X1 U9658 ( .A(n15830), .ZN(n15831) );
  INV_X1 U9659 ( .A(n1111), .ZN(n15881) );
  BUF_X1 U9660 ( .A(n15882), .Z(n15832) );
  INV_X1 U9661 ( .A(n7092), .ZN(n15833) );
  INV_X1 U9662 ( .A(n15833), .ZN(n15834) );
  INV_X1 U9663 ( .A(n1110), .ZN(n15888) );
  BUF_X1 U9664 ( .A(n15889), .Z(n15835) );
  INV_X1 U9665 ( .A(n7091), .ZN(n15836) );
  INV_X1 U9666 ( .A(n15836), .ZN(n15837) );
  INV_X1 U9667 ( .A(n1109), .ZN(n15895) );
  BUF_X1 U9668 ( .A(n15896), .Z(n15838) );
  INV_X1 U9669 ( .A(n7090), .ZN(n15839) );
  INV_X1 U9670 ( .A(n15839), .ZN(n15840) );
  BUF_X1 U9671 ( .A(n15843), .Z(n15841) );
  INV_X1 U9672 ( .A(n15845), .ZN(n15842) );
  INV_X1 U9673 ( .A(n15842), .ZN(n15843) );
  INV_X1 U9674 ( .A(n7089), .ZN(n15844) );
  INV_X1 U9675 ( .A(n15844), .ZN(n15845) );
  INV_X1 U9676 ( .A(n15846), .ZN(n15847) );
  BUF_X1 U9677 ( .A(n15850), .Z(n15848) );
  INV_X1 U9678 ( .A(n15852), .ZN(n15849) );
  INV_X1 U9679 ( .A(n15849), .ZN(n15850) );
  INV_X1 U9680 ( .A(n7088), .ZN(n15851) );
  INV_X1 U9681 ( .A(n15851), .ZN(n15852) );
  INV_X1 U9682 ( .A(n15853), .ZN(n15854) );
  BUF_X1 U9683 ( .A(n15857), .Z(n15855) );
  INV_X1 U9684 ( .A(n15859), .ZN(n15856) );
  INV_X1 U9685 ( .A(n15856), .ZN(n15857) );
  INV_X1 U9686 ( .A(n7087), .ZN(n15858) );
  INV_X1 U9687 ( .A(n15858), .ZN(n15859) );
  INV_X1 U9688 ( .A(n15860), .ZN(n15861) );
  BUF_X1 U9689 ( .A(n15864), .Z(n15862) );
  INV_X1 U9690 ( .A(n15866), .ZN(n15863) );
  INV_X1 U9691 ( .A(n15863), .ZN(n15864) );
  INV_X1 U9692 ( .A(n7086), .ZN(n15865) );
  INV_X1 U9693 ( .A(n15865), .ZN(n15866) );
  INV_X1 U9694 ( .A(n15867), .ZN(n15868) );
  BUF_X1 U9695 ( .A(n15871), .Z(n15869) );
  INV_X1 U9696 ( .A(n15873), .ZN(n15870) );
  INV_X1 U9697 ( .A(n15870), .ZN(n15871) );
  INV_X1 U9698 ( .A(n7085), .ZN(n15872) );
  INV_X1 U9699 ( .A(n15872), .ZN(n15873) );
  INV_X1 U9700 ( .A(n15874), .ZN(n15875) );
  BUF_X1 U9701 ( .A(n15878), .Z(n15876) );
  INV_X1 U9702 ( .A(n15880), .ZN(n15877) );
  INV_X1 U9703 ( .A(n15877), .ZN(n15878) );
  INV_X1 U9704 ( .A(n7084), .ZN(n15879) );
  INV_X1 U9705 ( .A(n15879), .ZN(n15880) );
  INV_X1 U9706 ( .A(n15881), .ZN(n15882) );
  BUF_X1 U9707 ( .A(n15885), .Z(n15883) );
  INV_X1 U9708 ( .A(n15887), .ZN(n15884) );
  INV_X1 U9709 ( .A(n15884), .ZN(n15885) );
  INV_X1 U9710 ( .A(n7083), .ZN(n15886) );
  INV_X1 U9711 ( .A(n15886), .ZN(n15887) );
  INV_X1 U9712 ( .A(n15888), .ZN(n15889) );
  BUF_X1 U9713 ( .A(n15892), .Z(n15890) );
  INV_X1 U9714 ( .A(n15894), .ZN(n15891) );
  INV_X1 U9715 ( .A(n15891), .ZN(n15892) );
  INV_X1 U9716 ( .A(n7082), .ZN(n15893) );
  INV_X1 U9717 ( .A(n15893), .ZN(n15894) );
  INV_X1 U9718 ( .A(n15895), .ZN(n15896) );
  BUF_X1 U9719 ( .A(n15899), .Z(n15897) );
  INV_X1 U9720 ( .A(n15901), .ZN(n15898) );
  INV_X1 U9721 ( .A(n15898), .ZN(n15899) );
  INV_X1 U9722 ( .A(n7081), .ZN(n15900) );
  INV_X1 U9723 ( .A(n15900), .ZN(n15901) );
  BUF_X1 U9724 ( .A(n15904), .Z(n15902) );
  INV_X1 U9725 ( .A(n15906), .ZN(n15903) );
  INV_X1 U9726 ( .A(n15903), .ZN(n15904) );
  INV_X1 U9727 ( .A(n7080), .ZN(n15905) );
  INV_X1 U9728 ( .A(n15905), .ZN(n15906) );
  BUF_X1 U9729 ( .A(n15909), .Z(n15907) );
  INV_X1 U9730 ( .A(n15911), .ZN(n15908) );
  INV_X1 U9731 ( .A(n15908), .ZN(n15909) );
  INV_X1 U9732 ( .A(n7079), .ZN(n15910) );
  INV_X1 U9733 ( .A(n15910), .ZN(n15911) );
  BUF_X1 U9734 ( .A(n15914), .Z(n15912) );
  INV_X1 U9735 ( .A(n15916), .ZN(n15913) );
  INV_X1 U9736 ( .A(n15913), .ZN(n15914) );
  INV_X1 U9737 ( .A(n7078), .ZN(n15915) );
  INV_X1 U9738 ( .A(n15915), .ZN(n15916) );
  BUF_X1 U9739 ( .A(n15919), .Z(n15917) );
  INV_X1 U9740 ( .A(n15921), .ZN(n15918) );
  INV_X1 U9741 ( .A(n15918), .ZN(n15919) );
  INV_X1 U9742 ( .A(n7077), .ZN(n15920) );
  INV_X1 U9743 ( .A(n15920), .ZN(n15921) );
  BUF_X1 U9744 ( .A(n15924), .Z(n15922) );
  INV_X1 U9745 ( .A(n15926), .ZN(n15923) );
  INV_X1 U9746 ( .A(n15923), .ZN(n15924) );
  INV_X1 U9747 ( .A(n7076), .ZN(n15925) );
  INV_X1 U9748 ( .A(n15925), .ZN(n15926) );
  BUF_X1 U9749 ( .A(n15929), .Z(n15927) );
  INV_X1 U9750 ( .A(n15931), .ZN(n15928) );
  INV_X1 U9751 ( .A(n15928), .ZN(n15929) );
  INV_X1 U9752 ( .A(n7075), .ZN(n15930) );
  INV_X1 U9753 ( .A(n15930), .ZN(n15931) );
  BUF_X1 U9754 ( .A(n15934), .Z(n15932) );
  INV_X1 U9755 ( .A(n15936), .ZN(n15933) );
  INV_X1 U9756 ( .A(n15933), .ZN(n15934) );
  INV_X1 U9757 ( .A(n7074), .ZN(n15935) );
  INV_X1 U9758 ( .A(n15935), .ZN(n15936) );
  BUF_X1 U9759 ( .A(n15939), .Z(n15937) );
  INV_X1 U9760 ( .A(n15941), .ZN(n15938) );
  INV_X1 U9761 ( .A(n15938), .ZN(n15939) );
  INV_X1 U9762 ( .A(n7073), .ZN(n15940) );
  INV_X1 U9763 ( .A(n15940), .ZN(n15941) );
  BUF_X1 U9764 ( .A(n15944), .Z(n15942) );
  INV_X1 U9765 ( .A(n15946), .ZN(n15943) );
  INV_X1 U9766 ( .A(n15943), .ZN(n15944) );
  INV_X1 U9767 ( .A(n7072), .ZN(n15945) );
  INV_X1 U9768 ( .A(n15945), .ZN(n15946) );
  BUF_X1 U9769 ( .A(n15949), .Z(n15947) );
  INV_X1 U9770 ( .A(n15951), .ZN(n15948) );
  INV_X1 U9771 ( .A(n15948), .ZN(n15949) );
  INV_X1 U9772 ( .A(n7071), .ZN(n15950) );
  INV_X1 U9773 ( .A(n15950), .ZN(n15951) );
  BUF_X1 U9774 ( .A(n15954), .Z(n15952) );
  INV_X1 U9775 ( .A(n15956), .ZN(n15953) );
  INV_X1 U9776 ( .A(n15953), .ZN(n15954) );
  INV_X1 U9777 ( .A(n7070), .ZN(n15955) );
  INV_X1 U9778 ( .A(n15955), .ZN(n15956) );
  BUF_X1 U9779 ( .A(n15959), .Z(n15957) );
  INV_X1 U9780 ( .A(n15961), .ZN(n15958) );
  INV_X1 U9781 ( .A(n15958), .ZN(n15959) );
  INV_X1 U9782 ( .A(n7069), .ZN(n15960) );
  INV_X1 U9783 ( .A(n15960), .ZN(n15961) );
  BUF_X1 U9784 ( .A(n15964), .Z(n15962) );
  INV_X1 U9785 ( .A(n15966), .ZN(n15963) );
  INV_X1 U9786 ( .A(n15963), .ZN(n15964) );
  INV_X1 U9787 ( .A(n70680), .ZN(n15965) );
  INV_X1 U9788 ( .A(n15965), .ZN(n15966) );
  BUF_X1 U9789 ( .A(n15969), .Z(n15967) );
  INV_X1 U9790 ( .A(n15971), .ZN(n15968) );
  INV_X1 U9791 ( .A(n15968), .ZN(n15969) );
  INV_X1 U9792 ( .A(n70670), .ZN(n15970) );
  INV_X1 U9793 ( .A(n15970), .ZN(n15971) );
  BUF_X1 U9794 ( .A(n15974), .Z(n15972) );
  INV_X1 U9795 ( .A(n15976), .ZN(n15973) );
  INV_X1 U9796 ( .A(n15973), .ZN(n15974) );
  INV_X1 U9797 ( .A(n70660), .ZN(n15975) );
  INV_X1 U9798 ( .A(n15975), .ZN(n15976) );
  BUF_X1 U9799 ( .A(n15979), .Z(n15977) );
  INV_X1 U9800 ( .A(n15981), .ZN(n15978) );
  INV_X1 U9801 ( .A(n15978), .ZN(n15979) );
  INV_X1 U9802 ( .A(n70650), .ZN(n15980) );
  INV_X1 U9803 ( .A(n15980), .ZN(n15981) );
  BUF_X1 U9804 ( .A(n15984), .Z(n15982) );
  INV_X1 U9805 ( .A(n15986), .ZN(n15983) );
  INV_X1 U9806 ( .A(n15983), .ZN(n15984) );
  INV_X1 U9807 ( .A(n70640), .ZN(n15985) );
  INV_X1 U9808 ( .A(n15985), .ZN(n15986) );
  BUF_X1 U9809 ( .A(n15989), .Z(n15987) );
  INV_X1 U9810 ( .A(n15991), .ZN(n15988) );
  INV_X1 U9811 ( .A(n15988), .ZN(n15989) );
  INV_X1 U9812 ( .A(n70630), .ZN(n15990) );
  INV_X1 U9813 ( .A(n15990), .ZN(n15991) );
  BUF_X1 U9814 ( .A(n15994), .Z(n15992) );
  INV_X1 U9815 ( .A(n15996), .ZN(n15993) );
  INV_X1 U9816 ( .A(n15993), .ZN(n15994) );
  INV_X1 U9817 ( .A(n70620), .ZN(n15995) );
  INV_X1 U9818 ( .A(n15995), .ZN(n15996) );
  BUF_X1 U9819 ( .A(n15999), .Z(n15997) );
  INV_X1 U9820 ( .A(n16001), .ZN(n15998) );
  INV_X1 U9821 ( .A(n15998), .ZN(n15999) );
  INV_X1 U9822 ( .A(n70610), .ZN(n16000) );
  INV_X1 U9823 ( .A(n16000), .ZN(n16001) );
  BUF_X1 U9824 ( .A(n16004), .Z(n16002) );
  INV_X1 U9825 ( .A(n16006), .ZN(n16003) );
  INV_X1 U9826 ( .A(n16003), .ZN(n16004) );
  INV_X1 U9827 ( .A(n70600), .ZN(n16005) );
  INV_X1 U9828 ( .A(n16005), .ZN(n16006) );
  BUF_X1 U9829 ( .A(n16009), .Z(n16007) );
  INV_X1 U9830 ( .A(n16011), .ZN(n16008) );
  INV_X1 U9831 ( .A(n16008), .ZN(n16009) );
  INV_X1 U9832 ( .A(n70590), .ZN(n16010) );
  INV_X1 U9833 ( .A(n16010), .ZN(n16011) );
  BUF_X1 U9834 ( .A(n16014), .Z(n16012) );
  INV_X1 U9835 ( .A(n16016), .ZN(n16013) );
  INV_X1 U9836 ( .A(n16013), .ZN(n16014) );
  INV_X1 U9837 ( .A(n70580), .ZN(n16015) );
  INV_X1 U9838 ( .A(n16015), .ZN(n16016) );
  BUF_X1 U9839 ( .A(n16019), .Z(n16017) );
  INV_X1 U9840 ( .A(n16021), .ZN(n16018) );
  INV_X1 U9841 ( .A(n16018), .ZN(n16019) );
  INV_X1 U9842 ( .A(n70570), .ZN(n16020) );
  INV_X1 U9843 ( .A(n16020), .ZN(n16021) );
  BUF_X1 U9844 ( .A(n16024), .Z(n16022) );
  INV_X1 U9845 ( .A(n16026), .ZN(n16023) );
  INV_X1 U9846 ( .A(n16023), .ZN(n16024) );
  INV_X1 U9847 ( .A(n70560), .ZN(n16025) );
  INV_X1 U9848 ( .A(n16025), .ZN(n16026) );
  BUF_X1 U9849 ( .A(n16029), .Z(n16027) );
  INV_X1 U9850 ( .A(n16031), .ZN(n16028) );
  INV_X1 U9851 ( .A(n16028), .ZN(n16029) );
  INV_X1 U9852 ( .A(n70550), .ZN(n16030) );
  INV_X1 U9853 ( .A(n16030), .ZN(n16031) );
  BUF_X1 U9854 ( .A(n16034), .Z(n16032) );
  INV_X1 U9855 ( .A(n16036), .ZN(n16033) );
  INV_X1 U9856 ( .A(n16033), .ZN(n16034) );
  INV_X1 U9857 ( .A(n70540), .ZN(n16035) );
  INV_X1 U9858 ( .A(n16035), .ZN(n16036) );
  BUF_X1 U9859 ( .A(n16039), .Z(n16037) );
  INV_X1 U9860 ( .A(n16041), .ZN(n16038) );
  INV_X1 U9861 ( .A(n16038), .ZN(n16039) );
  INV_X1 U9862 ( .A(n70530), .ZN(n16040) );
  INV_X1 U9863 ( .A(n16040), .ZN(n16041) );
  BUF_X1 U9864 ( .A(n16044), .Z(n16042) );
  INV_X1 U9865 ( .A(n16046), .ZN(n16043) );
  INV_X1 U9866 ( .A(n16043), .ZN(n16044) );
  INV_X1 U9867 ( .A(n70520), .ZN(n16045) );
  INV_X1 U9868 ( .A(n16045), .ZN(n16046) );
  BUF_X1 U9869 ( .A(n16049), .Z(n16047) );
  INV_X1 U9870 ( .A(n16051), .ZN(n16048) );
  INV_X1 U9871 ( .A(n16048), .ZN(n16049) );
  INV_X1 U9872 ( .A(n70510), .ZN(n16050) );
  INV_X1 U9873 ( .A(n16050), .ZN(n16051) );
  BUF_X1 U9874 ( .A(n16054), .Z(n16052) );
  INV_X1 U9875 ( .A(n16056), .ZN(n16053) );
  INV_X1 U9876 ( .A(n16053), .ZN(n16054) );
  INV_X1 U9877 ( .A(n70500), .ZN(n16055) );
  INV_X1 U9878 ( .A(n16055), .ZN(n16056) );
  BUF_X1 U9879 ( .A(n16059), .Z(n16057) );
  INV_X1 U9880 ( .A(n16061), .ZN(n16058) );
  INV_X1 U9881 ( .A(n16058), .ZN(n16059) );
  INV_X1 U9882 ( .A(n70490), .ZN(n16060) );
  INV_X1 U9883 ( .A(n16060), .ZN(n16061) );
  BUF_X1 U9884 ( .A(n16064), .Z(n16062) );
  INV_X1 U9885 ( .A(n16066), .ZN(n16063) );
  INV_X1 U9886 ( .A(n16063), .ZN(n16064) );
  INV_X1 U9887 ( .A(n70480), .ZN(n16065) );
  INV_X1 U9888 ( .A(n16065), .ZN(n16066) );
  BUF_X1 U9889 ( .A(n16069), .Z(n16067) );
  INV_X1 U9890 ( .A(n16071), .ZN(n16068) );
  INV_X1 U9891 ( .A(n16068), .ZN(n16069) );
  INV_X1 U9892 ( .A(n7047), .ZN(n16070) );
  INV_X1 U9893 ( .A(n16070), .ZN(n16071) );
  BUF_X1 U9894 ( .A(n16074), .Z(n16072) );
  INV_X1 U9895 ( .A(n16076), .ZN(n16073) );
  INV_X1 U9896 ( .A(n16073), .ZN(n16074) );
  INV_X1 U9897 ( .A(n7046), .ZN(n16075) );
  INV_X1 U9898 ( .A(n16075), .ZN(n16076) );
  BUF_X1 U9899 ( .A(n16079), .Z(n16077) );
  INV_X1 U9900 ( .A(n16081), .ZN(n16078) );
  INV_X1 U9901 ( .A(n16078), .ZN(n16079) );
  INV_X1 U9902 ( .A(n7045), .ZN(n16080) );
  INV_X1 U9903 ( .A(n16080), .ZN(n16081) );
  BUF_X1 U9904 ( .A(n16084), .Z(n16082) );
  INV_X1 U9905 ( .A(n16086), .ZN(n16083) );
  INV_X1 U9906 ( .A(n16083), .ZN(n16084) );
  INV_X1 U9907 ( .A(n7044), .ZN(n16085) );
  INV_X1 U9908 ( .A(n16085), .ZN(n16086) );
  BUF_X1 U9909 ( .A(n16089), .Z(n16087) );
  INV_X1 U9910 ( .A(n16091), .ZN(n16088) );
  INV_X1 U9911 ( .A(n16088), .ZN(n16089) );
  INV_X1 U9912 ( .A(n7043), .ZN(n16090) );
  INV_X1 U9913 ( .A(n16090), .ZN(n16091) );
  BUF_X1 U9914 ( .A(n16094), .Z(n16092) );
  INV_X1 U9915 ( .A(n16096), .ZN(n16093) );
  INV_X1 U9916 ( .A(n16093), .ZN(n16094) );
  INV_X1 U9917 ( .A(n7042), .ZN(n16095) );
  INV_X1 U9918 ( .A(n16095), .ZN(n16096) );
  BUF_X1 U9919 ( .A(n16099), .Z(n16097) );
  INV_X1 U9920 ( .A(n16101), .ZN(n16098) );
  INV_X1 U9921 ( .A(n16098), .ZN(n16099) );
  INV_X1 U9922 ( .A(n7041), .ZN(n16100) );
  INV_X1 U9923 ( .A(n16100), .ZN(n16101) );
  BUF_X1 U9924 ( .A(n16104), .Z(n16102) );
  INV_X1 U9925 ( .A(n16106), .ZN(n16103) );
  INV_X1 U9926 ( .A(n16103), .ZN(n16104) );
  INV_X1 U9927 ( .A(n7040), .ZN(n16105) );
  INV_X1 U9928 ( .A(n16105), .ZN(n16106) );
  BUF_X1 U9929 ( .A(n16109), .Z(n16107) );
  INV_X1 U9930 ( .A(n16111), .ZN(n16108) );
  INV_X1 U9931 ( .A(n16108), .ZN(n16109) );
  INV_X1 U9932 ( .A(n7039), .ZN(n16110) );
  INV_X1 U9933 ( .A(n16110), .ZN(n16111) );
  BUF_X1 U9934 ( .A(n16114), .Z(n16112) );
  INV_X1 U9935 ( .A(n16116), .ZN(n16113) );
  INV_X1 U9936 ( .A(n16113), .ZN(n16114) );
  INV_X1 U9937 ( .A(n7038), .ZN(n16115) );
  INV_X1 U9938 ( .A(n16115), .ZN(n16116) );
  BUF_X1 U9939 ( .A(n16119), .Z(n16117) );
  INV_X1 U9940 ( .A(n16121), .ZN(n16118) );
  INV_X1 U9941 ( .A(n16118), .ZN(n16119) );
  INV_X1 U9942 ( .A(n7037), .ZN(n16120) );
  INV_X1 U9943 ( .A(n16120), .ZN(n16121) );
  BUF_X1 U9944 ( .A(n16124), .Z(n16122) );
  INV_X1 U9945 ( .A(n16126), .ZN(n16123) );
  INV_X1 U9946 ( .A(n16123), .ZN(n16124) );
  INV_X1 U9947 ( .A(n7036), .ZN(n16125) );
  INV_X1 U9948 ( .A(n16125), .ZN(n16126) );
  BUF_X1 U9949 ( .A(n16129), .Z(n16127) );
  INV_X1 U9950 ( .A(n16131), .ZN(n16128) );
  INV_X1 U9951 ( .A(n16128), .ZN(n16129) );
  INV_X1 U9952 ( .A(n7035), .ZN(n16130) );
  INV_X1 U9953 ( .A(n16130), .ZN(n16131) );
  BUF_X1 U9954 ( .A(n16134), .Z(n16132) );
  INV_X1 U9955 ( .A(n16136), .ZN(n16133) );
  INV_X1 U9956 ( .A(n16133), .ZN(n16134) );
  INV_X1 U9957 ( .A(n7034), .ZN(n16135) );
  INV_X1 U9958 ( .A(n16135), .ZN(n16136) );
  INV_X1 U9959 ( .A(n1060), .ZN(n16166) );
  BUF_X1 U9960 ( .A(n16167), .Z(n16137) );
  INV_X1 U9961 ( .A(n7033), .ZN(n16138) );
  INV_X1 U9962 ( .A(n16138), .ZN(n16139) );
  INV_X1 U9963 ( .A(n1059), .ZN(n16173) );
  BUF_X1 U9964 ( .A(n16174), .Z(n16140) );
  INV_X1 U9965 ( .A(n7032), .ZN(n16141) );
  INV_X1 U9966 ( .A(n16141), .ZN(n16142) );
  INV_X1 U9967 ( .A(n1058), .ZN(n16180) );
  BUF_X1 U9968 ( .A(n16181), .Z(n16143) );
  INV_X1 U9969 ( .A(n7031), .ZN(n16144) );
  INV_X1 U9970 ( .A(n16144), .ZN(n16145) );
  INV_X1 U9971 ( .A(n1057), .ZN(n16187) );
  BUF_X1 U9972 ( .A(n16188), .Z(n16146) );
  INV_X1 U9973 ( .A(n70300), .ZN(n16147) );
  INV_X1 U9974 ( .A(n16147), .ZN(n16148) );
  INV_X1 U9975 ( .A(n1056), .ZN(n16194) );
  BUF_X1 U9976 ( .A(n16195), .Z(n16149) );
  INV_X1 U9977 ( .A(n70290), .ZN(n16150) );
  INV_X1 U9978 ( .A(n16150), .ZN(n16151) );
  INV_X1 U9979 ( .A(n1055), .ZN(n16201) );
  BUF_X1 U9980 ( .A(n16202), .Z(n16152) );
  INV_X1 U9981 ( .A(n70280), .ZN(n16153) );
  INV_X1 U9982 ( .A(n16153), .ZN(n16154) );
  INV_X1 U9983 ( .A(n1054), .ZN(n16208) );
  BUF_X1 U9984 ( .A(n16209), .Z(n16155) );
  INV_X1 U9985 ( .A(n70270), .ZN(n16156) );
  INV_X1 U9986 ( .A(n16156), .ZN(n16157) );
  INV_X1 U9987 ( .A(n1053), .ZN(n16215) );
  BUF_X1 U9988 ( .A(n16216), .Z(n16158) );
  INV_X1 U9989 ( .A(n70260), .ZN(n16159) );
  INV_X1 U9990 ( .A(n16159), .ZN(n16160) );
  BUF_X1 U9991 ( .A(n16163), .Z(n16161) );
  INV_X1 U9992 ( .A(n16165), .ZN(n16162) );
  INV_X1 U9993 ( .A(n16162), .ZN(n16163) );
  INV_X1 U9994 ( .A(n70250), .ZN(n16164) );
  INV_X1 U9995 ( .A(n16164), .ZN(n16165) );
  INV_X1 U9996 ( .A(n16166), .ZN(n16167) );
  BUF_X1 U9997 ( .A(n16170), .Z(n16168) );
  INV_X1 U9998 ( .A(n16172), .ZN(n16169) );
  INV_X1 U9999 ( .A(n16169), .ZN(n16170) );
  INV_X1 U10000 ( .A(n70240), .ZN(n16171) );
  INV_X1 U10001 ( .A(n16171), .ZN(n16172) );
  INV_X1 U10002 ( .A(n16173), .ZN(n16174) );
  BUF_X1 U10003 ( .A(n16177), .Z(n16175) );
  INV_X1 U10004 ( .A(n16179), .ZN(n16176) );
  INV_X1 U10005 ( .A(n16176), .ZN(n16177) );
  INV_X1 U10006 ( .A(n70230), .ZN(n16178) );
  INV_X1 U10007 ( .A(n16178), .ZN(n16179) );
  INV_X1 U10008 ( .A(n16180), .ZN(n16181) );
  BUF_X1 U10009 ( .A(n16184), .Z(n16182) );
  INV_X1 U10010 ( .A(n16186), .ZN(n16183) );
  INV_X1 U10011 ( .A(n16183), .ZN(n16184) );
  INV_X1 U10012 ( .A(n70220), .ZN(n16185) );
  INV_X1 U10013 ( .A(n16185), .ZN(n16186) );
  INV_X1 U10014 ( .A(n16187), .ZN(n16188) );
  BUF_X1 U10015 ( .A(n16191), .Z(n16189) );
  INV_X1 U10016 ( .A(n16193), .ZN(n16190) );
  INV_X1 U10017 ( .A(n16190), .ZN(n16191) );
  INV_X1 U10018 ( .A(n70210), .ZN(n16192) );
  INV_X1 U10019 ( .A(n16192), .ZN(n16193) );
  INV_X1 U10020 ( .A(n16194), .ZN(n16195) );
  BUF_X1 U10021 ( .A(n16198), .Z(n16196) );
  INV_X1 U10022 ( .A(n16200), .ZN(n16197) );
  INV_X1 U10023 ( .A(n16197), .ZN(n16198) );
  INV_X1 U10024 ( .A(n70200), .ZN(n16199) );
  INV_X1 U10025 ( .A(n16199), .ZN(n16200) );
  INV_X1 U10026 ( .A(n16201), .ZN(n16202) );
  BUF_X1 U10027 ( .A(n16205), .Z(n16203) );
  INV_X1 U10028 ( .A(n16207), .ZN(n16204) );
  INV_X1 U10029 ( .A(n16204), .ZN(n16205) );
  INV_X1 U10030 ( .A(n70190), .ZN(n16206) );
  INV_X1 U10031 ( .A(n16206), .ZN(n16207) );
  INV_X1 U10032 ( .A(n16208), .ZN(n16209) );
  BUF_X1 U10033 ( .A(n16212), .Z(n16210) );
  INV_X1 U10034 ( .A(n16214), .ZN(n16211) );
  INV_X1 U10035 ( .A(n16211), .ZN(n16212) );
  INV_X1 U10036 ( .A(n70180), .ZN(n16213) );
  INV_X1 U10037 ( .A(n16213), .ZN(n16214) );
  INV_X1 U10038 ( .A(n16215), .ZN(n16216) );
  BUF_X1 U10039 ( .A(n16219), .Z(n16217) );
  INV_X1 U10040 ( .A(n16221), .ZN(n16218) );
  INV_X1 U10041 ( .A(n16218), .ZN(n16219) );
  INV_X1 U10042 ( .A(n70170), .ZN(n16220) );
  INV_X1 U10043 ( .A(n16220), .ZN(n16221) );
  BUF_X1 U10044 ( .A(n16224), .Z(n16222) );
  INV_X1 U10045 ( .A(n16226), .ZN(n16223) );
  INV_X1 U10046 ( .A(n16223), .ZN(n16224) );
  INV_X1 U10047 ( .A(n70160), .ZN(n16225) );
  INV_X1 U10048 ( .A(n16225), .ZN(n16226) );
  BUF_X1 U10049 ( .A(n16229), .Z(n16227) );
  INV_X1 U10050 ( .A(n16231), .ZN(n16228) );
  INV_X1 U10051 ( .A(n16228), .ZN(n16229) );
  INV_X1 U10052 ( .A(n70150), .ZN(n16230) );
  INV_X1 U10053 ( .A(n16230), .ZN(n16231) );
  BUF_X1 U10054 ( .A(n16234), .Z(n16232) );
  INV_X1 U10055 ( .A(n16236), .ZN(n16233) );
  INV_X1 U10056 ( .A(n16233), .ZN(n16234) );
  INV_X1 U10057 ( .A(n7014), .ZN(n16235) );
  INV_X1 U10058 ( .A(n16235), .ZN(n16236) );
  BUF_X1 U10059 ( .A(n16239), .Z(n16237) );
  INV_X1 U10060 ( .A(n16241), .ZN(n16238) );
  INV_X1 U10061 ( .A(n16238), .ZN(n16239) );
  INV_X1 U10062 ( .A(n7013), .ZN(n16240) );
  INV_X1 U10063 ( .A(n16240), .ZN(n16241) );
  BUF_X1 U10064 ( .A(n16244), .Z(n16242) );
  INV_X1 U10065 ( .A(n16246), .ZN(n16243) );
  INV_X1 U10066 ( .A(n16243), .ZN(n16244) );
  INV_X1 U10067 ( .A(n7012), .ZN(n16245) );
  INV_X1 U10068 ( .A(n16245), .ZN(n16246) );
  BUF_X1 U10069 ( .A(n16249), .Z(n16247) );
  INV_X1 U10070 ( .A(n16251), .ZN(n16248) );
  INV_X1 U10071 ( .A(n16248), .ZN(n16249) );
  INV_X1 U10072 ( .A(n7011), .ZN(n16250) );
  INV_X1 U10073 ( .A(n16250), .ZN(n16251) );
  BUF_X1 U10074 ( .A(n16254), .Z(n16252) );
  INV_X1 U10075 ( .A(n16256), .ZN(n16253) );
  INV_X1 U10076 ( .A(n16253), .ZN(n16254) );
  INV_X1 U10077 ( .A(n7010), .ZN(n16255) );
  INV_X1 U10078 ( .A(n16255), .ZN(n16256) );
  BUF_X1 U10079 ( .A(n16259), .Z(n16257) );
  INV_X1 U10080 ( .A(n16261), .ZN(n16258) );
  INV_X1 U10081 ( .A(n16258), .ZN(n16259) );
  INV_X1 U10082 ( .A(n7009), .ZN(n16260) );
  INV_X1 U10083 ( .A(n16260), .ZN(n16261) );
  BUF_X1 U10084 ( .A(n16264), .Z(n16262) );
  INV_X1 U10085 ( .A(n16266), .ZN(n16263) );
  INV_X1 U10086 ( .A(n16263), .ZN(n16264) );
  INV_X1 U10087 ( .A(n7008), .ZN(n16265) );
  INV_X1 U10088 ( .A(n16265), .ZN(n16266) );
  BUF_X1 U10089 ( .A(n16269), .Z(n16267) );
  INV_X1 U10090 ( .A(n16271), .ZN(n16268) );
  INV_X1 U10091 ( .A(n16268), .ZN(n16269) );
  INV_X1 U10092 ( .A(n7007), .ZN(n16270) );
  INV_X1 U10093 ( .A(n16270), .ZN(n16271) );
  BUF_X1 U10094 ( .A(n16274), .Z(n16272) );
  INV_X1 U10095 ( .A(n16276), .ZN(n16273) );
  INV_X1 U10096 ( .A(n16273), .ZN(n16274) );
  INV_X1 U10097 ( .A(n7006), .ZN(n16275) );
  INV_X1 U10098 ( .A(n16275), .ZN(n16276) );
  BUF_X1 U10099 ( .A(n16279), .Z(n16277) );
  INV_X1 U10100 ( .A(n16281), .ZN(n16278) );
  INV_X1 U10101 ( .A(n16278), .ZN(n16279) );
  INV_X1 U10102 ( .A(n7005), .ZN(n16280) );
  INV_X1 U10103 ( .A(n16280), .ZN(n16281) );
  BUF_X1 U10104 ( .A(n16284), .Z(n16282) );
  INV_X1 U10105 ( .A(n16286), .ZN(n16283) );
  INV_X1 U10106 ( .A(n16283), .ZN(n16284) );
  INV_X1 U10107 ( .A(n7004), .ZN(n16285) );
  INV_X1 U10108 ( .A(n16285), .ZN(n16286) );
  BUF_X1 U10109 ( .A(n16289), .Z(n16287) );
  INV_X1 U10110 ( .A(n16291), .ZN(n16288) );
  INV_X1 U10111 ( .A(n16288), .ZN(n16289) );
  INV_X1 U10112 ( .A(n7003), .ZN(n16290) );
  INV_X1 U10113 ( .A(n16290), .ZN(n16291) );
  BUF_X1 U10114 ( .A(n16294), .Z(n16292) );
  INV_X1 U10115 ( .A(n16296), .ZN(n16293) );
  INV_X1 U10116 ( .A(n16293), .ZN(n16294) );
  INV_X1 U10117 ( .A(n7002), .ZN(n16295) );
  INV_X1 U10118 ( .A(n16295), .ZN(n16296) );
  BUF_X1 U10119 ( .A(n16299), .Z(n16297) );
  INV_X1 U10120 ( .A(n16301), .ZN(n16298) );
  INV_X1 U10121 ( .A(n16298), .ZN(n16299) );
  INV_X1 U10122 ( .A(n7001), .ZN(n16300) );
  INV_X1 U10123 ( .A(n16300), .ZN(n16301) );
  BUF_X1 U10124 ( .A(n16304), .Z(n16302) );
  INV_X1 U10125 ( .A(n16306), .ZN(n16303) );
  INV_X1 U10126 ( .A(n16303), .ZN(n16304) );
  INV_X1 U10127 ( .A(n7000), .ZN(n16305) );
  INV_X1 U10128 ( .A(n16305), .ZN(n16306) );
  BUF_X1 U10129 ( .A(n16309), .Z(n16307) );
  INV_X1 U10130 ( .A(n16311), .ZN(n16308) );
  INV_X1 U10131 ( .A(n16308), .ZN(n16309) );
  INV_X1 U10132 ( .A(n6999), .ZN(n16310) );
  INV_X1 U10133 ( .A(n16310), .ZN(n16311) );
  BUF_X1 U10134 ( .A(n16314), .Z(n16312) );
  INV_X1 U10135 ( .A(n16316), .ZN(n16313) );
  INV_X1 U10136 ( .A(n16313), .ZN(n16314) );
  INV_X1 U10137 ( .A(n6998), .ZN(n16315) );
  INV_X1 U10138 ( .A(n16315), .ZN(n16316) );
  BUF_X1 U10139 ( .A(n16319), .Z(n16317) );
  INV_X1 U10140 ( .A(n16321), .ZN(n16318) );
  INV_X1 U10141 ( .A(n16318), .ZN(n16319) );
  INV_X1 U10142 ( .A(n6997), .ZN(n16320) );
  INV_X1 U10143 ( .A(n16320), .ZN(n16321) );
  BUF_X1 U10144 ( .A(n16324), .Z(n16322) );
  INV_X1 U10145 ( .A(n16326), .ZN(n16323) );
  INV_X1 U10146 ( .A(n16323), .ZN(n16324) );
  INV_X1 U10147 ( .A(n6996), .ZN(n16325) );
  INV_X1 U10148 ( .A(n16325), .ZN(n16326) );
  BUF_X1 U10149 ( .A(n16329), .Z(n16327) );
  INV_X1 U10150 ( .A(n16331), .ZN(n16328) );
  INV_X1 U10151 ( .A(n16328), .ZN(n16329) );
  INV_X1 U10152 ( .A(n6995), .ZN(n16330) );
  INV_X1 U10153 ( .A(n16330), .ZN(n16331) );
  BUF_X1 U10154 ( .A(n16334), .Z(n16332) );
  INV_X1 U10155 ( .A(n16336), .ZN(n16333) );
  INV_X1 U10156 ( .A(n16333), .ZN(n16334) );
  INV_X1 U10157 ( .A(n6994), .ZN(n16335) );
  INV_X1 U10158 ( .A(n16335), .ZN(n16336) );
  BUF_X1 U10159 ( .A(n16339), .Z(n16337) );
  INV_X1 U10160 ( .A(n16341), .ZN(n16338) );
  INV_X1 U10161 ( .A(n16338), .ZN(n16339) );
  INV_X1 U10162 ( .A(n6993), .ZN(n16340) );
  INV_X1 U10163 ( .A(n16340), .ZN(n16341) );
  BUF_X1 U10164 ( .A(n16344), .Z(n16342) );
  INV_X1 U10165 ( .A(n16346), .ZN(n16343) );
  INV_X1 U10166 ( .A(n16343), .ZN(n16344) );
  INV_X1 U10167 ( .A(n6992), .ZN(n16345) );
  INV_X1 U10168 ( .A(n16345), .ZN(n16346) );
  BUF_X1 U10169 ( .A(n16349), .Z(n16347) );
  INV_X1 U10170 ( .A(n16351), .ZN(n16348) );
  INV_X1 U10171 ( .A(n16348), .ZN(n16349) );
  INV_X1 U10172 ( .A(n6991), .ZN(n16350) );
  INV_X1 U10173 ( .A(n16350), .ZN(n16351) );
  BUF_X1 U10174 ( .A(n16354), .Z(n16352) );
  INV_X1 U10175 ( .A(n16356), .ZN(n16353) );
  INV_X1 U10176 ( .A(n16353), .ZN(n16354) );
  INV_X1 U10177 ( .A(n6990), .ZN(n16355) );
  INV_X1 U10178 ( .A(n16355), .ZN(n16356) );
  BUF_X1 U10179 ( .A(n16359), .Z(n16357) );
  INV_X1 U10180 ( .A(n16361), .ZN(n16358) );
  INV_X1 U10181 ( .A(n16358), .ZN(n16359) );
  INV_X1 U10182 ( .A(n6989), .ZN(n16360) );
  INV_X1 U10183 ( .A(n16360), .ZN(n16361) );
  BUF_X1 U10184 ( .A(n16364), .Z(n16362) );
  INV_X1 U10185 ( .A(n16366), .ZN(n16363) );
  INV_X1 U10186 ( .A(n16363), .ZN(n16364) );
  INV_X1 U10187 ( .A(n6988), .ZN(n16365) );
  INV_X1 U10188 ( .A(n16365), .ZN(n16366) );
  BUF_X1 U10189 ( .A(n16369), .Z(n16367) );
  INV_X1 U10190 ( .A(n16371), .ZN(n16368) );
  INV_X1 U10191 ( .A(n16368), .ZN(n16369) );
  INV_X1 U10192 ( .A(n6987), .ZN(n16370) );
  INV_X1 U10193 ( .A(n16370), .ZN(n16371) );
  BUF_X1 U10194 ( .A(n16374), .Z(n16372) );
  INV_X1 U10195 ( .A(n16376), .ZN(n16373) );
  INV_X1 U10196 ( .A(n16373), .ZN(n16374) );
  INV_X1 U10197 ( .A(n6986), .ZN(n16375) );
  INV_X1 U10198 ( .A(n16375), .ZN(n16376) );
  BUF_X1 U10199 ( .A(n16379), .Z(n16377) );
  INV_X1 U10200 ( .A(n16381), .ZN(n16378) );
  INV_X1 U10201 ( .A(n16378), .ZN(n16379) );
  INV_X1 U10202 ( .A(n6985), .ZN(n16380) );
  INV_X1 U10203 ( .A(n16380), .ZN(n16381) );
  BUF_X1 U10204 ( .A(n16384), .Z(n16382) );
  INV_X1 U10205 ( .A(n16386), .ZN(n16383) );
  INV_X1 U10206 ( .A(n16383), .ZN(n16384) );
  INV_X1 U10207 ( .A(n6984), .ZN(n16385) );
  INV_X1 U10208 ( .A(n16385), .ZN(n16386) );
  BUF_X1 U10209 ( .A(n16389), .Z(n16387) );
  INV_X1 U10210 ( .A(n16391), .ZN(n16388) );
  INV_X1 U10211 ( .A(n16388), .ZN(n16389) );
  INV_X1 U10212 ( .A(n6983), .ZN(n16390) );
  INV_X1 U10213 ( .A(n16390), .ZN(n16391) );
  BUF_X1 U10214 ( .A(n16394), .Z(n16392) );
  INV_X1 U10215 ( .A(n16396), .ZN(n16393) );
  INV_X1 U10216 ( .A(n16393), .ZN(n16394) );
  INV_X1 U10217 ( .A(n6982), .ZN(n16395) );
  INV_X1 U10218 ( .A(n16395), .ZN(n16396) );
  BUF_X1 U10219 ( .A(n16399), .Z(n16397) );
  INV_X1 U10220 ( .A(n16401), .ZN(n16398) );
  INV_X1 U10221 ( .A(n16398), .ZN(n16399) );
  INV_X1 U10222 ( .A(n6981), .ZN(n16400) );
  INV_X1 U10223 ( .A(n16400), .ZN(n16401) );
  BUF_X1 U10224 ( .A(n16404), .Z(n16402) );
  INV_X1 U10225 ( .A(n16406), .ZN(n16403) );
  INV_X1 U10226 ( .A(n16403), .ZN(n16404) );
  INV_X1 U10227 ( .A(n6980), .ZN(n16405) );
  INV_X1 U10228 ( .A(n16405), .ZN(n16406) );
  BUF_X1 U10229 ( .A(n16409), .Z(n16407) );
  INV_X1 U10230 ( .A(n16411), .ZN(n16408) );
  INV_X1 U10231 ( .A(n16408), .ZN(n16409) );
  INV_X1 U10232 ( .A(n6979), .ZN(n16410) );
  INV_X1 U10233 ( .A(n16410), .ZN(n16411) );
  BUF_X1 U10234 ( .A(n16414), .Z(n16412) );
  INV_X1 U10235 ( .A(n16416), .ZN(n16413) );
  INV_X1 U10236 ( .A(n16413), .ZN(n16414) );
  INV_X1 U10237 ( .A(n6978), .ZN(n16415) );
  INV_X1 U10238 ( .A(n16415), .ZN(n16416) );
  BUF_X1 U10239 ( .A(n16419), .Z(n16417) );
  INV_X1 U10240 ( .A(n16421), .ZN(n16418) );
  INV_X1 U10241 ( .A(n16418), .ZN(n16419) );
  INV_X1 U10242 ( .A(n6977), .ZN(n16420) );
  INV_X1 U10243 ( .A(n16420), .ZN(n16421) );
  BUF_X1 U10244 ( .A(n16424), .Z(n16422) );
  INV_X1 U10245 ( .A(n16426), .ZN(n16423) );
  INV_X1 U10246 ( .A(n16423), .ZN(n16424) );
  INV_X1 U10247 ( .A(n69760), .ZN(n16425) );
  INV_X1 U10248 ( .A(n16425), .ZN(n16426) );
  BUF_X1 U10249 ( .A(n16429), .Z(n16427) );
  INV_X1 U10250 ( .A(n16431), .ZN(n16428) );
  INV_X1 U10251 ( .A(n16428), .ZN(n16429) );
  INV_X1 U10252 ( .A(n69750), .ZN(n16430) );
  INV_X1 U10253 ( .A(n16430), .ZN(n16431) );
  BUF_X1 U10254 ( .A(n16434), .Z(n16432) );
  INV_X1 U10255 ( .A(n16436), .ZN(n16433) );
  INV_X1 U10256 ( .A(n16433), .ZN(n16434) );
  INV_X1 U10257 ( .A(n69740), .ZN(n16435) );
  INV_X1 U10258 ( .A(n16435), .ZN(n16436) );
  BUF_X1 U10259 ( .A(n16439), .Z(n16437) );
  INV_X1 U10260 ( .A(n16441), .ZN(n16438) );
  INV_X1 U10261 ( .A(n16438), .ZN(n16439) );
  INV_X1 U10262 ( .A(n69730), .ZN(n16440) );
  INV_X1 U10263 ( .A(n16440), .ZN(n16441) );
  BUF_X1 U10264 ( .A(n16444), .Z(n16442) );
  INV_X1 U10265 ( .A(n16446), .ZN(n16443) );
  INV_X1 U10266 ( .A(n16443), .ZN(n16444) );
  INV_X1 U10267 ( .A(n69720), .ZN(n16445) );
  INV_X1 U10268 ( .A(n16445), .ZN(n16446) );
  BUF_X1 U10269 ( .A(n16449), .Z(n16447) );
  INV_X1 U10270 ( .A(n16451), .ZN(n16448) );
  INV_X1 U10271 ( .A(n16448), .ZN(n16449) );
  INV_X1 U10272 ( .A(n69710), .ZN(n16450) );
  INV_X1 U10273 ( .A(n16450), .ZN(n16451) );
  BUF_X1 U10274 ( .A(n16454), .Z(n16452) );
  INV_X1 U10275 ( .A(n16456), .ZN(n16453) );
  INV_X1 U10276 ( .A(n16453), .ZN(n16454) );
  INV_X1 U10277 ( .A(n69700), .ZN(n16455) );
  INV_X1 U10278 ( .A(n16455), .ZN(n16456) );
  INV_X1 U10279 ( .A(n1004), .ZN(n16486) );
  BUF_X1 U10280 ( .A(n16487), .Z(n16457) );
  INV_X1 U10281 ( .A(n69690), .ZN(n16458) );
  INV_X1 U10282 ( .A(n16458), .ZN(n16459) );
  INV_X1 U10283 ( .A(n1003), .ZN(n16493) );
  BUF_X1 U10284 ( .A(n16494), .Z(n16460) );
  INV_X1 U10285 ( .A(n69680), .ZN(n16461) );
  INV_X1 U10286 ( .A(n16461), .ZN(n16462) );
  INV_X1 U10287 ( .A(n1002), .ZN(n16500) );
  BUF_X1 U10288 ( .A(n16501), .Z(n16463) );
  INV_X1 U10289 ( .A(n69670), .ZN(n16464) );
  INV_X1 U10290 ( .A(n16464), .ZN(n16465) );
  INV_X1 U10291 ( .A(n1001), .ZN(n16507) );
  BUF_X1 U10292 ( .A(n16508), .Z(n16466) );
  INV_X1 U10293 ( .A(n69660), .ZN(n16467) );
  INV_X1 U10294 ( .A(n16467), .ZN(n16468) );
  INV_X1 U10295 ( .A(n1000), .ZN(n16514) );
  BUF_X1 U10296 ( .A(n16515), .Z(n16469) );
  INV_X1 U10297 ( .A(n69650), .ZN(n16470) );
  INV_X1 U10298 ( .A(n16470), .ZN(n16471) );
  INV_X1 U10299 ( .A(n999), .ZN(n16521) );
  BUF_X1 U10300 ( .A(n16522), .Z(n16472) );
  INV_X1 U10301 ( .A(n69640), .ZN(n16473) );
  INV_X1 U10302 ( .A(n16473), .ZN(n16474) );
  INV_X1 U10303 ( .A(n998), .ZN(n16528) );
  BUF_X1 U10304 ( .A(n16529), .Z(n16475) );
  INV_X1 U10305 ( .A(n69630), .ZN(n16476) );
  INV_X1 U10306 ( .A(n16476), .ZN(n16477) );
  INV_X1 U10307 ( .A(n997), .ZN(n16535) );
  BUF_X1 U10308 ( .A(n16536), .Z(n16478) );
  INV_X1 U10309 ( .A(n69620), .ZN(n16479) );
  INV_X1 U10310 ( .A(n16479), .ZN(n16480) );
  BUF_X1 U10311 ( .A(n16483), .Z(n16481) );
  INV_X1 U10312 ( .A(n16485), .ZN(n16482) );
  INV_X1 U10313 ( .A(n16482), .ZN(n16483) );
  INV_X1 U10314 ( .A(n69610), .ZN(n16484) );
  INV_X1 U10315 ( .A(n16484), .ZN(n16485) );
  INV_X1 U10316 ( .A(n16486), .ZN(n16487) );
  BUF_X1 U10317 ( .A(n16490), .Z(n16488) );
  INV_X1 U10318 ( .A(n16492), .ZN(n16489) );
  INV_X1 U10319 ( .A(n16489), .ZN(n16490) );
  INV_X1 U10320 ( .A(n69600), .ZN(n16491) );
  INV_X1 U10321 ( .A(n16491), .ZN(n16492) );
  INV_X1 U10322 ( .A(n16493), .ZN(n16494) );
  BUF_X1 U10323 ( .A(n16497), .Z(n16495) );
  INV_X1 U10324 ( .A(n16499), .ZN(n16496) );
  INV_X1 U10325 ( .A(n16496), .ZN(n16497) );
  INV_X1 U10326 ( .A(n69590), .ZN(n16498) );
  INV_X1 U10327 ( .A(n16498), .ZN(n16499) );
  INV_X1 U10328 ( .A(n16500), .ZN(n16501) );
  BUF_X1 U10329 ( .A(n16504), .Z(n16502) );
  INV_X1 U10330 ( .A(n16506), .ZN(n16503) );
  INV_X1 U10331 ( .A(n16503), .ZN(n16504) );
  INV_X1 U10332 ( .A(n69580), .ZN(n16505) );
  INV_X1 U10333 ( .A(n16505), .ZN(n16506) );
  INV_X1 U10334 ( .A(n16507), .ZN(n16508) );
  BUF_X1 U10335 ( .A(n16511), .Z(n16509) );
  INV_X1 U10336 ( .A(n16513), .ZN(n16510) );
  INV_X1 U10337 ( .A(n16510), .ZN(n16511) );
  INV_X1 U10338 ( .A(n69570), .ZN(n16512) );
  INV_X1 U10339 ( .A(n16512), .ZN(n16513) );
  INV_X1 U10340 ( .A(n16514), .ZN(n16515) );
  BUF_X1 U10341 ( .A(n16518), .Z(n16516) );
  INV_X1 U10342 ( .A(n16520), .ZN(n16517) );
  INV_X1 U10343 ( .A(n16517), .ZN(n16518) );
  INV_X1 U10344 ( .A(n69560), .ZN(n16519) );
  INV_X1 U10345 ( .A(n16519), .ZN(n16520) );
  INV_X1 U10346 ( .A(n16521), .ZN(n16522) );
  BUF_X1 U10347 ( .A(n16525), .Z(n16523) );
  INV_X1 U10348 ( .A(n16527), .ZN(n16524) );
  INV_X1 U10349 ( .A(n16524), .ZN(n16525) );
  INV_X1 U10350 ( .A(n6955), .ZN(n16526) );
  INV_X1 U10351 ( .A(n16526), .ZN(n16527) );
  INV_X1 U10352 ( .A(n16528), .ZN(n16529) );
  BUF_X1 U10353 ( .A(n16532), .Z(n16530) );
  INV_X1 U10354 ( .A(n16534), .ZN(n16531) );
  INV_X1 U10355 ( .A(n16531), .ZN(n16532) );
  INV_X1 U10356 ( .A(n6954), .ZN(n16533) );
  INV_X1 U10357 ( .A(n16533), .ZN(n16534) );
  INV_X1 U10358 ( .A(n16535), .ZN(n16536) );
  BUF_X1 U10359 ( .A(n16539), .Z(n16537) );
  INV_X1 U10360 ( .A(n16541), .ZN(n16538) );
  INV_X1 U10361 ( .A(n16538), .ZN(n16539) );
  INV_X1 U10362 ( .A(n6953), .ZN(n16540) );
  INV_X1 U10363 ( .A(n16540), .ZN(n16541) );
  BUF_X1 U10364 ( .A(n16544), .Z(n16542) );
  INV_X1 U10365 ( .A(n16546), .ZN(n16543) );
  INV_X1 U10366 ( .A(n16543), .ZN(n16544) );
  INV_X1 U10367 ( .A(n6952), .ZN(n16545) );
  INV_X1 U10368 ( .A(n16545), .ZN(n16546) );
  BUF_X1 U10369 ( .A(n16549), .Z(n16547) );
  INV_X1 U10370 ( .A(n16551), .ZN(n16548) );
  INV_X1 U10371 ( .A(n16548), .ZN(n16549) );
  INV_X1 U10372 ( .A(n6951), .ZN(n16550) );
  INV_X1 U10373 ( .A(n16550), .ZN(n16551) );
  BUF_X1 U10374 ( .A(n16554), .Z(n16552) );
  INV_X1 U10375 ( .A(n16556), .ZN(n16553) );
  INV_X1 U10376 ( .A(n16553), .ZN(n16554) );
  INV_X1 U10377 ( .A(n6950), .ZN(n16555) );
  INV_X1 U10378 ( .A(n16555), .ZN(n16556) );
  BUF_X1 U10379 ( .A(n16559), .Z(n16557) );
  INV_X1 U10380 ( .A(n16561), .ZN(n16558) );
  INV_X1 U10381 ( .A(n16558), .ZN(n16559) );
  INV_X1 U10382 ( .A(n6949), .ZN(n16560) );
  INV_X1 U10383 ( .A(n16560), .ZN(n16561) );
  BUF_X1 U10384 ( .A(n16564), .Z(n16562) );
  INV_X1 U10385 ( .A(n16566), .ZN(n16563) );
  INV_X1 U10386 ( .A(n16563), .ZN(n16564) );
  INV_X1 U10387 ( .A(n6948), .ZN(n16565) );
  INV_X1 U10388 ( .A(n16565), .ZN(n16566) );
  BUF_X1 U10389 ( .A(n16569), .Z(n16567) );
  INV_X1 U10390 ( .A(n16571), .ZN(n16568) );
  INV_X1 U10391 ( .A(n16568), .ZN(n16569) );
  INV_X1 U10392 ( .A(n6947), .ZN(n16570) );
  INV_X1 U10393 ( .A(n16570), .ZN(n16571) );
  BUF_X1 U10394 ( .A(n16574), .Z(n16572) );
  INV_X1 U10395 ( .A(n16576), .ZN(n16573) );
  INV_X1 U10396 ( .A(n16573), .ZN(n16574) );
  INV_X1 U10397 ( .A(n6946), .ZN(n16575) );
  INV_X1 U10398 ( .A(n16575), .ZN(n16576) );
  BUF_X1 U10399 ( .A(n16579), .Z(n16577) );
  INV_X1 U10400 ( .A(n16581), .ZN(n16578) );
  INV_X1 U10401 ( .A(n16578), .ZN(n16579) );
  INV_X1 U10402 ( .A(n6945), .ZN(n16580) );
  INV_X1 U10403 ( .A(n16580), .ZN(n16581) );
  BUF_X1 U10404 ( .A(n16584), .Z(n16582) );
  INV_X1 U10405 ( .A(n16586), .ZN(n16583) );
  INV_X1 U10406 ( .A(n16583), .ZN(n16584) );
  INV_X1 U10407 ( .A(n6944), .ZN(n16585) );
  INV_X1 U10408 ( .A(n16585), .ZN(n16586) );
  BUF_X1 U10409 ( .A(n16589), .Z(n16587) );
  INV_X1 U10410 ( .A(n16591), .ZN(n16588) );
  INV_X1 U10411 ( .A(n16588), .ZN(n16589) );
  INV_X1 U10412 ( .A(n6943), .ZN(n16590) );
  INV_X1 U10413 ( .A(n16590), .ZN(n16591) );
  BUF_X1 U10414 ( .A(n16594), .Z(n16592) );
  INV_X1 U10415 ( .A(n16596), .ZN(n16593) );
  INV_X1 U10416 ( .A(n16593), .ZN(n16594) );
  INV_X1 U10417 ( .A(n6942), .ZN(n16595) );
  INV_X1 U10418 ( .A(n16595), .ZN(n16596) );
  BUF_X1 U10419 ( .A(n16599), .Z(n16597) );
  INV_X1 U10420 ( .A(n16601), .ZN(n16598) );
  INV_X1 U10421 ( .A(n16598), .ZN(n16599) );
  INV_X1 U10422 ( .A(n6941), .ZN(n16600) );
  INV_X1 U10423 ( .A(n16600), .ZN(n16601) );
  BUF_X1 U10424 ( .A(n16604), .Z(n16602) );
  INV_X1 U10425 ( .A(n16606), .ZN(n16603) );
  INV_X1 U10426 ( .A(n16603), .ZN(n16604) );
  INV_X1 U10427 ( .A(n6940), .ZN(n16605) );
  INV_X1 U10428 ( .A(n16605), .ZN(n16606) );
  BUF_X1 U10429 ( .A(n16609), .Z(n16607) );
  INV_X1 U10430 ( .A(n16611), .ZN(n16608) );
  INV_X1 U10431 ( .A(n16608), .ZN(n16609) );
  INV_X1 U10432 ( .A(n6939), .ZN(n16610) );
  INV_X1 U10433 ( .A(n16610), .ZN(n16611) );
  BUF_X1 U10434 ( .A(n16614), .Z(n16612) );
  INV_X1 U10435 ( .A(n16616), .ZN(n16613) );
  INV_X1 U10436 ( .A(n16613), .ZN(n16614) );
  INV_X1 U10437 ( .A(n69380), .ZN(n16615) );
  INV_X1 U10438 ( .A(n16615), .ZN(n16616) );
  BUF_X1 U10439 ( .A(n16619), .Z(n16617) );
  INV_X1 U10440 ( .A(n16621), .ZN(n16618) );
  INV_X1 U10441 ( .A(n16618), .ZN(n16619) );
  INV_X1 U10442 ( .A(n69370), .ZN(n16620) );
  INV_X1 U10443 ( .A(n16620), .ZN(n16621) );
  BUF_X1 U10444 ( .A(n16624), .Z(n16622) );
  INV_X1 U10445 ( .A(n16626), .ZN(n16623) );
  INV_X1 U10446 ( .A(n16623), .ZN(n16624) );
  INV_X1 U10447 ( .A(n69360), .ZN(n16625) );
  INV_X1 U10448 ( .A(n16625), .ZN(n16626) );
  BUF_X1 U10449 ( .A(n16629), .Z(n16627) );
  INV_X1 U10450 ( .A(n16631), .ZN(n16628) );
  INV_X1 U10451 ( .A(n16628), .ZN(n16629) );
  INV_X1 U10452 ( .A(n69350), .ZN(n16630) );
  INV_X1 U10453 ( .A(n16630), .ZN(n16631) );
  BUF_X1 U10454 ( .A(n16634), .Z(n16632) );
  INV_X1 U10455 ( .A(n16636), .ZN(n16633) );
  INV_X1 U10456 ( .A(n16633), .ZN(n16634) );
  INV_X1 U10457 ( .A(n69340), .ZN(n16635) );
  INV_X1 U10458 ( .A(n16635), .ZN(n16636) );
  BUF_X1 U10459 ( .A(n16639), .Z(n16637) );
  INV_X1 U10460 ( .A(n16641), .ZN(n16638) );
  INV_X1 U10461 ( .A(n16638), .ZN(n16639) );
  INV_X1 U10462 ( .A(n69330), .ZN(n16640) );
  INV_X1 U10463 ( .A(n16640), .ZN(n16641) );
  BUF_X1 U10464 ( .A(n16644), .Z(n16642) );
  INV_X1 U10465 ( .A(n16646), .ZN(n16643) );
  INV_X1 U10466 ( .A(n16643), .ZN(n16644) );
  INV_X1 U10467 ( .A(n69320), .ZN(n16645) );
  INV_X1 U10468 ( .A(n16645), .ZN(n16646) );
  BUF_X1 U10469 ( .A(n16649), .Z(n16647) );
  INV_X1 U10470 ( .A(n16651), .ZN(n16648) );
  INV_X1 U10471 ( .A(n16648), .ZN(n16649) );
  INV_X1 U10472 ( .A(n69310), .ZN(n16650) );
  INV_X1 U10473 ( .A(n16650), .ZN(n16651) );
  BUF_X1 U10474 ( .A(n16654), .Z(n16652) );
  INV_X1 U10475 ( .A(n16656), .ZN(n16653) );
  INV_X1 U10476 ( .A(n16653), .ZN(n16654) );
  INV_X1 U10477 ( .A(n69300), .ZN(n16655) );
  INV_X1 U10478 ( .A(n16655), .ZN(n16656) );
  BUF_X1 U10479 ( .A(n16659), .Z(n16657) );
  INV_X1 U10480 ( .A(n16661), .ZN(n16658) );
  INV_X1 U10481 ( .A(n16658), .ZN(n16659) );
  INV_X1 U10482 ( .A(n69290), .ZN(n16660) );
  INV_X1 U10483 ( .A(n16660), .ZN(n16661) );
  BUF_X1 U10484 ( .A(n16664), .Z(n16662) );
  INV_X1 U10485 ( .A(n16666), .ZN(n16663) );
  INV_X1 U10486 ( .A(n16663), .ZN(n16664) );
  INV_X1 U10487 ( .A(n69280), .ZN(n16665) );
  INV_X1 U10488 ( .A(n16665), .ZN(n16666) );
  BUF_X1 U10489 ( .A(n16669), .Z(n16667) );
  INV_X1 U10490 ( .A(n16671), .ZN(n16668) );
  INV_X1 U10491 ( .A(n16668), .ZN(n16669) );
  INV_X1 U10492 ( .A(n69270), .ZN(n16670) );
  INV_X1 U10493 ( .A(n16670), .ZN(n16671) );
  BUF_X1 U10494 ( .A(n16674), .Z(n16672) );
  INV_X1 U10495 ( .A(n16676), .ZN(n16673) );
  INV_X1 U10496 ( .A(n16673), .ZN(n16674) );
  INV_X1 U10497 ( .A(n69260), .ZN(n16675) );
  INV_X1 U10498 ( .A(n16675), .ZN(n16676) );
  BUF_X1 U10499 ( .A(n16679), .Z(n16677) );
  INV_X1 U10500 ( .A(n16681), .ZN(n16678) );
  INV_X1 U10501 ( .A(n16678), .ZN(n16679) );
  INV_X1 U10502 ( .A(n69250), .ZN(n16680) );
  INV_X1 U10503 ( .A(n16680), .ZN(n16681) );
  BUF_X1 U10504 ( .A(n16684), .Z(n16682) );
  INV_X1 U10505 ( .A(n16686), .ZN(n16683) );
  INV_X1 U10506 ( .A(n16683), .ZN(n16684) );
  INV_X1 U10507 ( .A(n69240), .ZN(n16685) );
  INV_X1 U10508 ( .A(n16685), .ZN(n16686) );
  BUF_X1 U10509 ( .A(n16689), .Z(n16687) );
  INV_X1 U10510 ( .A(n16691), .ZN(n16688) );
  INV_X1 U10511 ( .A(n16688), .ZN(n16689) );
  INV_X1 U10512 ( .A(n69230), .ZN(n16690) );
  INV_X1 U10513 ( .A(n16690), .ZN(n16691) );
  BUF_X1 U10514 ( .A(n16694), .Z(n16692) );
  INV_X1 U10515 ( .A(n16696), .ZN(n16693) );
  INV_X1 U10516 ( .A(n16693), .ZN(n16694) );
  INV_X1 U10517 ( .A(n6922), .ZN(n16695) );
  INV_X1 U10518 ( .A(n16695), .ZN(n16696) );
  BUF_X1 U10519 ( .A(n16699), .Z(n16697) );
  INV_X1 U10520 ( .A(n16701), .ZN(n16698) );
  INV_X1 U10521 ( .A(n16698), .ZN(n16699) );
  INV_X1 U10522 ( .A(n6921), .ZN(n16700) );
  INV_X1 U10523 ( .A(n16700), .ZN(n16701) );
  BUF_X1 U10524 ( .A(n16704), .Z(n16702) );
  INV_X1 U10525 ( .A(n16706), .ZN(n16703) );
  INV_X1 U10526 ( .A(n16703), .ZN(n16704) );
  INV_X1 U10527 ( .A(n6920), .ZN(n16705) );
  INV_X1 U10528 ( .A(n16705), .ZN(n16706) );
  BUF_X1 U10529 ( .A(n16709), .Z(n16707) );
  INV_X1 U10530 ( .A(n16711), .ZN(n16708) );
  INV_X1 U10531 ( .A(n16708), .ZN(n16709) );
  INV_X1 U10532 ( .A(n6919), .ZN(n16710) );
  INV_X1 U10533 ( .A(n16710), .ZN(n16711) );
  BUF_X1 U10534 ( .A(n16714), .Z(n16712) );
  INV_X1 U10535 ( .A(n16716), .ZN(n16713) );
  INV_X1 U10536 ( .A(n16713), .ZN(n16714) );
  INV_X1 U10537 ( .A(n6918), .ZN(n16715) );
  INV_X1 U10538 ( .A(n16715), .ZN(n16716) );
  BUF_X1 U10539 ( .A(n16719), .Z(n16717) );
  INV_X1 U10540 ( .A(n16721), .ZN(n16718) );
  INV_X1 U10541 ( .A(n16718), .ZN(n16719) );
  INV_X1 U10542 ( .A(n6917), .ZN(n16720) );
  INV_X1 U10543 ( .A(n16720), .ZN(n16721) );
  BUF_X1 U10544 ( .A(n16724), .Z(n16722) );
  INV_X1 U10545 ( .A(n16726), .ZN(n16723) );
  INV_X1 U10546 ( .A(n16723), .ZN(n16724) );
  INV_X1 U10547 ( .A(n6916), .ZN(n16725) );
  INV_X1 U10548 ( .A(n16725), .ZN(n16726) );
  BUF_X1 U10549 ( .A(n16729), .Z(n16727) );
  INV_X1 U10550 ( .A(n16731), .ZN(n16728) );
  INV_X1 U10551 ( .A(n16728), .ZN(n16729) );
  INV_X1 U10552 ( .A(n6915), .ZN(n16730) );
  INV_X1 U10553 ( .A(n16730), .ZN(n16731) );
  BUF_X1 U10554 ( .A(n16734), .Z(n16732) );
  INV_X1 U10555 ( .A(n16736), .ZN(n16733) );
  INV_X1 U10556 ( .A(n16733), .ZN(n16734) );
  INV_X1 U10557 ( .A(n6914), .ZN(n16735) );
  INV_X1 U10558 ( .A(n16735), .ZN(n16736) );
  BUF_X1 U10559 ( .A(n16739), .Z(n16737) );
  INV_X1 U10560 ( .A(n16741), .ZN(n16738) );
  INV_X1 U10561 ( .A(n16738), .ZN(n16739) );
  INV_X1 U10562 ( .A(n6913), .ZN(n16740) );
  INV_X1 U10563 ( .A(n16740), .ZN(n16741) );
  BUF_X1 U10564 ( .A(n16744), .Z(n16742) );
  INV_X1 U10565 ( .A(n16746), .ZN(n16743) );
  INV_X1 U10566 ( .A(n16743), .ZN(n16744) );
  INV_X1 U10567 ( .A(n6912), .ZN(n16745) );
  INV_X1 U10568 ( .A(n16745), .ZN(n16746) );
  BUF_X1 U10569 ( .A(n16749), .Z(n16747) );
  INV_X1 U10570 ( .A(n16751), .ZN(n16748) );
  INV_X1 U10571 ( .A(n16748), .ZN(n16749) );
  INV_X1 U10572 ( .A(n6911), .ZN(n16750) );
  INV_X1 U10573 ( .A(n16750), .ZN(n16751) );
  BUF_X1 U10574 ( .A(n16754), .Z(n16752) );
  INV_X1 U10575 ( .A(n16756), .ZN(n16753) );
  INV_X1 U10576 ( .A(n16753), .ZN(n16754) );
  INV_X1 U10577 ( .A(n6910), .ZN(n16755) );
  INV_X1 U10578 ( .A(n16755), .ZN(n16756) );
  BUF_X1 U10579 ( .A(n16759), .Z(n16757) );
  INV_X1 U10580 ( .A(n16761), .ZN(n16758) );
  INV_X1 U10581 ( .A(n16758), .ZN(n16759) );
  INV_X1 U10582 ( .A(n6909), .ZN(n16760) );
  INV_X1 U10583 ( .A(n16760), .ZN(n16761) );
  BUF_X1 U10584 ( .A(n16764), .Z(n16762) );
  INV_X1 U10585 ( .A(n16766), .ZN(n16763) );
  INV_X1 U10586 ( .A(n16763), .ZN(n16764) );
  INV_X1 U10587 ( .A(n6908), .ZN(n16765) );
  INV_X1 U10588 ( .A(n16765), .ZN(n16766) );
  BUF_X1 U10589 ( .A(n16769), .Z(n16767) );
  INV_X1 U10590 ( .A(n16771), .ZN(n16768) );
  INV_X1 U10591 ( .A(n16768), .ZN(n16769) );
  INV_X1 U10592 ( .A(n6907), .ZN(n16770) );
  INV_X1 U10593 ( .A(n16770), .ZN(n16771) );
  BUF_X1 U10594 ( .A(n16774), .Z(n16772) );
  INV_X1 U10595 ( .A(n16776), .ZN(n16773) );
  INV_X1 U10596 ( .A(n16773), .ZN(n16774) );
  INV_X1 U10597 ( .A(n6906), .ZN(n16775) );
  INV_X1 U10598 ( .A(n16775), .ZN(n16776) );
  BUF_X1 U10599 ( .A(n16781), .Z(n16777) );
  INV_X1 U10600 ( .A(n2872), .ZN(n16778) );
  INV_X1 U10601 ( .A(n16778), .ZN(n16779) );
  INV_X1 U10602 ( .A(n6375), .ZN(n16780) );
  INV_X1 U10603 ( .A(n16780), .ZN(n16781) );
  BUF_X1 U10604 ( .A(n16786), .Z(n16782) );
  INV_X1 U10605 ( .A(n2873), .ZN(n16783) );
  INV_X1 U10606 ( .A(n16783), .ZN(n16784) );
  INV_X1 U10607 ( .A(n6376), .ZN(n16785) );
  INV_X1 U10608 ( .A(n16785), .ZN(n16786) );
  BUF_X1 U10609 ( .A(n16791), .Z(n16787) );
  INV_X1 U10610 ( .A(n1847), .ZN(n16788) );
  INV_X1 U10611 ( .A(n16788), .ZN(n16789) );
  INV_X1 U10612 ( .A(n54280), .ZN(n16790) );
  INV_X1 U10613 ( .A(n16790), .ZN(n16791) );
  BUF_X1 U10614 ( .A(n16796), .Z(n16792) );
  INV_X1 U10615 ( .A(n2871), .ZN(n16793) );
  INV_X1 U10616 ( .A(n16793), .ZN(n16794) );
  INV_X1 U10617 ( .A(n6374), .ZN(n16795) );
  INV_X1 U10618 ( .A(n16795), .ZN(n16796) );
  BUF_X1 U10619 ( .A(n16801), .Z(n16797) );
  INV_X1 U10620 ( .A(n1845), .ZN(n16798) );
  INV_X1 U10621 ( .A(n16798), .ZN(n16799) );
  INV_X1 U10622 ( .A(n54260), .ZN(n16800) );
  INV_X1 U10623 ( .A(n16800), .ZN(n16801) );
  BUF_X1 U10624 ( .A(n16806), .Z(n16802) );
  INV_X1 U10625 ( .A(n1846), .ZN(n16803) );
  INV_X1 U10626 ( .A(n16803), .ZN(n16804) );
  INV_X1 U10627 ( .A(n54270), .ZN(n16805) );
  INV_X1 U10628 ( .A(n16805), .ZN(n16806) );
  BUF_X1 U10629 ( .A(n16811), .Z(n16807) );
  INV_X1 U10630 ( .A(n1849), .ZN(n16808) );
  INV_X1 U10631 ( .A(n16808), .ZN(n16809) );
  INV_X1 U10632 ( .A(n54300), .ZN(n16810) );
  INV_X1 U10633 ( .A(n16810), .ZN(n16811) );
  BUF_X1 U10634 ( .A(n16816), .Z(n16812) );
  INV_X1 U10635 ( .A(n1848), .ZN(n16813) );
  INV_X1 U10636 ( .A(n16813), .ZN(n16814) );
  INV_X1 U10637 ( .A(n54290), .ZN(n16815) );
  INV_X1 U10638 ( .A(n16815), .ZN(n16816) );
  BUF_X1 U10639 ( .A(n16821), .Z(n16817) );
  INV_X1 U10640 ( .A(n1852), .ZN(n16818) );
  INV_X1 U10641 ( .A(n16818), .ZN(n16819) );
  INV_X1 U10642 ( .A(n54330), .ZN(n16820) );
  INV_X1 U10643 ( .A(n16820), .ZN(n16821) );
  BUF_X1 U10644 ( .A(n16826), .Z(n16822) );
  INV_X1 U10645 ( .A(n1851), .ZN(n16823) );
  INV_X1 U10646 ( .A(n16823), .ZN(n16824) );
  INV_X1 U10647 ( .A(n54320), .ZN(n16825) );
  INV_X1 U10648 ( .A(n16825), .ZN(n16826) );
  BUF_X1 U10649 ( .A(n16831), .Z(n16827) );
  INV_X1 U10650 ( .A(n1850), .ZN(n16828) );
  INV_X1 U10651 ( .A(n16828), .ZN(n16829) );
  INV_X1 U10652 ( .A(n54310), .ZN(n16830) );
  INV_X1 U10653 ( .A(n16830), .ZN(n16831) );
  BUF_X1 U10654 ( .A(n16836), .Z(n16832) );
  INV_X1 U10655 ( .A(n1855), .ZN(n16833) );
  INV_X1 U10656 ( .A(n16833), .ZN(n16834) );
  INV_X1 U10657 ( .A(n54360), .ZN(n16835) );
  INV_X1 U10658 ( .A(n16835), .ZN(n16836) );
  BUF_X1 U10659 ( .A(n16841), .Z(n16837) );
  INV_X1 U10660 ( .A(n1858), .ZN(n16838) );
  INV_X1 U10661 ( .A(n16838), .ZN(n16839) );
  INV_X1 U10662 ( .A(n5439), .ZN(n16840) );
  INV_X1 U10663 ( .A(n16840), .ZN(n16841) );
  BUF_X1 U10664 ( .A(n16846), .Z(n16842) );
  INV_X1 U10665 ( .A(n1853), .ZN(n16843) );
  INV_X1 U10666 ( .A(n16843), .ZN(n16844) );
  INV_X1 U10667 ( .A(n54340), .ZN(n16845) );
  INV_X1 U10668 ( .A(n16845), .ZN(n16846) );
  BUF_X1 U10669 ( .A(n16851), .Z(n16847) );
  INV_X1 U10670 ( .A(n1854), .ZN(n16848) );
  INV_X1 U10671 ( .A(n16848), .ZN(n16849) );
  INV_X1 U10672 ( .A(n54350), .ZN(n16850) );
  INV_X1 U10673 ( .A(n16850), .ZN(n16851) );
  BUF_X1 U10674 ( .A(n16856), .Z(n16852) );
  INV_X1 U10675 ( .A(n28610), .ZN(n16853) );
  INV_X1 U10676 ( .A(n16853), .ZN(n16854) );
  INV_X1 U10677 ( .A(n63640), .ZN(n16855) );
  INV_X1 U10678 ( .A(n16855), .ZN(n16856) );
  BUF_X1 U10679 ( .A(n16861), .Z(n16857) );
  INV_X1 U10680 ( .A(n1856), .ZN(n16858) );
  INV_X1 U10681 ( .A(n16858), .ZN(n16859) );
  INV_X1 U10682 ( .A(n54370), .ZN(n16860) );
  INV_X1 U10683 ( .A(n16860), .ZN(n16861) );
  BUF_X1 U10684 ( .A(n16866), .Z(n16862) );
  INV_X1 U10685 ( .A(n1857), .ZN(n16863) );
  INV_X1 U10686 ( .A(n16863), .ZN(n16864) );
  INV_X1 U10687 ( .A(n54380), .ZN(n16865) );
  INV_X1 U10688 ( .A(n16865), .ZN(n16866) );
  BUF_X1 U10689 ( .A(n16871), .Z(n16867) );
  INV_X1 U10690 ( .A(n274700), .ZN(n16868) );
  INV_X1 U10691 ( .A(n16868), .ZN(n16869) );
  INV_X1 U10692 ( .A(n62620), .ZN(n16870) );
  INV_X1 U10693 ( .A(n16870), .ZN(n16871) );
  BUF_X1 U10694 ( .A(n16875), .Z(n16872) );
  INV_X1 U10695 ( .A(matrix_mul_2D_0__0__0_), .ZN(n16873) );
  INV_X1 U10696 ( .A(n5440), .ZN(n16874) );
  INV_X1 U10697 ( .A(n16874), .ZN(n16875) );
  BUF_X1 U10698 ( .A(n16880), .Z(n16876) );
  INV_X1 U10699 ( .A(n28600), .ZN(n16877) );
  INV_X1 U10700 ( .A(n16877), .ZN(n16878) );
  INV_X1 U10701 ( .A(n63630), .ZN(n16879) );
  INV_X1 U10702 ( .A(n16879), .ZN(n16880) );
  BUF_X1 U10703 ( .A(n16884), .Z(n16881) );
  INV_X1 U10704 ( .A(matrix_mul_2D_6__7__0_), .ZN(n16882) );
  INV_X1 U10705 ( .A(n62650), .ZN(n16883) );
  INV_X1 U10706 ( .A(n16883), .ZN(n16884) );
  BUF_X1 U10707 ( .A(n16889), .Z(n16885) );
  INV_X1 U10708 ( .A(n28650), .ZN(n16886) );
  INV_X1 U10709 ( .A(n16886), .ZN(n16887) );
  INV_X1 U10710 ( .A(n63680), .ZN(n16888) );
  INV_X1 U10711 ( .A(n16888), .ZN(n16889) );
  BUF_X1 U10712 ( .A(n16894), .Z(n16890) );
  INV_X1 U10713 ( .A(n274500), .ZN(n16891) );
  INV_X1 U10714 ( .A(n16891), .ZN(n16892) );
  INV_X1 U10715 ( .A(n6260), .ZN(n16893) );
  INV_X1 U10716 ( .A(n16893), .ZN(n16894) );
  BUF_X1 U10717 ( .A(n16899), .Z(n16895) );
  INV_X1 U10718 ( .A(n28580), .ZN(n16896) );
  INV_X1 U10719 ( .A(n16896), .ZN(n16897) );
  INV_X1 U10720 ( .A(n63610), .ZN(n16898) );
  INV_X1 U10721 ( .A(n16898), .ZN(n16899) );
  BUF_X1 U10722 ( .A(n16904), .Z(n16900) );
  INV_X1 U10723 ( .A(n28620), .ZN(n16901) );
  INV_X1 U10724 ( .A(n16901), .ZN(n16902) );
  INV_X1 U10725 ( .A(n63650), .ZN(n16903) );
  INV_X1 U10726 ( .A(n16903), .ZN(n16904) );
  BUF_X1 U10727 ( .A(n16909), .Z(n16905) );
  INV_X1 U10728 ( .A(n274800), .ZN(n16906) );
  INV_X1 U10729 ( .A(n16906), .ZN(n16907) );
  INV_X1 U10730 ( .A(n62630), .ZN(n16908) );
  INV_X1 U10731 ( .A(n16908), .ZN(n16909) );
  BUF_X1 U10732 ( .A(n16914), .Z(n16910) );
  INV_X1 U10733 ( .A(n273900), .ZN(n16911) );
  INV_X1 U10734 ( .A(n16911), .ZN(n16912) );
  INV_X1 U10735 ( .A(n6254), .ZN(n16913) );
  INV_X1 U10736 ( .A(n16913), .ZN(n16914) );
  BUF_X1 U10737 ( .A(n16919), .Z(n16915) );
  INV_X1 U10738 ( .A(n274200), .ZN(n16916) );
  INV_X1 U10739 ( .A(n16916), .ZN(n16917) );
  INV_X1 U10740 ( .A(n6257), .ZN(n16918) );
  INV_X1 U10741 ( .A(n16918), .ZN(n16919) );
  BUF_X1 U10742 ( .A(n16924), .Z(n16920) );
  INV_X1 U10743 ( .A(n28530), .ZN(n16921) );
  INV_X1 U10744 ( .A(n16921), .ZN(n16922) );
  INV_X1 U10745 ( .A(n63560), .ZN(n16923) );
  INV_X1 U10746 ( .A(n16923), .ZN(n16924) );
  BUF_X1 U10747 ( .A(n16929), .Z(n16925) );
  INV_X1 U10748 ( .A(n2749), .ZN(n16926) );
  INV_X1 U10749 ( .A(n16926), .ZN(n16927) );
  INV_X1 U10750 ( .A(n62640), .ZN(n16928) );
  INV_X1 U10751 ( .A(n16928), .ZN(n16929) );
  BUF_X1 U10752 ( .A(n16934), .Z(n16930) );
  INV_X1 U10753 ( .A(n28660), .ZN(n16931) );
  INV_X1 U10754 ( .A(n16931), .ZN(n16932) );
  INV_X1 U10755 ( .A(n63690), .ZN(n16933) );
  INV_X1 U10756 ( .A(n16933), .ZN(n16934) );
  BUF_X1 U10757 ( .A(n16939), .Z(n16935) );
  INV_X1 U10758 ( .A(n273800), .ZN(n16936) );
  INV_X1 U10759 ( .A(n16936), .ZN(n16937) );
  INV_X1 U10760 ( .A(n6253), .ZN(n16938) );
  INV_X1 U10761 ( .A(n16938), .ZN(n16939) );
  BUF_X1 U10762 ( .A(n16944), .Z(n16940) );
  INV_X1 U10763 ( .A(n28640), .ZN(n16941) );
  INV_X1 U10764 ( .A(n16941), .ZN(n16942) );
  INV_X1 U10765 ( .A(n63670), .ZN(n16943) );
  INV_X1 U10766 ( .A(n16943), .ZN(n16944) );
  BUF_X1 U10767 ( .A(n16949), .Z(n16945) );
  INV_X1 U10768 ( .A(n28590), .ZN(n16946) );
  INV_X1 U10769 ( .A(n16946), .ZN(n16947) );
  INV_X1 U10770 ( .A(n63620), .ZN(n16948) );
  INV_X1 U10771 ( .A(n16948), .ZN(n16949) );
  BUF_X1 U10772 ( .A(n16954), .Z(n16950) );
  INV_X1 U10773 ( .A(n274100), .ZN(n16951) );
  INV_X1 U10774 ( .A(n16951), .ZN(n16952) );
  INV_X1 U10775 ( .A(n6256), .ZN(n16953) );
  INV_X1 U10776 ( .A(n16953), .ZN(n16954) );
  BUF_X1 U10777 ( .A(n16958), .Z(n16955) );
  INV_X1 U10778 ( .A(matrix_mul_2D_7__6__0_), .ZN(n16956) );
  INV_X1 U10779 ( .A(n63700), .ZN(n16957) );
  INV_X1 U10780 ( .A(n16957), .ZN(n16958) );
  BUF_X1 U10781 ( .A(n16963), .Z(n16959) );
  INV_X1 U10782 ( .A(n28630), .ZN(n16960) );
  INV_X1 U10783 ( .A(n16960), .ZN(n16961) );
  INV_X1 U10784 ( .A(n63660), .ZN(n16962) );
  INV_X1 U10785 ( .A(n16962), .ZN(n16963) );
  BUF_X1 U10786 ( .A(n16968), .Z(n16964) );
  INV_X1 U10787 ( .A(n274300), .ZN(n16965) );
  INV_X1 U10788 ( .A(n16965), .ZN(n16966) );
  INV_X1 U10789 ( .A(n6258), .ZN(n16967) );
  INV_X1 U10790 ( .A(n16967), .ZN(n16968) );
  BUF_X1 U10791 ( .A(n16973), .Z(n16969) );
  INV_X1 U10792 ( .A(n273600), .ZN(n16970) );
  INV_X1 U10793 ( .A(n16970), .ZN(n16971) );
  INV_X1 U10794 ( .A(n6251), .ZN(n16972) );
  INV_X1 U10795 ( .A(n16972), .ZN(n16973) );
  BUF_X1 U10796 ( .A(n16978), .Z(n16974) );
  INV_X1 U10797 ( .A(n274400), .ZN(n16975) );
  INV_X1 U10798 ( .A(n16975), .ZN(n16976) );
  INV_X1 U10799 ( .A(n6259), .ZN(n16977) );
  INV_X1 U10800 ( .A(n16977), .ZN(n16978) );
  BUF_X1 U10801 ( .A(n16983), .Z(n16979) );
  INV_X1 U10802 ( .A(n274600), .ZN(n16980) );
  INV_X1 U10803 ( .A(n16980), .ZN(n16981) );
  INV_X1 U10804 ( .A(n62610), .ZN(n16982) );
  INV_X1 U10805 ( .A(n16982), .ZN(n16983) );
  BUF_X1 U10806 ( .A(n16988), .Z(n16984) );
  INV_X1 U10807 ( .A(n28570), .ZN(n16985) );
  INV_X1 U10808 ( .A(n16985), .ZN(n16986) );
  INV_X1 U10809 ( .A(n63600), .ZN(n16987) );
  INV_X1 U10810 ( .A(n16987), .ZN(n16988) );
  BUF_X1 U10811 ( .A(n16993), .Z(n16989) );
  INV_X1 U10812 ( .A(n28540), .ZN(n16990) );
  INV_X1 U10813 ( .A(n16990), .ZN(n16991) );
  INV_X1 U10814 ( .A(n63570), .ZN(n16992) );
  INV_X1 U10815 ( .A(n16992), .ZN(n16993) );
  BUF_X1 U10816 ( .A(n16998), .Z(n16994) );
  INV_X1 U10817 ( .A(n28560), .ZN(n16995) );
  INV_X1 U10818 ( .A(n16995), .ZN(n16996) );
  INV_X1 U10819 ( .A(n63590), .ZN(n16997) );
  INV_X1 U10820 ( .A(n16997), .ZN(n16998) );
  BUF_X1 U10821 ( .A(n17003), .Z(n16999) );
  INV_X1 U10822 ( .A(n274000), .ZN(n17000) );
  INV_X1 U10823 ( .A(n17000), .ZN(n17001) );
  INV_X1 U10824 ( .A(n6255), .ZN(n17002) );
  INV_X1 U10825 ( .A(n17002), .ZN(n17003) );
  BUF_X1 U10826 ( .A(n17008), .Z(n17004) );
  INV_X1 U10827 ( .A(n28550), .ZN(n17005) );
  INV_X1 U10828 ( .A(n17005), .ZN(n17006) );
  INV_X1 U10829 ( .A(n63580), .ZN(n17007) );
  INV_X1 U10830 ( .A(n17007), .ZN(n17008) );
  BUF_X1 U10831 ( .A(n17013), .Z(n17009) );
  INV_X1 U10832 ( .A(n2870), .ZN(n17010) );
  INV_X1 U10833 ( .A(n17010), .ZN(n17011) );
  INV_X1 U10834 ( .A(n6373), .ZN(n17012) );
  INV_X1 U10835 ( .A(n17012), .ZN(n17013) );
  BUF_X1 U10836 ( .A(n17017), .Z(n17014) );
  INV_X1 U10837 ( .A(matrix_mul_2D_7__7__0_), .ZN(n17015) );
  INV_X1 U10838 ( .A(n6385), .ZN(n17016) );
  INV_X1 U10839 ( .A(n17016), .ZN(n17017) );
  BUF_X1 U10840 ( .A(n17022), .Z(n17018) );
  INV_X1 U10841 ( .A(n28680), .ZN(n17019) );
  INV_X1 U10842 ( .A(n17019), .ZN(n17020) );
  INV_X1 U10843 ( .A(n6371), .ZN(n17021) );
  INV_X1 U10844 ( .A(n17021), .ZN(n17022) );
  BUF_X1 U10845 ( .A(n17027), .Z(n17023) );
  INV_X1 U10846 ( .A(n2869), .ZN(n17024) );
  INV_X1 U10847 ( .A(n17024), .ZN(n17025) );
  INV_X1 U10848 ( .A(n6372), .ZN(n17026) );
  INV_X1 U10849 ( .A(n17026), .ZN(n17027) );
  BUF_X1 U10850 ( .A(n17032), .Z(n17028) );
  INV_X1 U10851 ( .A(n2879), .ZN(n17029) );
  INV_X1 U10852 ( .A(n17029), .ZN(n17030) );
  INV_X1 U10853 ( .A(n6382), .ZN(n17031) );
  INV_X1 U10854 ( .A(n17031), .ZN(n17032) );
  BUF_X1 U10855 ( .A(n17037), .Z(n17033) );
  INV_X1 U10856 ( .A(n2880), .ZN(n17034) );
  INV_X1 U10857 ( .A(n17034), .ZN(n17035) );
  INV_X1 U10858 ( .A(n6383), .ZN(n17036) );
  INV_X1 U10859 ( .A(n17036), .ZN(n17037) );
  BUF_X1 U10860 ( .A(n17042), .Z(n17038) );
  INV_X1 U10861 ( .A(n2881), .ZN(n17039) );
  INV_X1 U10862 ( .A(n17039), .ZN(n17040) );
  INV_X1 U10863 ( .A(n6384), .ZN(n17041) );
  INV_X1 U10864 ( .A(n17041), .ZN(n17042) );
  BUF_X1 U10865 ( .A(n17047), .Z(n17043) );
  INV_X1 U10866 ( .A(n2876), .ZN(n17044) );
  INV_X1 U10867 ( .A(n17044), .ZN(n17045) );
  INV_X1 U10868 ( .A(n6379), .ZN(n17046) );
  INV_X1 U10869 ( .A(n17046), .ZN(n17047) );
  BUF_X1 U10870 ( .A(n17052), .Z(n17048) );
  INV_X1 U10871 ( .A(n2877), .ZN(n17049) );
  INV_X1 U10872 ( .A(n17049), .ZN(n17050) );
  INV_X1 U10873 ( .A(n6380), .ZN(n17051) );
  INV_X1 U10874 ( .A(n17051), .ZN(n17052) );
  BUF_X1 U10875 ( .A(n17057), .Z(n17053) );
  INV_X1 U10876 ( .A(n2878), .ZN(n17054) );
  INV_X1 U10877 ( .A(n17054), .ZN(n17055) );
  INV_X1 U10878 ( .A(n6381), .ZN(n17056) );
  INV_X1 U10879 ( .A(n17056), .ZN(n17057) );
  BUF_X1 U10880 ( .A(n17062), .Z(n17058) );
  INV_X1 U10881 ( .A(n2874), .ZN(n17059) );
  INV_X1 U10882 ( .A(n17059), .ZN(n17060) );
  INV_X1 U10883 ( .A(n6377), .ZN(n17061) );
  INV_X1 U10884 ( .A(n17061), .ZN(n17062) );
  BUF_X1 U10885 ( .A(n17067), .Z(n17063) );
  INV_X1 U10886 ( .A(n2875), .ZN(n17064) );
  INV_X1 U10887 ( .A(n17064), .ZN(n17065) );
  INV_X1 U10888 ( .A(n6378), .ZN(n17066) );
  INV_X1 U10889 ( .A(n17066), .ZN(n17067) );
  CLKBUF_X1 U10890 ( .A(n22694), .Z(n17068) );
  CLKBUF_X1 U10891 ( .A(r899_B_7_), .Z(n17069) );
  CLKBUF_X1 U10892 ( .A(n17071), .Z(n17070) );
  CLKBUF_X1 U10893 ( .A(n23937), .Z(n17071) );
  NAND2_X1 U10894 ( .A1(n26637), .A2(n27298), .ZN(n17072) );
  CLKBUF_X1 U10895 ( .A(n23650), .Z(n17073) );
  CLKBUF_X1 U10896 ( .A(n18611), .Z(n17074) );
  CLKBUF_X1 U10897 ( .A(n18610), .Z(n17075) );
  CLKBUF_X1 U10898 ( .A(n18595), .Z(n17076) );
  CLKBUF_X1 U10899 ( .A(n18593), .Z(n17077) );
  CLKBUF_X1 U10900 ( .A(n18984), .Z(n17078) );
  CLKBUF_X1 U10901 ( .A(n18566), .Z(n17079) );
  CLKBUF_X1 U10902 ( .A(n18559), .Z(n17080) );
  CLKBUF_X1 U10903 ( .A(n23014), .Z(n17081) );
  CLKBUF_X1 U10904 ( .A(n3186), .Z(n17082) );
  CLKBUF_X1 U10905 ( .A(n54220), .Z(n17083) );
  CLKBUF_X1 U10906 ( .A(n18162), .Z(n17084) );
  CLKBUF_X1 U10907 ( .A(n27293), .Z(n17085) );
  CLKBUF_X1 U10908 ( .A(n54240), .Z(n17086) );
  CLKBUF_X1 U10909 ( .A(n24101), .Z(n17087) );
  CLKBUF_X1 U10910 ( .A(n22752), .Z(n17088) );
  CLKBUF_X1 U10911 ( .A(n26688), .Z(n17089) );
  CLKBUF_X1 U10912 ( .A(n22766), .Z(n17090) );
  CLKBUF_X1 U10913 ( .A(n20644), .Z(n17091) );
  CLKBUF_X1 U10914 ( .A(n20635), .Z(n17092) );
  CLKBUF_X1 U10915 ( .A(n20634), .Z(n17093) );
  CLKBUF_X1 U10916 ( .A(n20626), .Z(n17094) );
  CLKBUF_X1 U10917 ( .A(n27148), .Z(n17095) );
  CLKBUF_X1 U10918 ( .A(n27270), .Z(n17096) );
  CLKBUF_X1 U10919 ( .A(n27219), .Z(n17097) );
  CLKBUF_X1 U10920 ( .A(n20535), .Z(n17098) );
  CLKBUF_X1 U10921 ( .A(n20906), .Z(n17099) );
  CLKBUF_X1 U10922 ( .A(n20901), .Z(n17100) );
  CLKBUF_X1 U10923 ( .A(n20538), .Z(n17101) );
  CLKBUF_X1 U10924 ( .A(n5200), .Z(n17102) );
  CLKBUF_X1 U10925 ( .A(n22879), .Z(n17103) );
  CLKBUF_X1 U10926 ( .A(n24649), .Z(n17104) );
  CLKBUF_X1 U10927 ( .A(n17068), .Z(n17105) );
  CLKBUF_X1 U10928 ( .A(n26897), .Z(n17106) );
  CLKBUF_X1 U10929 ( .A(n26895), .Z(n17107) );
  CLKBUF_X1 U10930 ( .A(n26899), .Z(n17108) );
  CLKBUF_X1 U10931 ( .A(n26898), .Z(n17109) );
  CLKBUF_X1 U10932 ( .A(n22711), .Z(n17110) );
  CLKBUF_X1 U10933 ( .A(n20785), .Z(n17111) );
  CLKBUF_X1 U10934 ( .A(n21864), .Z(n17112) );
  CLKBUF_X1 U10935 ( .A(n17124), .Z(n17113) );
  CLKBUF_X1 U10936 ( .A(n26514), .Z(n17114) );
  CLKBUF_X1 U10937 ( .A(n23644), .Z(n17115) );
  CLKBUF_X1 U10938 ( .A(n26497), .Z(n17116) );
  CLKBUF_X1 U10939 ( .A(n26379), .Z(n17117) );
  CLKBUF_X1 U10940 ( .A(n26323), .Z(n17118) );
  CLKBUF_X1 U10941 ( .A(n25918), .Z(n17119) );
  CLKBUF_X1 U10942 ( .A(n26727), .Z(n17120) );
  CLKBUF_X1 U10943 ( .A(n25517), .Z(n17121) );
  CLKBUF_X1 U10944 ( .A(n25513), .Z(n17122) );
  CLKBUF_X1 U10945 ( .A(n25245), .Z(n17123) );
  NAND3_X1 U10946 ( .A1(n21438), .A2(n25662), .A3(n17083), .ZN(n17124) );
  INV_X1 U10947 ( .A(n25942), .ZN(n17125) );
  INV_X1 U10948 ( .A(n17125), .ZN(n17126) );
  INV_X1 U10949 ( .A(n17125), .ZN(n17127) );
  INV_X1 U10950 ( .A(n17124), .ZN(n17128) );
  NAND4_X1 U10951 ( .A1(n17086), .A2(n24714), .A3(n24711), .A4(n19755), .ZN(
        n17129) );
  CLKBUF_X1 U10952 ( .A(n27333), .Z(n17130) );
  NAND3_X1 U10953 ( .A1(n22432), .A2(n3097), .A3(n22468), .ZN(n17131) );
  INV_X1 U10954 ( .A(n17131), .ZN(n17132) );
  INV_X1 U10955 ( .A(n17131), .ZN(n17133) );
  INV_X1 U10956 ( .A(n17129), .ZN(n17134) );
  INV_X1 U10957 ( .A(n17129), .ZN(n17135) );
  CLKBUF_X1 U10958 ( .A(n18985), .Z(n17136) );
  CLKBUF_X1 U10959 ( .A(n42090), .Z(n17265) );
  CLKBUF_X1 U10960 ( .A(n45660), .Z(n17266) );
  NOR4_X1 U10961 ( .A1(n542), .A2(n553), .A3(n17996), .A4(n4570), .ZN(n17267)
         );
  CLKBUF_X1 U10962 ( .A(n26987), .Z(n17268) );
  NAND3_X1 U10963 ( .A1(n877), .A2(n25957), .A3(n19109), .ZN(n17269) );
  INV_X1 U10964 ( .A(n17270), .ZN(n17271) );
  INV_X1 U10965 ( .A(n17272), .ZN(n17273) );
  INV_X1 U10966 ( .A(n17274), .ZN(n17275) );
  INV_X1 U10967 ( .A(n17276), .ZN(n17277) );
  INV_X1 U10968 ( .A(n17278), .ZN(n17279) );
  INV_X1 U10969 ( .A(n17280), .ZN(n17281) );
  INV_X1 U10970 ( .A(n17282), .ZN(n17283) );
  INV_X1 U10971 ( .A(n17284), .ZN(n17285) );
  INV_X1 U10972 ( .A(n17286), .ZN(n17287) );
  INV_X1 U10973 ( .A(n17288), .ZN(n17289) );
  INV_X1 U10974 ( .A(n17290), .ZN(n17291) );
  INV_X1 U10975 ( .A(n17292), .ZN(n17293) );
  INV_X1 U10976 ( .A(n17294), .ZN(n17295) );
  INV_X1 U10977 ( .A(n17296), .ZN(n17297) );
  INV_X1 U10978 ( .A(n17298), .ZN(n17299) );
  INV_X1 U10979 ( .A(n17300), .ZN(n17301) );
  INV_X1 U10980 ( .A(n17302), .ZN(n17303) );
  INV_X1 U10981 ( .A(n17304), .ZN(n17305) );
  INV_X1 U10982 ( .A(n17306), .ZN(n17307) );
  INV_X1 U10983 ( .A(n17308), .ZN(n17309) );
  INV_X1 U10984 ( .A(n17310), .ZN(n17311) );
  INV_X1 U10985 ( .A(n17312), .ZN(n17313) );
  INV_X1 U10986 ( .A(n17314), .ZN(n17315) );
  INV_X1 U10987 ( .A(n17316), .ZN(n17317) );
  INV_X1 U10988 ( .A(n17318), .ZN(n17319) );
  INV_X1 U10989 ( .A(n17320), .ZN(n17321) );
  INV_X1 U10990 ( .A(n17322), .ZN(n17323) );
  INV_X1 U10991 ( .A(n17324), .ZN(n17325) );
  INV_X1 U10992 ( .A(n17326), .ZN(n17327) );
  INV_X1 U10993 ( .A(n17328), .ZN(n17329) );
  INV_X1 U10994 ( .A(n17330), .ZN(n17331) );
  INV_X1 U10995 ( .A(n17332), .ZN(n17333) );
  INV_X1 U10996 ( .A(n17334), .ZN(n17335) );
  INV_X1 U10997 ( .A(n17336), .ZN(n17337) );
  INV_X1 U10998 ( .A(n17338), .ZN(n17339) );
  INV_X1 U10999 ( .A(n17340), .ZN(n17341) );
  INV_X1 U11000 ( .A(n17342), .ZN(n17343) );
  INV_X1 U11001 ( .A(n17344), .ZN(n17345) );
  INV_X1 U11002 ( .A(n17346), .ZN(n17347) );
  INV_X1 U11003 ( .A(n17348), .ZN(n17349) );
  INV_X1 U11004 ( .A(n17350), .ZN(n17351) );
  INV_X1 U11005 ( .A(n17352), .ZN(n17353) );
  INV_X1 U11006 ( .A(n17354), .ZN(n17355) );
  INV_X1 U11007 ( .A(n17356), .ZN(n17357) );
  INV_X1 U11008 ( .A(n17358), .ZN(n17359) );
  INV_X1 U11009 ( .A(n17360), .ZN(n17361) );
  INV_X1 U11010 ( .A(n17362), .ZN(n17363) );
  INV_X1 U11011 ( .A(n17364), .ZN(n17365) );
  INV_X1 U11012 ( .A(n17366), .ZN(n17367) );
  INV_X1 U11013 ( .A(n17368), .ZN(n17369) );
  INV_X1 U11014 ( .A(n17370), .ZN(n17371) );
  INV_X1 U11015 ( .A(n17372), .ZN(n17373) );
  INV_X1 U11016 ( .A(n17374), .ZN(n17375) );
  INV_X1 U11017 ( .A(n17376), .ZN(n17377) );
  INV_X1 U11018 ( .A(n17378), .ZN(n17379) );
  INV_X1 U11019 ( .A(n17380), .ZN(n17381) );
  INV_X1 U11020 ( .A(n17382), .ZN(n17383) );
  INV_X1 U11021 ( .A(n17384), .ZN(n17385) );
  INV_X1 U11022 ( .A(n17386), .ZN(n17387) );
  INV_X1 U11023 ( .A(n17388), .ZN(n17389) );
  INV_X1 U11024 ( .A(n17390), .ZN(n17391) );
  INV_X1 U11025 ( .A(n17392), .ZN(n17393) );
  INV_X1 U11026 ( .A(n17394), .ZN(n17395) );
  INV_X1 U11027 ( .A(n17396), .ZN(n17397) );
  INV_X1 U11028 ( .A(n17398), .ZN(n17399) );
  INV_X1 U11029 ( .A(n17400), .ZN(n17401) );
  INV_X1 U11030 ( .A(n17402), .ZN(n17403) );
  INV_X1 U11031 ( .A(n17404), .ZN(n17405) );
  INV_X1 U11032 ( .A(n17406), .ZN(n17407) );
  INV_X1 U11033 ( .A(n17408), .ZN(n17409) );
  INV_X1 U11034 ( .A(n17410), .ZN(n17411) );
  INV_X1 U11035 ( .A(n17412), .ZN(n17413) );
  INV_X1 U11036 ( .A(n17414), .ZN(n17415) );
  INV_X1 U11037 ( .A(n17416), .ZN(n17417) );
  INV_X1 U11038 ( .A(n17418), .ZN(n17419) );
  INV_X1 U11039 ( .A(n17420), .ZN(n17421) );
  INV_X1 U11040 ( .A(n17422), .ZN(n17423) );
  INV_X1 U11041 ( .A(n17424), .ZN(n17425) );
  INV_X1 U11042 ( .A(n17426), .ZN(n17427) );
  INV_X1 U11043 ( .A(n17428), .ZN(n17429) );
  INV_X1 U11044 ( .A(n17430), .ZN(n17431) );
  INV_X1 U11045 ( .A(n17432), .ZN(n17433) );
  INV_X1 U11046 ( .A(n17434), .ZN(n17435) );
  INV_X1 U11047 ( .A(n17436), .ZN(n17437) );
  INV_X1 U11048 ( .A(n17438), .ZN(n17439) );
  INV_X1 U11049 ( .A(n17440), .ZN(n17441) );
  INV_X1 U11050 ( .A(n17442), .ZN(n17443) );
  INV_X1 U11051 ( .A(n17444), .ZN(n17445) );
  INV_X1 U11052 ( .A(n17446), .ZN(n17447) );
  INV_X1 U11053 ( .A(n17448), .ZN(n17449) );
  INV_X1 U11054 ( .A(n17450), .ZN(n17451) );
  INV_X1 U11055 ( .A(n17452), .ZN(n17453) );
  INV_X1 U11056 ( .A(n17454), .ZN(n17455) );
  INV_X1 U11057 ( .A(n17456), .ZN(n17457) );
  INV_X1 U11058 ( .A(n17458), .ZN(n17459) );
  INV_X1 U11059 ( .A(n17460), .ZN(n17461) );
  INV_X1 U11060 ( .A(n17462), .ZN(n17463) );
  INV_X1 U11061 ( .A(n17464), .ZN(n17465) );
  INV_X1 U11062 ( .A(n17466), .ZN(n17467) );
  INV_X1 U11063 ( .A(n17468), .ZN(n17469) );
  INV_X1 U11064 ( .A(n17470), .ZN(n17471) );
  INV_X1 U11065 ( .A(n17472), .ZN(n17473) );
  INV_X1 U11066 ( .A(n17474), .ZN(n17475) );
  INV_X1 U11067 ( .A(n17476), .ZN(n17477) );
  INV_X1 U11068 ( .A(n17478), .ZN(n17479) );
  INV_X1 U11069 ( .A(n17480), .ZN(n17481) );
  INV_X1 U11070 ( .A(n17482), .ZN(n17483) );
  INV_X1 U11071 ( .A(n17484), .ZN(n17485) );
  INV_X1 U11072 ( .A(n17486), .ZN(n17487) );
  INV_X1 U11073 ( .A(n17488), .ZN(n17489) );
  INV_X1 U11074 ( .A(n17490), .ZN(n17491) );
  INV_X1 U11075 ( .A(n17492), .ZN(n17493) );
  INV_X1 U11076 ( .A(n17494), .ZN(n17495) );
  INV_X1 U11077 ( .A(n17496), .ZN(n17497) );
  INV_X1 U11078 ( .A(n17498), .ZN(n17499) );
  INV_X1 U11079 ( .A(n17500), .ZN(n17501) );
  INV_X1 U11080 ( .A(n17502), .ZN(n17503) );
  INV_X1 U11081 ( .A(n17504), .ZN(n17505) );
  INV_X1 U11082 ( .A(n17506), .ZN(n17507) );
  INV_X1 U11083 ( .A(n17508), .ZN(n17509) );
  INV_X1 U11084 ( .A(n17510), .ZN(n17511) );
  INV_X1 U11085 ( .A(n17512), .ZN(n17513) );
  INV_X1 U11086 ( .A(n17514), .ZN(n17515) );
  INV_X1 U11087 ( .A(n17516), .ZN(n17517) );
  INV_X1 U11088 ( .A(n17518), .ZN(n17519) );
  INV_X1 U11089 ( .A(n17520), .ZN(n17521) );
  INV_X1 U11090 ( .A(n17522), .ZN(n17523) );
  INV_X1 U11091 ( .A(n17524), .ZN(n17525) );
  INV_X1 U11092 ( .A(n17526), .ZN(n17527) );
  INV_X1 U11093 ( .A(n17528), .ZN(n17529) );
  INV_X1 U11094 ( .A(n17530), .ZN(n17531) );
  INV_X1 U11095 ( .A(n17532), .ZN(n17533) );
  INV_X1 U11096 ( .A(n17534), .ZN(n17535) );
  INV_X1 U11097 ( .A(n17536), .ZN(n17537) );
  INV_X1 U11098 ( .A(n17538), .ZN(n17539) );
  INV_X1 U11099 ( .A(n17540), .ZN(n17541) );
  INV_X1 U11100 ( .A(n17542), .ZN(n17543) );
  INV_X1 U11101 ( .A(n17544), .ZN(n17545) );
  INV_X1 U11102 ( .A(n17546), .ZN(n17547) );
  INV_X1 U11103 ( .A(n17548), .ZN(n17549) );
  INV_X1 U11104 ( .A(n17550), .ZN(n17551) );
  INV_X1 U11105 ( .A(n17552), .ZN(n17553) );
  INV_X1 U11106 ( .A(n17554), .ZN(n17555) );
  INV_X1 U11107 ( .A(n17556), .ZN(n17557) );
  INV_X1 U11108 ( .A(n17558), .ZN(n17559) );
  INV_X1 U11109 ( .A(n17560), .ZN(n17561) );
  INV_X1 U11110 ( .A(n17562), .ZN(n17563) );
  INV_X1 U11111 ( .A(n17564), .ZN(n17565) );
  INV_X1 U11112 ( .A(n17566), .ZN(n17567) );
  INV_X1 U11113 ( .A(n17568), .ZN(n17569) );
  INV_X1 U11114 ( .A(n17570), .ZN(n17571) );
  INV_X1 U11115 ( .A(n17572), .ZN(n17573) );
  INV_X1 U11116 ( .A(n17574), .ZN(n17575) );
  INV_X1 U11117 ( .A(n17576), .ZN(n17577) );
  INV_X1 U11118 ( .A(n17578), .ZN(n17579) );
  INV_X1 U11119 ( .A(n17580), .ZN(n17581) );
  INV_X1 U11120 ( .A(n17582), .ZN(n17583) );
  INV_X1 U11121 ( .A(n17584), .ZN(n17585) );
  INV_X1 U11122 ( .A(n17586), .ZN(n17587) );
  INV_X1 U11123 ( .A(n17588), .ZN(n17589) );
  INV_X1 U11124 ( .A(n17590), .ZN(n17591) );
  INV_X1 U11125 ( .A(n17592), .ZN(n17593) );
  INV_X1 U11126 ( .A(n17594), .ZN(n17595) );
  INV_X1 U11127 ( .A(n17596), .ZN(n17597) );
  INV_X1 U11128 ( .A(n17598), .ZN(n17599) );
  INV_X1 U11129 ( .A(n17600), .ZN(n17601) );
  INV_X1 U11130 ( .A(n17602), .ZN(n17603) );
  INV_X1 U11131 ( .A(n17604), .ZN(n17605) );
  INV_X1 U11132 ( .A(n17606), .ZN(n17607) );
  INV_X1 U11133 ( .A(n17608), .ZN(n17609) );
  INV_X1 U11134 ( .A(n17610), .ZN(n17611) );
  INV_X1 U11135 ( .A(n17612), .ZN(n17613) );
  INV_X1 U11136 ( .A(n17614), .ZN(n17615) );
  INV_X1 U11137 ( .A(n17616), .ZN(n17617) );
  INV_X1 U11138 ( .A(n17618), .ZN(n17619) );
  INV_X1 U11139 ( .A(n17620), .ZN(n17621) );
  INV_X1 U11140 ( .A(n17622), .ZN(n17623) );
  INV_X1 U11141 ( .A(n17624), .ZN(n17625) );
  INV_X1 U11142 ( .A(n17626), .ZN(n17627) );
  INV_X1 U11143 ( .A(n17628), .ZN(n17629) );
  INV_X1 U11144 ( .A(n17630), .ZN(n17631) );
  INV_X1 U11145 ( .A(n17632), .ZN(n17633) );
  INV_X1 U11146 ( .A(n17634), .ZN(n17635) );
  INV_X1 U11147 ( .A(n17636), .ZN(n17637) );
  INV_X1 U11148 ( .A(n17638), .ZN(n17639) );
  INV_X1 U11149 ( .A(n17640), .ZN(n17641) );
  INV_X1 U11150 ( .A(n17642), .ZN(n17643) );
  INV_X1 U11151 ( .A(n17644), .ZN(n17645) );
  INV_X1 U11152 ( .A(n17646), .ZN(n17647) );
  INV_X1 U11153 ( .A(n17648), .ZN(n17649) );
  INV_X1 U11154 ( .A(n17650), .ZN(n17651) );
  INV_X1 U11155 ( .A(n17652), .ZN(n17653) );
  INV_X1 U11156 ( .A(n17654), .ZN(n17655) );
  INV_X1 U11157 ( .A(n17656), .ZN(n17657) );
  INV_X1 U11158 ( .A(n17658), .ZN(n17659) );
  INV_X1 U11159 ( .A(n17660), .ZN(n17661) );
  INV_X1 U11160 ( .A(n17662), .ZN(n17663) );
  INV_X1 U11161 ( .A(n17664), .ZN(n17665) );
  INV_X1 U11162 ( .A(n17666), .ZN(n17667) );
  INV_X1 U11163 ( .A(n17668), .ZN(n17669) );
  INV_X1 U11164 ( .A(n17670), .ZN(n17671) );
  INV_X1 U11165 ( .A(n17672), .ZN(n17673) );
  INV_X1 U11166 ( .A(n17674), .ZN(n17675) );
  INV_X1 U11167 ( .A(n17676), .ZN(n17677) );
  INV_X1 U11168 ( .A(n17678), .ZN(n17679) );
  INV_X1 U11169 ( .A(n17680), .ZN(n17681) );
  INV_X1 U11170 ( .A(n17682), .ZN(n17683) );
  INV_X1 U11171 ( .A(n17684), .ZN(n17685) );
  INV_X1 U11172 ( .A(n17686), .ZN(n17687) );
  INV_X1 U11173 ( .A(n17688), .ZN(n17689) );
  INV_X1 U11174 ( .A(n17690), .ZN(n17691) );
  INV_X1 U11175 ( .A(n17692), .ZN(n17693) );
  INV_X1 U11176 ( .A(n17694), .ZN(n17695) );
  INV_X1 U11177 ( .A(n17696), .ZN(n17697) );
  INV_X1 U11178 ( .A(n17698), .ZN(n17699) );
  INV_X1 U11179 ( .A(n17700), .ZN(n17701) );
  INV_X1 U11180 ( .A(n17702), .ZN(n17703) );
  INV_X1 U11181 ( .A(n17704), .ZN(n17705) );
  INV_X1 U11182 ( .A(n17706), .ZN(n17707) );
  INV_X1 U11183 ( .A(n17708), .ZN(n17709) );
  INV_X1 U11184 ( .A(n17710), .ZN(n17711) );
  INV_X1 U11185 ( .A(n17712), .ZN(n17713) );
  INV_X1 U11186 ( .A(n17714), .ZN(n17715) );
  INV_X1 U11187 ( .A(n17716), .ZN(n17717) );
  INV_X1 U11188 ( .A(n17718), .ZN(n17719) );
  INV_X1 U11189 ( .A(n17720), .ZN(n17721) );
  INV_X1 U11190 ( .A(n17722), .ZN(n17723) );
  INV_X1 U11191 ( .A(n17724), .ZN(n17725) );
  INV_X1 U11192 ( .A(n17726), .ZN(n17727) );
  INV_X1 U11193 ( .A(n17728), .ZN(n17729) );
  INV_X1 U11194 ( .A(n17730), .ZN(n17731) );
  INV_X1 U11195 ( .A(n17732), .ZN(n17733) );
  INV_X1 U11196 ( .A(n17734), .ZN(n17735) );
  INV_X1 U11197 ( .A(n17736), .ZN(n17737) );
  INV_X1 U11198 ( .A(n17738), .ZN(n17739) );
  INV_X1 U11199 ( .A(n17740), .ZN(n17741) );
  INV_X1 U11200 ( .A(n17742), .ZN(n17743) );
  INV_X1 U11201 ( .A(n17744), .ZN(n17745) );
  INV_X1 U11202 ( .A(n17746), .ZN(n17747) );
  INV_X1 U11203 ( .A(n17748), .ZN(n17749) );
  INV_X1 U11204 ( .A(n17750), .ZN(n17751) );
  INV_X1 U11205 ( .A(n17752), .ZN(n17753) );
  INV_X1 U11206 ( .A(n17754), .ZN(n17755) );
  INV_X1 U11207 ( .A(n17756), .ZN(n17757) );
  INV_X1 U11208 ( .A(n17758), .ZN(n17759) );
  INV_X1 U11209 ( .A(n17760), .ZN(n17761) );
  INV_X1 U11210 ( .A(n17762), .ZN(n17763) );
  INV_X1 U11211 ( .A(n17764), .ZN(n17765) );
  INV_X1 U11212 ( .A(n17766), .ZN(n17767) );
  INV_X1 U11213 ( .A(n17768), .ZN(n17769) );
  INV_X1 U11214 ( .A(n17770), .ZN(n17771) );
  INV_X1 U11215 ( .A(n17772), .ZN(n17773) );
  INV_X1 U11216 ( .A(n17774), .ZN(n17775) );
  INV_X1 U11217 ( .A(n17776), .ZN(n17777) );
  INV_X1 U11218 ( .A(n17778), .ZN(n17779) );
  INV_X1 U11219 ( .A(n17780), .ZN(n17781) );
  INV_X1 U11220 ( .A(n17782), .ZN(n17783) );
  INV_X1 U11221 ( .A(n17784), .ZN(n17785) );
  INV_X1 U11222 ( .A(n17786), .ZN(n17787) );
  INV_X1 U11223 ( .A(n17788), .ZN(n17789) );
  INV_X1 U11224 ( .A(n17790), .ZN(n17791) );
  INV_X1 U11225 ( .A(n17792), .ZN(n17793) );
  INV_X1 U11226 ( .A(n17794), .ZN(n17795) );
  INV_X1 U11227 ( .A(n17796), .ZN(n17797) );
  INV_X1 U11228 ( .A(n17798), .ZN(n17799) );
  INV_X1 U11229 ( .A(n17800), .ZN(n17801) );
  INV_X1 U11230 ( .A(n17802), .ZN(n17803) );
  INV_X1 U11231 ( .A(n17804), .ZN(n17805) );
  INV_X1 U11232 ( .A(n17806), .ZN(n17807) );
  INV_X1 U11233 ( .A(n17808), .ZN(n17809) );
  INV_X1 U11234 ( .A(n17810), .ZN(n17811) );
  INV_X1 U11235 ( .A(n17812), .ZN(n17813) );
  INV_X1 U11236 ( .A(n17814), .ZN(n17815) );
  INV_X1 U11237 ( .A(n17816), .ZN(n17817) );
  INV_X1 U11238 ( .A(n17818), .ZN(n17819) );
  INV_X1 U11239 ( .A(n17820), .ZN(n17821) );
  INV_X1 U11240 ( .A(n17822), .ZN(n17823) );
  INV_X1 U11241 ( .A(n17824), .ZN(n17825) );
  INV_X1 U11242 ( .A(n17826), .ZN(n17827) );
  INV_X1 U11243 ( .A(n17828), .ZN(n17829) );
  INV_X1 U11244 ( .A(n17830), .ZN(n17831) );
  INV_X1 U11245 ( .A(n17832), .ZN(n17833) );
  INV_X1 U11246 ( .A(n17834), .ZN(n17835) );
  INV_X1 U11247 ( .A(n17836), .ZN(n17837) );
  INV_X1 U11248 ( .A(n17838), .ZN(n17839) );
  INV_X1 U11249 ( .A(n17840), .ZN(n17841) );
  INV_X1 U11250 ( .A(n17842), .ZN(n17843) );
  INV_X1 U11251 ( .A(n17844), .ZN(n17845) );
  INV_X1 U11252 ( .A(n17846), .ZN(n17847) );
  INV_X1 U11253 ( .A(n17848), .ZN(n17849) );
  INV_X1 U11254 ( .A(n17850), .ZN(n17851) );
  INV_X1 U11255 ( .A(n17852), .ZN(n17853) );
  INV_X1 U11256 ( .A(n17854), .ZN(n17855) );
  INV_X1 U11257 ( .A(n17856), .ZN(n17857) );
  INV_X1 U11258 ( .A(n17858), .ZN(n17859) );
  INV_X1 U11259 ( .A(n17860), .ZN(n17861) );
  INV_X1 U11260 ( .A(n17862), .ZN(n17863) );
  INV_X1 U11261 ( .A(n17864), .ZN(n17865) );
  INV_X1 U11262 ( .A(n17866), .ZN(n17867) );
  INV_X1 U11263 ( .A(n17868), .ZN(n17869) );
  INV_X1 U11264 ( .A(n17870), .ZN(n17871) );
  INV_X1 U11265 ( .A(n17872), .ZN(n17873) );
  INV_X1 U11266 ( .A(n17874), .ZN(n17875) );
  INV_X1 U11267 ( .A(n17876), .ZN(n17877) );
  INV_X1 U11268 ( .A(n17878), .ZN(n17879) );
  INV_X1 U11269 ( .A(n17880), .ZN(n17881) );
  INV_X1 U11270 ( .A(n17882), .ZN(n17883) );
  INV_X1 U11271 ( .A(n17884), .ZN(n17885) );
  INV_X1 U11272 ( .A(n17886), .ZN(n17887) );
  INV_X1 U11273 ( .A(n17888), .ZN(n17889) );
  INV_X1 U11274 ( .A(n17890), .ZN(n17891) );
  INV_X1 U11275 ( .A(n17892), .ZN(n17893) );
  INV_X1 U11276 ( .A(n17894), .ZN(n17895) );
  INV_X1 U11277 ( .A(n17896), .ZN(n17897) );
  INV_X1 U11278 ( .A(n17898), .ZN(n17899) );
  INV_X1 U11279 ( .A(n17900), .ZN(n17901) );
  INV_X1 U11280 ( .A(n17902), .ZN(n17903) );
  INV_X1 U11281 ( .A(n17904), .ZN(n17905) );
  INV_X1 U11282 ( .A(n17906), .ZN(n17907) );
  INV_X1 U11283 ( .A(n17908), .ZN(n17909) );
  INV_X1 U11284 ( .A(n17910), .ZN(n17911) );
  INV_X1 U11285 ( .A(n17912), .ZN(n17913) );
  INV_X1 U11286 ( .A(n17914), .ZN(n17915) );
  INV_X1 U11287 ( .A(n17916), .ZN(n17917) );
  INV_X1 U11288 ( .A(n17918), .ZN(n17919) );
  INV_X1 U11289 ( .A(n17920), .ZN(n17921) );
  INV_X1 U11290 ( .A(n17922), .ZN(n17923) );
  INV_X1 U11291 ( .A(n17924), .ZN(n17925) );
  INV_X1 U11292 ( .A(n17926), .ZN(n17927) );
  INV_X1 U11293 ( .A(n17928), .ZN(n17929) );
  INV_X1 U11294 ( .A(n17930), .ZN(n17931) );
  INV_X1 U11295 ( .A(n17932), .ZN(n17933) );
  INV_X1 U11296 ( .A(n17934), .ZN(n17935) );
  INV_X1 U11297 ( .A(n17936), .ZN(n17937) );
  INV_X1 U11298 ( .A(n17938), .ZN(n17939) );
  INV_X1 U11299 ( .A(n17940), .ZN(n17941) );
  INV_X1 U11300 ( .A(n17942), .ZN(n17943) );
  INV_X1 U11301 ( .A(n17944), .ZN(n17945) );
  INV_X1 U11302 ( .A(n17946), .ZN(n17947) );
  INV_X1 U11303 ( .A(n17948), .ZN(n17949) );
  INV_X1 U11304 ( .A(n17950), .ZN(n17951) );
  INV_X1 U11305 ( .A(n17952), .ZN(n17953) );
  INV_X1 U11306 ( .A(n17954), .ZN(n17955) );
  INV_X1 U11307 ( .A(n17956), .ZN(n17957) );
  INV_X1 U11308 ( .A(n17958), .ZN(n17959) );
  INV_X1 U11309 ( .A(n17960), .ZN(n17961) );
  INV_X1 U11310 ( .A(n17962), .ZN(n17963) );
  INV_X1 U11311 ( .A(n17964), .ZN(n17965) );
  INV_X1 U11312 ( .A(n17966), .ZN(n17967) );
  INV_X1 U11313 ( .A(n17968), .ZN(n17969) );
  INV_X1 U11314 ( .A(n17970), .ZN(n17971) );
  INV_X1 U11315 ( .A(n17972), .ZN(n17973) );
  INV_X1 U11316 ( .A(n17974), .ZN(n17975) );
  INV_X1 U11317 ( .A(n17976), .ZN(n17977) );
  INV_X1 U11318 ( .A(n17978), .ZN(n17979) );
  INV_X1 U11319 ( .A(n17980), .ZN(n17981) );
  INV_X1 U11320 ( .A(n17982), .ZN(n17983) );
  INV_X1 U11321 ( .A(n17984), .ZN(n17985) );
  INV_X1 U11322 ( .A(n17986), .ZN(n17987) );
  INV_X1 U11323 ( .A(n17988), .ZN(n17989) );
  CLKBUF_X1 U11324 ( .A(n4986), .Z(n17990) );
  NAND2_X1 U11325 ( .A1(n26499), .A2(n25326), .ZN(n17991) );
  CLKBUF_X1 U11326 ( .A(n47880), .Z(n17992) );
  NAND2_X1 U11327 ( .A1(n20895), .A2(n21023), .ZN(n17993) );
  OR2_X1 U11328 ( .A1(n25607), .A2(n3482), .ZN(n17994) );
  OR2_X1 U11329 ( .A1(n22796), .A2(n45160), .ZN(n17995) );
  CLKBUF_X1 U11330 ( .A(n4569), .Z(n17996) );
  CLKBUF_X1 U11331 ( .A(n4028), .Z(n17997) );
  CLKBUF_X1 U11332 ( .A(n26973), .Z(n17998) );
  CLKBUF_X1 U11333 ( .A(n27297), .Z(n17999) );
  CLKBUF_X1 U11334 ( .A(n23423), .Z(n18000) );
  CLKBUF_X1 U11335 ( .A(n25832), .Z(n18001) );
  CLKBUF_X1 U11336 ( .A(n25846), .Z(n18002) );
  CLKBUF_X1 U11337 ( .A(n24732), .Z(n18003) );
  CLKBUF_X1 U11338 ( .A(n24734), .Z(n18004) );
  CLKBUF_X1 U11339 ( .A(n24736), .Z(n18005) );
  CLKBUF_X1 U11340 ( .A(n18946), .Z(n18006) );
  CLKBUF_X1 U11341 ( .A(n18947), .Z(n18007) );
  CLKBUF_X1 U11342 ( .A(n18948), .Z(n18008) );
  CLKBUF_X1 U11343 ( .A(n24750), .Z(n18009) );
  CLKBUF_X1 U11344 ( .A(n24753), .Z(n18010) );
  CLKBUF_X1 U11345 ( .A(n24761), .Z(n18011) );
  CLKBUF_X1 U11346 ( .A(n24763), .Z(n18012) );
  CLKBUF_X1 U11347 ( .A(n24765), .Z(n18013) );
  CLKBUF_X1 U11348 ( .A(n24770), .Z(n18014) );
  CLKBUF_X1 U11349 ( .A(n24777), .Z(n18015) );
  CLKBUF_X1 U11350 ( .A(n24779), .Z(n18016) );
  CLKBUF_X1 U11351 ( .A(n24784), .Z(n18017) );
  CLKBUF_X1 U11352 ( .A(n24787), .Z(n18018) );
  CLKBUF_X1 U11353 ( .A(n24795), .Z(n18019) );
  CLKBUF_X1 U11354 ( .A(n24797), .Z(n18020) );
  CLKBUF_X1 U11355 ( .A(n24799), .Z(n18021) );
  CLKBUF_X1 U11356 ( .A(n18952), .Z(n18022) );
  CLKBUF_X1 U11357 ( .A(n18953), .Z(n18023) );
  CLKBUF_X1 U11358 ( .A(n24803), .Z(n18024) );
  CLKBUF_X1 U11359 ( .A(n24805), .Z(n18025) );
  CLKBUF_X1 U11360 ( .A(n24807), .Z(n18026) );
  CLKBUF_X1 U11361 ( .A(n18954), .Z(n18027) );
  CLKBUF_X1 U11362 ( .A(n24812), .Z(n18028) );
  CLKBUF_X1 U11363 ( .A(n18956), .Z(n18029) );
  CLKBUF_X1 U11364 ( .A(n24816), .Z(n18030) );
  CLKBUF_X1 U11365 ( .A(n18957), .Z(n18031) );
  CLKBUF_X1 U11366 ( .A(n18958), .Z(n18032) );
  CLKBUF_X1 U11367 ( .A(n24820), .Z(n18033) );
  CLKBUF_X1 U11368 ( .A(n18959), .Z(n18034) );
  CLKBUF_X1 U11369 ( .A(n18961), .Z(n18035) );
  CLKBUF_X1 U11370 ( .A(n18964), .Z(n18036) );
  CLKBUF_X1 U11371 ( .A(n18967), .Z(n18037) );
  CLKBUF_X1 U11372 ( .A(n18970), .Z(n18038) );
  CLKBUF_X1 U11373 ( .A(n18972), .Z(n18039) );
  CLKBUF_X1 U11374 ( .A(n18975), .Z(n18040) );
  CLKBUF_X1 U11375 ( .A(n18977), .Z(n18041) );
  CLKBUF_X1 U11376 ( .A(n18980), .Z(n18042) );
  CLKBUF_X1 U11377 ( .A(n18981), .Z(n18043) );
  CLKBUF_X1 U11378 ( .A(n18982), .Z(n18044) );
  CLKBUF_X1 U11379 ( .A(n26903), .Z(n18045) );
  CLKBUF_X1 U11380 ( .A(n18983), .Z(n18046) );
  CLKBUF_X1 U11381 ( .A(n24865), .Z(n18047) );
  CLKBUF_X1 U11382 ( .A(n24867), .Z(n18048) );
  CLKBUF_X1 U11383 ( .A(n24869), .Z(n18049) );
  CLKBUF_X1 U11384 ( .A(n24871), .Z(n18050) );
  CLKBUF_X1 U11385 ( .A(n24887), .Z(n18051) );
  CLKBUF_X1 U11386 ( .A(n24892), .Z(n18052) );
  CLKBUF_X1 U11387 ( .A(n24895), .Z(n18053) );
  CLKBUF_X1 U11388 ( .A(n24897), .Z(n18054) );
  CLKBUF_X1 U11389 ( .A(n24899), .Z(n18055) );
  CLKBUF_X1 U11390 ( .A(n24901), .Z(n18056) );
  CLKBUF_X1 U11391 ( .A(n24903), .Z(n18057) );
  CLKBUF_X1 U11392 ( .A(n24905), .Z(n18058) );
  CLKBUF_X1 U11393 ( .A(n24909), .Z(n18059) );
  CLKBUF_X1 U11394 ( .A(n24911), .Z(n18060) );
  CLKBUF_X1 U11395 ( .A(n18987), .Z(n18061) );
  CLKBUF_X1 U11396 ( .A(n24916), .Z(n18062) );
  CLKBUF_X1 U11397 ( .A(n18988), .Z(n18063) );
  CLKBUF_X1 U11398 ( .A(n24946), .Z(n18064) );
  CLKBUF_X1 U11399 ( .A(n24948), .Z(n18065) );
  CLKBUF_X1 U11400 ( .A(n24950), .Z(n18066) );
  CLKBUF_X1 U11401 ( .A(n24953), .Z(n18067) );
  CLKBUF_X1 U11402 ( .A(n24955), .Z(n18068) );
  CLKBUF_X1 U11403 ( .A(n24957), .Z(n18069) );
  CLKBUF_X1 U11404 ( .A(n24960), .Z(n18070) );
  CLKBUF_X1 U11405 ( .A(n24962), .Z(n18071) );
  CLKBUF_X1 U11406 ( .A(n24964), .Z(n18072) );
  CLKBUF_X1 U11407 ( .A(n24967), .Z(n18073) );
  CLKBUF_X1 U11408 ( .A(n24969), .Z(n18074) );
  CLKBUF_X1 U11409 ( .A(n24972), .Z(n18075) );
  CLKBUF_X1 U11410 ( .A(n24986), .Z(n18076) );
  CLKBUF_X1 U11411 ( .A(n24988), .Z(n18077) );
  CLKBUF_X1 U11412 ( .A(n24990), .Z(n18078) );
  CLKBUF_X1 U11413 ( .A(n24995), .Z(n18079) );
  CLKBUF_X1 U11414 ( .A(n19000), .Z(n18080) );
  CLKBUF_X1 U11415 ( .A(n24998), .Z(n18081) );
  CLKBUF_X1 U11416 ( .A(n25003), .Z(n18082) );
  CLKBUF_X1 U11417 ( .A(n25005), .Z(n18083) );
  CLKBUF_X1 U11418 ( .A(n25007), .Z(n18084) );
  CLKBUF_X1 U11419 ( .A(n25009), .Z(n18085) );
  CLKBUF_X1 U11420 ( .A(n25011), .Z(n18086) );
  CLKBUF_X1 U11421 ( .A(n19001), .Z(n18087) );
  CLKBUF_X1 U11422 ( .A(n25028), .Z(n18088) );
  CLKBUF_X1 U11423 ( .A(n25032), .Z(n18089) );
  CLKBUF_X1 U11424 ( .A(n25064), .Z(n18090) );
  CLKBUF_X1 U11425 ( .A(n25067), .Z(n18091) );
  CLKBUF_X1 U11426 ( .A(n25069), .Z(n18092) );
  CLKBUF_X1 U11427 ( .A(n25071), .Z(n18093) );
  CLKBUF_X1 U11428 ( .A(n25073), .Z(n18094) );
  CLKBUF_X1 U11429 ( .A(n27188), .Z(n18095) );
  CLKBUF_X1 U11430 ( .A(n25077), .Z(n18096) );
  CLKBUF_X1 U11431 ( .A(n27244), .Z(n18097) );
  CLKBUF_X1 U11432 ( .A(n19018), .Z(n18098) );
  NAND4_X1 U11433 ( .A1(N4509), .A2(n22472), .A3(n22435), .A4(n44420), .ZN(
        n18099) );
  NAND4_X1 U11434 ( .A1(N2985), .A2(n22469), .A3(n22433), .A4(n4026), .ZN(
        n18100) );
  CLKBUF_X1 U11435 ( .A(n26646), .Z(n18101) );
  CLKBUF_X1 U11436 ( .A(n25659), .Z(n18102) );
  CLKBUF_X1 U11437 ( .A(n20920), .Z(n18103) );
  CLKBUF_X1 U11438 ( .A(n27152), .Z(n18104) );
  CLKBUF_X1 U11439 ( .A(n20925), .Z(n18105) );
  CLKBUF_X1 U11440 ( .A(n26638), .Z(n18106) );
  CLKBUF_X1 U11441 ( .A(n26640), .Z(n18107) );
  CLKBUF_X1 U11442 ( .A(n27157), .Z(n18108) );
  CLKBUF_X1 U11443 ( .A(n27245), .Z(n18109) );
  CLKBUF_X1 U11444 ( .A(n27173), .Z(n18110) );
  CLKBUF_X1 U11445 ( .A(n27229), .Z(n18111) );
  CLKBUF_X1 U11446 ( .A(n27227), .Z(n18112) );
  CLKBUF_X1 U11447 ( .A(n27226), .Z(n18113) );
  CLKBUF_X1 U11448 ( .A(n27173), .Z(n18114) );
  CLKBUF_X1 U11449 ( .A(n17136), .Z(n18115) );
  CLKBUF_X1 U11450 ( .A(n24581), .Z(n18116) );
  CLKBUF_X1 U11451 ( .A(n24578), .Z(n18117) );
  CLKBUF_X1 U11452 ( .A(n24564), .Z(n18118) );
  CLKBUF_X1 U11453 ( .A(n25165), .Z(n18119) );
  CLKBUF_X1 U11454 ( .A(n25169), .Z(n18120) );
  CLKBUF_X1 U11455 ( .A(n24547), .Z(n18121) );
  CLKBUF_X1 U11456 ( .A(n27029), .Z(n18122) );
  CLKBUF_X1 U11457 ( .A(n22895), .Z(n18123) );
  CLKBUF_X1 U11458 ( .A(n27265), .Z(n18124) );
  CLKBUF_X1 U11459 ( .A(n27264), .Z(n18125) );
  CLKBUF_X1 U11460 ( .A(n27155), .Z(n18126) );
  CLKBUF_X1 U11461 ( .A(n24810), .Z(n18127) );
  CLKBUF_X1 U11462 ( .A(n26935), .Z(n18128) );
  CLKBUF_X1 U11463 ( .A(n26936), .Z(n18129) );
  CLKBUF_X1 U11464 ( .A(n26933), .Z(n18130) );
  CLKBUF_X1 U11465 ( .A(n26934), .Z(n18131) );
  CLKBUF_X1 U11466 ( .A(n26931), .Z(n18132) );
  CLKBUF_X1 U11467 ( .A(n26932), .Z(n18133) );
  CLKBUF_X1 U11468 ( .A(n26929), .Z(n18134) );
  CLKBUF_X1 U11469 ( .A(n269301), .Z(n18135) );
  CLKBUF_X1 U11470 ( .A(n20999), .Z(n18136) );
  CLKBUF_X1 U11471 ( .A(n26928), .Z(n18137) );
  CLKBUF_X1 U11472 ( .A(n21057), .Z(n18138) );
  CLKBUF_X1 U11473 ( .A(n26901), .Z(n18139) );
  CLKBUF_X1 U11474 ( .A(n26905), .Z(n18140) );
  CLKBUF_X1 U11475 ( .A(n22802), .Z(n18141) );
  CLKBUF_X1 U11476 ( .A(n18852), .Z(n18142) );
  CLKBUF_X1 U11477 ( .A(n25286), .Z(n18143) );
  CLKBUF_X1 U11478 ( .A(n24182), .Z(n18144) );
  CLKBUF_X1 U11479 ( .A(n25293), .Z(n18145) );
  CLKBUF_X1 U11480 ( .A(n24177), .Z(n18146) );
  CLKBUF_X1 U11481 ( .A(n25301), .Z(n18147) );
  CLKBUF_X1 U11482 ( .A(n22794), .Z(n18148) );
  CLKBUF_X1 U11483 ( .A(n19755), .Z(n18149) );
  CLKBUF_X1 U11484 ( .A(n22790), .Z(n18150) );
  CLKBUF_X1 U11485 ( .A(n22792), .Z(n18151) );
  CLKBUF_X1 U11486 ( .A(n27791), .Z(n18152) );
  CLKBUF_X1 U11487 ( .A(n22786), .Z(n18153) );
  CLKBUF_X1 U11488 ( .A(n26691), .Z(n18154) );
  CLKBUF_X1 U11489 ( .A(n26662), .Z(n18155) );
  CLKBUF_X1 U11490 ( .A(n26663), .Z(n18156) );
  CLKBUF_X1 U11491 ( .A(n26660), .Z(n18157) );
  CLKBUF_X1 U11492 ( .A(n26661), .Z(n18158) );
  CLKBUF_X1 U11493 ( .A(n26658), .Z(n18159) );
  CLKBUF_X1 U11494 ( .A(n26659), .Z(n18160) );
  CLKBUF_X1 U11495 ( .A(n26656), .Z(n18161) );
  CLKBUF_X1 U11496 ( .A(n26657), .Z(n18162) );
  CLKBUF_X1 U11497 ( .A(n21056), .Z(n18163) );
  CLKBUF_X1 U11498 ( .A(n26655), .Z(n18164) );
  CLKBUF_X1 U11499 ( .A(n26618), .Z(n18165) );
  CLKBUF_X1 U11500 ( .A(n21061), .Z(n18166) );
  CLKBUF_X1 U11501 ( .A(n21064), .Z(n18167) );
  CLKBUF_X1 U11502 ( .A(n26574), .Z(n18168) );
  CLKBUF_X1 U11503 ( .A(n26574), .Z(n18169) );
  CLKBUF_X1 U11504 ( .A(n265601), .Z(n18170) );
  CLKBUF_X1 U11505 ( .A(n26561), .Z(n18171) );
  CLKBUF_X1 U11506 ( .A(n22952), .Z(n18172) );
  CLKBUF_X1 U11507 ( .A(n21139), .Z(n18173) );
  CLKBUF_X1 U11508 ( .A(n21145), .Z(n18174) );
  CLKBUF_X1 U11509 ( .A(n26991), .Z(n18175) );
  CLKBUF_X1 U11510 ( .A(n21149), .Z(n18176) );
  CLKBUF_X1 U11511 ( .A(n27269), .Z(n18177) );
  CLKBUF_X1 U11512 ( .A(n21152), .Z(n18178) );
  CLKBUF_X1 U11513 ( .A(n21327), .Z(n18179) );
  CLKBUF_X1 U11514 ( .A(n21155), .Z(n18180) );
  CLKBUF_X1 U11515 ( .A(n27147), .Z(n18181) );
  CLKBUF_X1 U11516 ( .A(n21158), .Z(n18182) );
  CLKBUF_X1 U11517 ( .A(n21166), .Z(n18183) );
  CLKBUF_X1 U11518 ( .A(n27156), .Z(n18184) );
  CLKBUF_X1 U11519 ( .A(n21169), .Z(n18185) );
  CLKBUF_X1 U11520 ( .A(n17992), .Z(n18186) );
  CLKBUF_X1 U11521 ( .A(n21177), .Z(n18187) );
  CLKBUF_X1 U11522 ( .A(n21184), .Z(n18188) );
  CLKBUF_X1 U11523 ( .A(n24569), .Z(n18189) );
  CLKBUF_X1 U11524 ( .A(n21191), .Z(n18190) );
  CLKBUF_X1 U11525 ( .A(n25173), .Z(n18191) );
  CLKBUF_X1 U11526 ( .A(n21194), .Z(n18192) );
  CLKBUF_X1 U11527 ( .A(n25543), .Z(n18193) );
  CLKBUF_X1 U11528 ( .A(n21197), .Z(n18194) );
  CLKBUF_X1 U11529 ( .A(n24552), .Z(n18195) );
  CLKBUF_X1 U11530 ( .A(n21200), .Z(n18196) );
  CLKBUF_X1 U11531 ( .A(n25175), .Z(n18197) );
  CLKBUF_X1 U11532 ( .A(n21203), .Z(n18198) );
  CLKBUF_X1 U11533 ( .A(n25556), .Z(n18199) );
  CLKBUF_X1 U11534 ( .A(n21206), .Z(n18200) );
  CLKBUF_X1 U11535 ( .A(n21210), .Z(n18201) );
  CLKBUF_X1 U11536 ( .A(n21214), .Z(n18202) );
  CLKBUF_X1 U11537 ( .A(n25547), .Z(n18203) );
  CLKBUF_X1 U11538 ( .A(n21217), .Z(n18204) );
  CLKBUF_X1 U11539 ( .A(n4990), .Z(n18205) );
  CLKBUF_X1 U11540 ( .A(n21220), .Z(n18206) );
  CLKBUF_X1 U11541 ( .A(n25561), .Z(n18207) );
  CLKBUF_X1 U11542 ( .A(n21223), .Z(n18208) );
  CLKBUF_X1 U11543 ( .A(n21226), .Z(n18209) );
  CLKBUF_X1 U11544 ( .A(n20484), .Z(n18210) );
  CLKBUF_X1 U11545 ( .A(n21231), .Z(n18211) );
  CLKBUF_X1 U11546 ( .A(n21238), .Z(n18212) );
  CLKBUF_X1 U11547 ( .A(n4985), .Z(n18213) );
  CLKBUF_X1 U11548 ( .A(n21245), .Z(n18214) );
  CLKBUF_X1 U11549 ( .A(n20487), .Z(n18215) );
  CLKBUF_X1 U11550 ( .A(n27223), .Z(n18216) );
  CLKBUF_X1 U11551 ( .A(n21255), .Z(n18217) );
  CLKBUF_X1 U11552 ( .A(n21252), .Z(n18218) );
  CLKBUF_X1 U11553 ( .A(n27224), .Z(n18219) );
  CLKBUF_X1 U11554 ( .A(n4989), .Z(n18220) );
  CLKBUF_X1 U11555 ( .A(n21257), .Z(n18221) );
  CLKBUF_X1 U11556 ( .A(n20546), .Z(n18222) );
  CLKBUF_X1 U11557 ( .A(n21260), .Z(n18223) );
  CLKBUF_X1 U11558 ( .A(n21263), .Z(n18224) );
  CLKBUF_X1 U11559 ( .A(n20480), .Z(n18225) );
  CLKBUF_X1 U11560 ( .A(n27200), .Z(n18226) );
  CLKBUF_X1 U11561 ( .A(n27202), .Z(n18227) );
  CLKBUF_X1 U11562 ( .A(n21270), .Z(n18228) );
  CLKBUF_X1 U11563 ( .A(n21272), .Z(n18229) );
  CLKBUF_X1 U11564 ( .A(n20585), .Z(n18230) );
  CLKBUF_X1 U11565 ( .A(n21275), .Z(n18231) );
  CLKBUF_X1 U11566 ( .A(n24218), .Z(n18232) );
  CLKBUF_X1 U11567 ( .A(n21278), .Z(n18233) );
  CLKBUF_X1 U11568 ( .A(n21285), .Z(n18234) );
  CLKBUF_X1 U11569 ( .A(n21289), .Z(n18235) );
  CLKBUF_X1 U11570 ( .A(n24210), .Z(n18236) );
  CLKBUF_X1 U11571 ( .A(n21292), .Z(n18237) );
  CLKBUF_X1 U11572 ( .A(n25260), .Z(n18238) );
  CLKBUF_X1 U11573 ( .A(n21295), .Z(n18239) );
  CLKBUF_X1 U11574 ( .A(n26736), .Z(n18240) );
  CLKBUF_X1 U11575 ( .A(n21298), .Z(n18241) );
  CLKBUF_X1 U11576 ( .A(n26737), .Z(n18242) );
  CLKBUF_X1 U11577 ( .A(n21301), .Z(n18243) );
  CLKBUF_X1 U11578 ( .A(n24204), .Z(n18244) );
  CLKBUF_X1 U11579 ( .A(n21304), .Z(n18245) );
  CLKBUF_X1 U11580 ( .A(n25269), .Z(n18246) );
  CLKBUF_X1 U11581 ( .A(n21307), .Z(n18247) );
  CLKBUF_X1 U11582 ( .A(n24198), .Z(n18248) );
  CLKBUF_X1 U11583 ( .A(n21310), .Z(n18249) );
  CLKBUF_X1 U11584 ( .A(n25274), .Z(n18250) );
  CLKBUF_X1 U11585 ( .A(n21313), .Z(n18251) );
  CLKBUF_X1 U11586 ( .A(n24195), .Z(n18252) );
  CLKBUF_X1 U11587 ( .A(n21316), .Z(n18253) );
  CLKBUF_X1 U11588 ( .A(n25278), .Z(n18254) );
  CLKBUF_X1 U11589 ( .A(n21319), .Z(n18255) );
  CLKBUF_X1 U11590 ( .A(n22801), .Z(n18256) );
  CLKBUF_X1 U11591 ( .A(n21322), .Z(n18257) );
  NAND2_X1 U11592 ( .A1(n24705), .A2(n5297), .ZN(n18258) );
  CLKBUF_X1 U11593 ( .A(n4890), .Z(n18259) );
  CLKBUF_X1 U11594 ( .A(n21332), .Z(n18260) );
  CLKBUF_X1 U11595 ( .A(n27061), .Z(n18261) );
  CLKBUF_X1 U11596 ( .A(n21339), .Z(n18262) );
  NAND2_X1 U11597 ( .A1(n265001), .A2(n26328), .ZN(n18263) );
  CLKBUF_X1 U11598 ( .A(n27098), .Z(n18264) );
  CLKBUF_X1 U11599 ( .A(n21346), .Z(n18265) );
  CLKBUF_X1 U11600 ( .A(n4885), .Z(n18266) );
  CLKBUF_X1 U11601 ( .A(n21349), .Z(n18267) );
  NAND2_X1 U11602 ( .A1(n22422), .A2(n21510), .ZN(n18268) );
  CLKBUF_X1 U11603 ( .A(n5205), .Z(n18269) );
  CLKBUF_X1 U11604 ( .A(n21360), .Z(n18270) );
  NAND2_X1 U11605 ( .A1(n19227), .A2(n21631), .ZN(n18271) );
  NAND3_X1 U11606 ( .A1(n26376), .A2(n17102), .A3(n19227), .ZN(n18272) );
  CLKBUF_X1 U11607 ( .A(n27043), .Z(n18273) );
  CLKBUF_X1 U11608 ( .A(n21387), .Z(n18274) );
  CLKBUF_X1 U11609 ( .A(n17132), .Z(n18275) );
  CLKBUF_X1 U11610 ( .A(n21391), .Z(n18276) );
  NAND4_X1 U11611 ( .A1(N2811), .A2(n26083), .A3(n21868), .A4(n3663), .ZN(
        n18277) );
  CLKBUF_X1 U11612 ( .A(n20900), .Z(n18278) );
  CLKBUF_X1 U11613 ( .A(n20905), .Z(n18279) );
  CLKBUF_X1 U11614 ( .A(n23012), .Z(n18280) );
  CLKBUF_X1 U11615 ( .A(n21402), .Z(n18281) );
  CLKBUF_X1 U11616 ( .A(n23066), .Z(n18282) );
  CLKBUF_X1 U11617 ( .A(n25894), .Z(n18283) );
  CLKBUF_X1 U11618 ( .A(n23101), .Z(n18284) );
  CLKBUF_X1 U11619 ( .A(n23103), .Z(n18285) );
  CLKBUF_X1 U11620 ( .A(n23105), .Z(n18286) );
  CLKBUF_X1 U11621 ( .A(n23107), .Z(n18287) );
  CLKBUF_X1 U11622 ( .A(n23115), .Z(n18288) );
  CLKBUF_X1 U11623 ( .A(n23121), .Z(n18289) );
  CLKBUF_X1 U11624 ( .A(n23123), .Z(n18290) );
  CLKBUF_X1 U11625 ( .A(n23125), .Z(n18291) );
  CLKBUF_X1 U11626 ( .A(n23134), .Z(n18292) );
  CLKBUF_X1 U11627 ( .A(n23143), .Z(n18293) );
  CLKBUF_X1 U11628 ( .A(n23148), .Z(n18294) );
  CLKBUF_X1 U11629 ( .A(n23150), .Z(n18295) );
  CLKBUF_X1 U11630 ( .A(n23155), .Z(n18296) );
  CLKBUF_X1 U11631 ( .A(n23160), .Z(n18297) );
  CLKBUF_X1 U11632 ( .A(n23165), .Z(n18298) );
  CLKBUF_X1 U11633 ( .A(n23174), .Z(n18299) );
  CLKBUF_X1 U11634 ( .A(n23176), .Z(n18300) );
  CLKBUF_X1 U11635 ( .A(n23178), .Z(n18301) );
  CLKBUF_X1 U11636 ( .A(n23186), .Z(n18302) );
  CLKBUF_X1 U11637 ( .A(n23188), .Z(n18303) );
  CLKBUF_X1 U11638 ( .A(n23194), .Z(n18304) );
  CLKBUF_X1 U11639 ( .A(n26561), .Z(n18305) );
  CLKBUF_X1 U11640 ( .A(n23196), .Z(n18306) );
  CLKBUF_X1 U11641 ( .A(n23198), .Z(n18307) );
  CLKBUF_X1 U11642 ( .A(n23200), .Z(n18308) );
  CLKBUF_X1 U11643 ( .A(n23205), .Z(n18309) );
  CLKBUF_X1 U11644 ( .A(n23207), .Z(n18310) );
  CLKBUF_X1 U11645 ( .A(n23209), .Z(n18311) );
  CLKBUF_X1 U11646 ( .A(n23213), .Z(n18312) );
  CLKBUF_X1 U11647 ( .A(n23216), .Z(n18313) );
  CLKBUF_X1 U11648 ( .A(n17111), .Z(n18314) );
  CLKBUF_X1 U11649 ( .A(n23217), .Z(n18315) );
  CLKBUF_X1 U11650 ( .A(n23219), .Z(n18316) );
  CLKBUF_X1 U11651 ( .A(n23222), .Z(n18317) );
  CLKBUF_X1 U11652 ( .A(n23225), .Z(n18318) );
  CLKBUF_X1 U11653 ( .A(n23224), .Z(n18319) );
  CLKBUF_X1 U11654 ( .A(n23226), .Z(n18320) );
  CLKBUF_X1 U11655 ( .A(n23228), .Z(n18321) );
  CLKBUF_X1 U11656 ( .A(n23227), .Z(n18322) );
  CLKBUF_X1 U11657 ( .A(n23230), .Z(n18323) );
  CLKBUF_X1 U11658 ( .A(n23231), .Z(n18324) );
  CLKBUF_X1 U11659 ( .A(n23232), .Z(n18325) );
  CLKBUF_X1 U11660 ( .A(n23236), .Z(n18326) );
  CLKBUF_X1 U11661 ( .A(n23237), .Z(n18327) );
  CLKBUF_X1 U11662 ( .A(n23238), .Z(n18328) );
  CLKBUF_X1 U11663 ( .A(n23239), .Z(n18329) );
  CLKBUF_X1 U11664 ( .A(n23242), .Z(n18330) );
  CLKBUF_X1 U11665 ( .A(n23241), .Z(n18331) );
  CLKBUF_X1 U11666 ( .A(n23244), .Z(n18332) );
  CLKBUF_X1 U11667 ( .A(n23243), .Z(n18333) );
  CLKBUF_X1 U11668 ( .A(n23246), .Z(n18334) );
  CLKBUF_X1 U11669 ( .A(n23245), .Z(n18335) );
  CLKBUF_X1 U11670 ( .A(n23248), .Z(n18336) );
  CLKBUF_X1 U11671 ( .A(n23247), .Z(n18337) );
  CLKBUF_X1 U11672 ( .A(n23250), .Z(n18338) );
  CLKBUF_X1 U11673 ( .A(n23249), .Z(n18339) );
  CLKBUF_X1 U11674 ( .A(n23252), .Z(n18340) );
  CLKBUF_X1 U11675 ( .A(n23251), .Z(n18341) );
  CLKBUF_X1 U11676 ( .A(n23254), .Z(n18342) );
  CLKBUF_X1 U11677 ( .A(n23253), .Z(n18343) );
  CLKBUF_X1 U11678 ( .A(n23257), .Z(n18344) );
  CLKBUF_X1 U11679 ( .A(n23256), .Z(n18345) );
  CLKBUF_X1 U11680 ( .A(n23259), .Z(n18346) );
  CLKBUF_X1 U11681 ( .A(n23258), .Z(n18347) );
  CLKBUF_X1 U11682 ( .A(n23261), .Z(n18348) );
  CLKBUF_X1 U11683 ( .A(n23260), .Z(n18349) );
  CLKBUF_X1 U11684 ( .A(n23262), .Z(n18350) );
  CLKBUF_X1 U11685 ( .A(n23263), .Z(n18351) );
  CLKBUF_X1 U11686 ( .A(n23270), .Z(n18352) );
  CLKBUF_X1 U11687 ( .A(n23271), .Z(n18353) );
  CLKBUF_X1 U11688 ( .A(n23278), .Z(n18354) );
  CLKBUF_X1 U11689 ( .A(n23279), .Z(n18355) );
  CLKBUF_X1 U11690 ( .A(n23280), .Z(n18356) );
  CLKBUF_X1 U11691 ( .A(n23281), .Z(n18357) );
  CLKBUF_X1 U11692 ( .A(n23282), .Z(n18358) );
  CLKBUF_X1 U11693 ( .A(n23283), .Z(n18359) );
  CLKBUF_X1 U11694 ( .A(n23288), .Z(n18360) );
  CLKBUF_X1 U11695 ( .A(n23289), .Z(n18361) );
  CLKBUF_X1 U11696 ( .A(n23290), .Z(n18362) );
  CLKBUF_X1 U11697 ( .A(n23291), .Z(n18363) );
  CLKBUF_X1 U11698 ( .A(n23292), .Z(n18364) );
  CLKBUF_X1 U11699 ( .A(n23293), .Z(n18365) );
  CLKBUF_X1 U11700 ( .A(n23294), .Z(n18366) );
  CLKBUF_X1 U11701 ( .A(n23295), .Z(n18367) );
  CLKBUF_X1 U11702 ( .A(n23302), .Z(n18368) );
  CLKBUF_X1 U11703 ( .A(n23303), .Z(n18369) );
  CLKBUF_X1 U11704 ( .A(n23383), .Z(n18370) );
  CLKBUF_X1 U11705 ( .A(n23384), .Z(n18371) );
  CLKBUF_X1 U11706 ( .A(n23385), .Z(n18372) );
  CLKBUF_X1 U11707 ( .A(n23386), .Z(n18373) );
  CLKBUF_X1 U11708 ( .A(n23390), .Z(n18374) );
  CLKBUF_X1 U11709 ( .A(n23391), .Z(n18375) );
  CLKBUF_X1 U11710 ( .A(n23392), .Z(n18376) );
  CLKBUF_X1 U11711 ( .A(n23393), .Z(n18377) );
  CLKBUF_X1 U11712 ( .A(n23398), .Z(n18378) );
  CLKBUF_X1 U11713 ( .A(n23399), .Z(n18379) );
  CLKBUF_X1 U11714 ( .A(n23400), .Z(n18380) );
  CLKBUF_X1 U11715 ( .A(n23401), .Z(n18381) );
  CLKBUF_X1 U11716 ( .A(n23406), .Z(n18382) );
  CLKBUF_X1 U11717 ( .A(n23405), .Z(n18383) );
  CLKBUF_X1 U11718 ( .A(n23407), .Z(n18384) );
  CLKBUF_X1 U11719 ( .A(n23408), .Z(n18385) );
  CLKBUF_X1 U11720 ( .A(n23412), .Z(n18386) );
  CLKBUF_X1 U11721 ( .A(n23413), .Z(n18387) );
  CLKBUF_X1 U11722 ( .A(n23414), .Z(n18388) );
  CLKBUF_X1 U11723 ( .A(n23415), .Z(n18389) );
  CLKBUF_X1 U11724 ( .A(n23419), .Z(n18390) );
  CLKBUF_X1 U11725 ( .A(n23420), .Z(n18391) );
  CLKBUF_X1 U11726 ( .A(n23422), .Z(n18392) );
  CLKBUF_X1 U11727 ( .A(n23421), .Z(n18393) );
  CLKBUF_X1 U11728 ( .A(n23425), .Z(n18394) );
  CLKBUF_X1 U11729 ( .A(n23426), .Z(n18395) );
  CLKBUF_X1 U11730 ( .A(n23428), .Z(n18396) );
  CLKBUF_X1 U11731 ( .A(n23427), .Z(n18397) );
  CLKBUF_X1 U11732 ( .A(n23429), .Z(n18398) );
  CLKBUF_X1 U11733 ( .A(n23430), .Z(n18399) );
  CLKBUF_X1 U11734 ( .A(n23432), .Z(n18400) );
  CLKBUF_X1 U11735 ( .A(n23431), .Z(n18401) );
  CLKBUF_X1 U11736 ( .A(n23434), .Z(n18402) );
  CLKBUF_X1 U11737 ( .A(n23433), .Z(n18403) );
  CLKBUF_X1 U11738 ( .A(n23436), .Z(n18404) );
  CLKBUF_X1 U11739 ( .A(n23435), .Z(n18405) );
  CLKBUF_X1 U11740 ( .A(n23438), .Z(n18406) );
  CLKBUF_X1 U11741 ( .A(n23437), .Z(n18407) );
  CLKBUF_X1 U11742 ( .A(n23440), .Z(n18408) );
  CLKBUF_X1 U11743 ( .A(n23439), .Z(n18409) );
  CLKBUF_X1 U11744 ( .A(n23442), .Z(n18410) );
  CLKBUF_X1 U11745 ( .A(n23441), .Z(n18411) );
  CLKBUF_X1 U11746 ( .A(n23443), .Z(n18412) );
  CLKBUF_X1 U11747 ( .A(n23444), .Z(n18413) );
  CLKBUF_X1 U11748 ( .A(n23445), .Z(n18414) );
  CLKBUF_X1 U11749 ( .A(n26513), .Z(n18415) );
  CLKBUF_X1 U11750 ( .A(n23446), .Z(n18416) );
  CLKBUF_X1 U11751 ( .A(n23448), .Z(n18417) );
  CLKBUF_X1 U11752 ( .A(n23453), .Z(n18418) );
  CLKBUF_X1 U11753 ( .A(n23455), .Z(n18419) );
  CLKBUF_X1 U11754 ( .A(n23457), .Z(n18420) );
  CLKBUF_X1 U11755 ( .A(n23459), .Z(n18421) );
  CLKBUF_X1 U11756 ( .A(n23461), .Z(n18422) );
  CLKBUF_X1 U11757 ( .A(n23463), .Z(n18423) );
  CLKBUF_X1 U11758 ( .A(n23465), .Z(n18424) );
  CLKBUF_X1 U11759 ( .A(n23467), .Z(n18425) );
  CLKBUF_X1 U11760 ( .A(n23469), .Z(n18426) );
  CLKBUF_X1 U11761 ( .A(n23471), .Z(n18427) );
  CLKBUF_X1 U11762 ( .A(n23473), .Z(n18428) );
  CLKBUF_X1 U11763 ( .A(n23475), .Z(n18429) );
  CLKBUF_X1 U11764 ( .A(n23479), .Z(n18430) );
  CLKBUF_X1 U11765 ( .A(n26375), .Z(n18431) );
  CLKBUF_X1 U11766 ( .A(n23486), .Z(n18432) );
  CLKBUF_X1 U11767 ( .A(n27154), .Z(n18433) );
  CLKBUF_X1 U11768 ( .A(n23488), .Z(n18434) );
  CLKBUF_X1 U11769 ( .A(n23491), .Z(n18435) );
  CLKBUF_X1 U11770 ( .A(n23495), .Z(n18436) );
  CLKBUF_X1 U11771 ( .A(n23497), .Z(n18437) );
  CLKBUF_X1 U11772 ( .A(n23499), .Z(n18438) );
  CLKBUF_X1 U11773 ( .A(n23590), .Z(n18439) );
  CLKBUF_X1 U11774 ( .A(n23592), .Z(n18440) );
  CLKBUF_X1 U11775 ( .A(n23594), .Z(n18441) );
  CLKBUF_X1 U11776 ( .A(n23596), .Z(n18442) );
  CLKBUF_X1 U11777 ( .A(n23598), .Z(n18443) );
  CLKBUF_X1 U11778 ( .A(n23600), .Z(n18444) );
  CLKBUF_X1 U11779 ( .A(n23602), .Z(n18445) );
  CLKBUF_X1 U11780 ( .A(n23604), .Z(n18446) );
  CLKBUF_X1 U11781 ( .A(n23640), .Z(n18447) );
  CLKBUF_X1 U11782 ( .A(n23645), .Z(n18448) );
  CLKBUF_X1 U11783 ( .A(n23647), .Z(n18449) );
  CLKBUF_X1 U11784 ( .A(n23649), .Z(n18450) );
  CLKBUF_X1 U11785 ( .A(n23673), .Z(n18451) );
  CLKBUF_X1 U11786 ( .A(n23730), .Z(n18452) );
  CLKBUF_X1 U11787 ( .A(n24822), .Z(n18453) );
  CLKBUF_X1 U11788 ( .A(n26619), .Z(n18454) );
  CLKBUF_X1 U11789 ( .A(n21062), .Z(n18455) );
  CLKBUF_X1 U11790 ( .A(n21000), .Z(n18456) );
  CLKBUF_X1 U11791 ( .A(n26626), .Z(n18457) );
  CLKBUF_X1 U11792 ( .A(n17123), .Z(n18458) );
  CLKBUF_X1 U11793 ( .A(n21065), .Z(n18459) );
  CLKBUF_X1 U11794 ( .A(n21003), .Z(n18460) );
  CLKBUF_X1 U11795 ( .A(n21058), .Z(n18461) );
  CLKBUF_X1 U11796 ( .A(n22696), .Z(n18462) );
  CLKBUF_X1 U11797 ( .A(n22700), .Z(n18463) );
  CLKBUF_X1 U11798 ( .A(n3078), .Z(n18464) );
  CLKBUF_X1 U11799 ( .A(n22703), .Z(n18465) );
  CLKBUF_X1 U11800 ( .A(n45490), .Z(n18466) );
  CLKBUF_X1 U11801 ( .A(n22706), .Z(n18467) );
  CLKBUF_X1 U11802 ( .A(n22710), .Z(n18468) );
  CLKBUF_X1 U11803 ( .A(n25739), .Z(n18469) );
  CLKBUF_X1 U11804 ( .A(n22713), .Z(n18470) );
  CLKBUF_X1 U11805 ( .A(n20921), .Z(n18471) );
  CLKBUF_X1 U11806 ( .A(n22716), .Z(n18472) );
  CLKBUF_X1 U11807 ( .A(n21406), .Z(n18473) );
  CLKBUF_X1 U11808 ( .A(n22719), .Z(n18474) );
  CLKBUF_X1 U11809 ( .A(n20926), .Z(n18475) );
  CLKBUF_X1 U11810 ( .A(n22722), .Z(n18476) );
  CLKBUF_X1 U11811 ( .A(srstn), .Z(n18477) );
  CLKBUF_X1 U11812 ( .A(n21412), .Z(n18478) );
  CLKBUF_X1 U11813 ( .A(n22729), .Z(n18479) );
  CLKBUF_X1 U11814 ( .A(n4818), .Z(n18480) );
  CLKBUF_X1 U11815 ( .A(n22747), .Z(n18481) );
  CLKBUF_X1 U11816 ( .A(n22751), .Z(n18482) );
  CLKBUF_X1 U11817 ( .A(n51360), .Z(n18483) );
  CLKBUF_X1 U11818 ( .A(n21164), .Z(n18484) );
  CLKBUF_X1 U11819 ( .A(n21171), .Z(n18485) );
  CLKBUF_X1 U11820 ( .A(n22785), .Z(n18486) );
  CLKBUF_X1 U11821 ( .A(n24169), .Z(n18487) );
  CLKBUF_X1 U11822 ( .A(n24170), .Z(n18488) );
  CLKBUF_X1 U11823 ( .A(n24173), .Z(n18489) );
  CLKBUF_X1 U11824 ( .A(n24185), .Z(n18490) );
  CLKBUF_X1 U11825 ( .A(n20580), .Z(n18491) );
  CLKBUF_X1 U11826 ( .A(n22798), .Z(n18492) );
  CLKBUF_X1 U11827 ( .A(n24193), .Z(n18493) );
  CLKBUF_X1 U11828 ( .A(n24192), .Z(n18494) );
  CLKBUF_X1 U11829 ( .A(n24213), .Z(n18495) );
  CLKBUF_X1 U11830 ( .A(n26755), .Z(n18496) );
  CLKBUF_X1 U11831 ( .A(n20719), .Z(n18497) );
  CLKBUF_X1 U11832 ( .A(n20717), .Z(n18498) );
  CLKBUF_X1 U11833 ( .A(n20718), .Z(n18499) );
  CLKBUF_X1 U11834 ( .A(n20713), .Z(n18500) );
  CLKBUF_X1 U11835 ( .A(n20711), .Z(n18501) );
  CLKBUF_X1 U11836 ( .A(n20712), .Z(n18502) );
  CLKBUF_X1 U11837 ( .A(n20709), .Z(n18503) );
  CLKBUF_X1 U11838 ( .A(n20710), .Z(n18504) );
  CLKBUF_X1 U11839 ( .A(n20708), .Z(n18505) );
  CLKBUF_X1 U11840 ( .A(n24415), .Z(n18506) );
  CLKBUF_X1 U11841 ( .A(n20621), .Z(n18507) );
  CLKBUF_X1 U11842 ( .A(n24484), .Z(n18508) );
  CLKBUF_X1 U11843 ( .A(n20556), .Z(n18509) );
  CLKBUF_X1 U11844 ( .A(n24760), .Z(n18510) );
  CLKBUF_X1 U11845 ( .A(n24485), .Z(n18511) );
  CLKBUF_X1 U11846 ( .A(n24511), .Z(n18512) );
  CLKBUF_X1 U11847 ( .A(n24675), .Z(n18513) );
  CLKBUF_X1 U11848 ( .A(n27302), .Z(n18514) );
  CLKBUF_X1 U11849 ( .A(n456), .Z(n18515) );
  CLKBUF_X1 U11850 ( .A(n24658), .Z(n18516) );
  CLKBUF_X1 U11851 ( .A(n25524), .Z(n18517) );
  CLKBUF_X1 U11852 ( .A(n24632), .Z(n18518) );
  CLKBUF_X1 U11853 ( .A(n25955), .Z(n18519) );
  CLKBUF_X1 U11854 ( .A(n27268), .Z(n18520) );
  CLKBUF_X1 U11855 ( .A(n27267), .Z(n18521) );
  CLKBUF_X1 U11856 ( .A(n25945), .Z(n18522) );
  CLKBUF_X1 U11857 ( .A(n27266), .Z(n18523) );
  CLKBUF_X1 U11858 ( .A(n25947), .Z(n18524) );
  CLKBUF_X1 U11859 ( .A(n47880), .Z(n18525) );
  CLKBUF_X1 U11860 ( .A(n25112), .Z(n18526) );
  CLKBUF_X1 U11861 ( .A(n47890), .Z(n18527) );
  CLKBUF_X1 U11862 ( .A(n25549), .Z(n18528) );
  CLKBUF_X1 U11863 ( .A(n24531), .Z(n18529) );
  CLKBUF_X1 U11864 ( .A(n22927), .Z(n18530) );
  CLKBUF_X1 U11865 ( .A(n22924), .Z(n18531) );
  CLKBUF_X1 U11866 ( .A(n22921), .Z(n18532) );
  CLKBUF_X1 U11867 ( .A(n22918), .Z(n18533) );
  CLKBUF_X1 U11868 ( .A(n25551), .Z(n18534) );
  CLKBUF_X1 U11869 ( .A(n24526), .Z(n18535) );
  CLKBUF_X1 U11870 ( .A(n22915), .Z(n18536) );
  CLKBUF_X1 U11871 ( .A(n22912), .Z(n18537) );
  CLKBUF_X1 U11872 ( .A(n22909), .Z(n18538) );
  CLKBUF_X1 U11873 ( .A(n22906), .Z(n18539) );
  CLKBUF_X1 U11874 ( .A(n21416), .Z(n18540) );
  CLKBUF_X1 U11875 ( .A(n27232), .Z(n18541) );
  CLKBUF_X1 U11876 ( .A(n21419), .Z(n18542) );
  CLKBUF_X1 U11877 ( .A(n27177), .Z(n18543) );
  CLKBUF_X1 U11878 ( .A(n20548), .Z(n18544) );
  CLKBUF_X1 U11879 ( .A(n22890), .Z(n18545) );
  CLKBUF_X1 U11880 ( .A(n24755), .Z(n18546) );
  CLKBUF_X1 U11881 ( .A(n25870), .Z(n18547) );
  CLKBUF_X1 U11882 ( .A(n24782), .Z(n18548) );
  CLKBUF_X1 U11883 ( .A(n20587), .Z(n18549) );
  CLKBUF_X1 U11884 ( .A(n22881), .Z(n18550) );
  CLKBUF_X1 U11885 ( .A(n25892), .Z(n18551) );
  CLKBUF_X1 U11886 ( .A(n24791), .Z(n18552) );
  CLKBUF_X1 U11887 ( .A(n25596), .Z(n18553) );
  CLKBUF_X1 U11888 ( .A(n25601), .Z(n18554) );
  CLKBUF_X1 U11889 ( .A(n24228), .Z(n18555) );
  CLKBUF_X1 U11890 ( .A(n24216), .Z(n18556) );
  CLKBUF_X1 U11891 ( .A(n24224), .Z(n18557) );
  CLKBUF_X1 U11892 ( .A(n25942), .Z(n18558) );
  CLKBUF_X1 U11893 ( .A(n27794), .Z(n18559) );
  CLKBUF_X1 U11894 ( .A(n20534), .Z(n18560) );
  CLKBUF_X1 U11895 ( .A(n20537), .Z(n18561) );
  CLKBUF_X1 U11896 ( .A(n25674), .Z(n18562) );
  CLKBUF_X1 U11897 ( .A(n25676), .Z(n18563) );
  CLKBUF_X1 U11898 ( .A(n25099), .Z(n18564) );
  CLKBUF_X1 U11899 ( .A(n19025), .Z(n18565) );
  CLKBUF_X1 U11900 ( .A(n20882), .Z(n18566) );
  CLKBUF_X1 U11901 ( .A(n25105), .Z(n18567) );
  CLKBUF_X1 U11902 ( .A(n19029), .Z(n18568) );
  CLKBUF_X1 U11903 ( .A(n25978), .Z(n18569) );
  CLKBUF_X1 U11904 ( .A(n24513), .Z(n18570) );
  CLKBUF_X1 U11905 ( .A(n23132), .Z(n18571) );
  CLKBUF_X1 U11906 ( .A(n25191), .Z(n18572) );
  CLKBUF_X1 U11907 ( .A(n19054), .Z(n18573) );
  CLKBUF_X1 U11908 ( .A(n23141), .Z(n18574) );
  CLKBUF_X1 U11909 ( .A(n25189), .Z(n18575) );
  CLKBUF_X1 U11910 ( .A(n19053), .Z(n18576) );
  CLKBUF_X1 U11911 ( .A(n23146), .Z(n18577) );
  CLKBUF_X1 U11912 ( .A(n24258), .Z(n18578) );
  CLKBUF_X1 U11913 ( .A(n23153), .Z(n18579) );
  CLKBUF_X1 U11914 ( .A(n24252), .Z(n18580) );
  CLKBUF_X1 U11915 ( .A(n24249), .Z(n18581) );
  CLKBUF_X1 U11916 ( .A(n23168), .Z(n18582) );
  CLKBUF_X1 U11917 ( .A(n23171), .Z(n18583) );
  CLKBUF_X1 U11918 ( .A(n23181), .Z(n18584) );
  CLKBUF_X1 U11919 ( .A(n23184), .Z(n18585) );
  CLKBUF_X1 U11920 ( .A(n24237), .Z(n18586) );
  CLKBUF_X1 U11921 ( .A(n26531), .Z(n18587) );
  CLKBUF_X1 U11922 ( .A(n22838), .Z(n18588) );
  CLKBUF_X1 U11923 ( .A(n24231), .Z(n18589) );
  CLKBUF_X1 U11924 ( .A(n21436), .Z(n18590) );
  CLKBUF_X1 U11925 ( .A(n23203), .Z(n18591) );
  CLKBUF_X1 U11926 ( .A(n22826), .Z(n18592) );
  CLKBUF_X1 U11927 ( .A(n22828), .Z(n18593) );
  CLKBUF_X1 U11928 ( .A(n30950), .Z(n18594) );
  CLKBUF_X1 U11929 ( .A(n27273), .Z(n18595) );
  CLKBUF_X1 U11930 ( .A(n27125), .Z(n18596) );
  CLKBUF_X1 U11931 ( .A(n4983), .Z(n18597) );
  CLKBUF_X1 U11932 ( .A(n4987), .Z(n18598) );
  CLKBUF_X1 U11933 ( .A(n4982), .Z(n18599) );
  CLKBUF_X1 U11934 ( .A(n27214), .Z(n18600) );
  CLKBUF_X1 U11935 ( .A(n27215), .Z(n18601) );
  CLKBUF_X1 U11936 ( .A(n19315), .Z(n18602) );
  CLKBUF_X1 U11937 ( .A(n27193), .Z(n18603) );
  CLKBUF_X1 U11938 ( .A(n27216), .Z(n18604) );
  CLKBUF_X1 U11939 ( .A(n19314), .Z(n18605) );
  CLKBUF_X1 U11940 ( .A(n27195), .Z(n18606) );
  CLKBUF_X1 U11941 ( .A(n27194), .Z(n18607) );
  CLKBUF_X1 U11942 ( .A(n20558), .Z(n18608) );
  CLKBUF_X1 U11943 ( .A(n20563), .Z(n18609) );
  CLKBUF_X1 U11944 ( .A(n20565), .Z(n18610) );
  CLKBUF_X1 U11945 ( .A(n20560), .Z(n18611) );
  CLKBUF_X1 U11946 ( .A(n20591), .Z(n18612) );
  CLKBUF_X1 U11947 ( .A(n27766), .Z(n18613) );
  CLKBUF_X1 U11948 ( .A(n25196), .Z(n18614) );
  CLKBUF_X1 U11949 ( .A(n20593), .Z(n18615) );
  CLKBUF_X1 U11950 ( .A(n20879), .Z(n18616) );
  CLKBUF_X1 U11951 ( .A(n20603), .Z(n18617) );
  CLKBUF_X1 U11952 ( .A(n20874), .Z(n18618) );
  CLKBUF_X1 U11953 ( .A(n25193), .Z(n18619) );
  CLKBUF_X1 U11954 ( .A(n20601), .Z(n18620) );
  CLKBUF_X1 U11955 ( .A(n24306), .Z(n18621) );
  CLKBUF_X1 U11956 ( .A(n24300), .Z(n18622) );
  CLKBUF_X1 U11957 ( .A(n23388), .Z(n18623) );
  CLKBUF_X1 U11958 ( .A(n24294), .Z(n18624) );
  CLKBUF_X1 U11959 ( .A(n24288), .Z(n18625) );
  CLKBUF_X1 U11960 ( .A(n23403), .Z(n18626) );
  CLKBUF_X1 U11961 ( .A(n24282), .Z(n18627) );
  CLKBUF_X1 U11962 ( .A(n23410), .Z(n18628) );
  CLKBUF_X1 U11963 ( .A(n23417), .Z(n18629) );
  CLKBUF_X1 U11964 ( .A(n24276), .Z(n18630) );
  CLKBUF_X1 U11965 ( .A(n23424), .Z(n18631) );
  CLKBUF_X1 U11966 ( .A(n24270), .Z(n18632) );
  CLKBUF_X1 U11967 ( .A(n24261), .Z(n18633) );
  CLKBUF_X1 U11968 ( .A(n24264), .Z(n18634) );
  CLKBUF_X1 U11969 ( .A(n23158), .Z(n18635) );
  CLKBUF_X1 U11970 ( .A(n24255), .Z(n18636) );
  CLKBUF_X1 U11971 ( .A(n24246), .Z(n18637) );
  CLKBUF_X1 U11972 ( .A(n23163), .Z(n18638) );
  CLKBUF_X1 U11973 ( .A(n24240), .Z(n18639) );
  CLKBUF_X1 U11974 ( .A(n27210), .Z(n18640) );
  CLKBUF_X1 U11975 ( .A(n19315), .Z(n18641) );
  CLKBUF_X1 U11976 ( .A(n27211), .Z(n18642) );
  CLKBUF_X1 U11977 ( .A(n27213), .Z(n18643) );
  CLKBUF_X1 U11978 ( .A(n27212), .Z(n18644) );
  CLKBUF_X1 U11979 ( .A(n27190), .Z(n18645) );
  CLKBUF_X1 U11980 ( .A(n27189), .Z(n18646) );
  CLKBUF_X1 U11981 ( .A(n27191), .Z(n18647) );
  CLKBUF_X1 U11982 ( .A(n19314), .Z(n18648) );
  CLKBUF_X1 U11983 ( .A(n27192), .Z(n18649) );
  CLKBUF_X1 U11984 ( .A(n26666), .Z(n18650) );
  CLKBUF_X1 U11985 ( .A(n25198), .Z(n18651) );
  CLKBUF_X1 U11986 ( .A(n25248), .Z(n18652) );
  CLKBUF_X1 U11987 ( .A(n25204), .Z(n18653) );
  CLKBUF_X1 U11988 ( .A(n24399), .Z(n18654) );
  CLKBUF_X1 U11989 ( .A(n24395), .Z(n18655) );
  CLKBUF_X1 U11990 ( .A(n26893), .Z(n18656) );
  CLKBUF_X1 U11991 ( .A(n26894), .Z(n18657) );
  CLKBUF_X1 U11992 ( .A(n268901), .Z(n18658) );
  CLKBUF_X1 U11993 ( .A(n26891), .Z(n18659) );
  CLKBUF_X1 U11994 ( .A(n26887), .Z(n18660) );
  CLKBUF_X1 U11995 ( .A(n26889), .Z(n18661) );
  CLKBUF_X1 U11996 ( .A(n26885), .Z(n18662) );
  CLKBUF_X1 U11997 ( .A(n26886), .Z(n18663) );
  CLKBUF_X1 U11998 ( .A(n26839), .Z(n18664) );
  CLKBUF_X1 U11999 ( .A(n26828), .Z(n18665) );
  CLKBUF_X1 U12000 ( .A(n26831), .Z(n18666) );
  CLKBUF_X1 U12001 ( .A(n26832), .Z(n18667) );
  CLKBUF_X1 U12002 ( .A(n26864), .Z(n18668) );
  CLKBUF_X1 U12003 ( .A(n26863), .Z(n18669) );
  CLKBUF_X1 U12004 ( .A(n26862), .Z(n18670) );
  CLKBUF_X1 U12005 ( .A(n26861), .Z(n18671) );
  CLKBUF_X1 U12006 ( .A(n268601), .Z(n18672) );
  CLKBUF_X1 U12007 ( .A(n26859), .Z(n18673) );
  CLKBUF_X1 U12008 ( .A(n26858), .Z(n18674) );
  CLKBUF_X1 U12009 ( .A(n26857), .Z(n18675) );
  CLKBUF_X1 U12010 ( .A(n26856), .Z(n18676) );
  CLKBUF_X1 U12011 ( .A(n24861), .Z(n18677) );
  CLKBUF_X1 U12012 ( .A(n23585), .Z(n18678) );
  CLKBUF_X1 U12013 ( .A(n24360), .Z(n18679) );
  CLKBUF_X1 U12014 ( .A(n23333), .Z(n18680) );
  CLKBUF_X1 U12015 ( .A(n23336), .Z(n18681) );
  CLKBUF_X1 U12016 ( .A(n24351), .Z(n18682) );
  CLKBUF_X1 U12017 ( .A(n23339), .Z(n18683) );
  CLKBUF_X1 U12018 ( .A(n24345), .Z(n18684) );
  CLKBUF_X1 U12019 ( .A(n23342), .Z(n18685) );
  CLKBUF_X1 U12020 ( .A(n24339), .Z(n18686) );
  CLKBUF_X1 U12021 ( .A(n26838), .Z(n18687) );
  CLKBUF_X1 U12022 ( .A(n26837), .Z(n18688) );
  CLKBUF_X1 U12023 ( .A(n26834), .Z(n18689) );
  CLKBUF_X1 U12024 ( .A(n26833), .Z(n18690) );
  CLKBUF_X1 U12025 ( .A(n268301), .Z(n18691) );
  CLKBUF_X1 U12026 ( .A(n26829), .Z(n18692) );
  CLKBUF_X1 U12027 ( .A(n26826), .Z(n18693) );
  CLKBUF_X1 U12028 ( .A(n26825), .Z(n18694) );
  CLKBUF_X1 U12029 ( .A(n26822), .Z(n18695) );
  CLKBUF_X1 U12030 ( .A(n26821), .Z(n18696) );
  CLKBUF_X1 U12031 ( .A(n26818), .Z(n18697) );
  CLKBUF_X1 U12032 ( .A(n26817), .Z(n18698) );
  CLKBUF_X1 U12033 ( .A(n26814), .Z(n18699) );
  CLKBUF_X1 U12034 ( .A(n26813), .Z(n18700) );
  CLKBUF_X1 U12035 ( .A(n268101), .Z(n18701) );
  CLKBUF_X1 U12036 ( .A(n26809), .Z(n18702) );
  CLKBUF_X1 U12037 ( .A(n24309), .Z(n18703) );
  CLKBUF_X1 U12038 ( .A(n24664), .Z(n18704) );
  CLKBUF_X1 U12039 ( .A(n27795), .Z(n18705) );
  CLKBUF_X1 U12040 ( .A(n27805), .Z(n18706) );
  CLKBUF_X1 U12041 ( .A(n25249), .Z(n18707) );
  CLKBUF_X1 U12042 ( .A(n19068), .Z(n18708) );
  CLKBUF_X1 U12043 ( .A(n20689), .Z(n18709) );
  CLKBUF_X1 U12044 ( .A(n25140), .Z(n18710) );
  CLKBUF_X1 U12045 ( .A(n25134), .Z(n18711) );
  CLKBUF_X1 U12046 ( .A(n25137), .Z(n18712) );
  CLKBUF_X1 U12047 ( .A(n25158), .Z(n18713) );
  CLKBUF_X1 U12048 ( .A(n25152), .Z(n18714) );
  CLKBUF_X1 U12049 ( .A(n25155), .Z(n18715) );
  CLKBUF_X1 U12050 ( .A(n20607), .Z(n18716) );
  CLKBUF_X1 U12051 ( .A(n20861), .Z(n18717) );
  CLKBUF_X1 U12052 ( .A(n20691), .Z(n18718) );
  CLKBUF_X1 U12053 ( .A(n23730), .Z(n18719) );
  CLKBUF_X1 U12054 ( .A(n27296), .Z(n18720) );
  CLKBUF_X1 U12055 ( .A(r899_B_2_), .Z(n18721) );
  CLKBUF_X1 U12056 ( .A(n26921), .Z(n18722) );
  CLKBUF_X1 U12057 ( .A(n23744), .Z(n18723) );
  CLKBUF_X1 U12058 ( .A(n23743), .Z(n18724) );
  CLKBUF_X1 U12059 ( .A(n269201), .Z(n18725) );
  CLKBUF_X1 U12060 ( .A(n23749), .Z(n18726) );
  CLKBUF_X1 U12061 ( .A(n23750), .Z(n18727) );
  CLKBUF_X1 U12062 ( .A(n26919), .Z(n18728) );
  CLKBUF_X1 U12063 ( .A(n23756), .Z(n18729) );
  CLKBUF_X1 U12064 ( .A(n23755), .Z(n18730) );
  CLKBUF_X1 U12065 ( .A(n26918), .Z(n18731) );
  CLKBUF_X1 U12066 ( .A(n23761), .Z(n18732) );
  CLKBUF_X1 U12067 ( .A(n23762), .Z(n18733) );
  CLKBUF_X1 U12068 ( .A(n26917), .Z(n18734) );
  CLKBUF_X1 U12069 ( .A(n23768), .Z(n18735) );
  CLKBUF_X1 U12070 ( .A(n23767), .Z(n18736) );
  CLKBUF_X1 U12071 ( .A(n26916), .Z(n18737) );
  CLKBUF_X1 U12072 ( .A(n23774), .Z(n18738) );
  CLKBUF_X1 U12073 ( .A(n23773), .Z(n18739) );
  CLKBUF_X1 U12074 ( .A(n26915), .Z(n18740) );
  CLKBUF_X1 U12075 ( .A(n23780), .Z(n18741) );
  CLKBUF_X1 U12076 ( .A(n23779), .Z(n18742) );
  CLKBUF_X1 U12077 ( .A(n26914), .Z(n18743) );
  CLKBUF_X1 U12078 ( .A(n23786), .Z(n18744) );
  CLKBUF_X1 U12079 ( .A(n23785), .Z(n18745) );
  CLKBUF_X1 U12080 ( .A(n26913), .Z(n18746) );
  CLKBUF_X1 U12081 ( .A(n23792), .Z(n18747) );
  CLKBUF_X1 U12082 ( .A(n23791), .Z(n18748) );
  CLKBUF_X1 U12083 ( .A(n26912), .Z(n18749) );
  CLKBUF_X1 U12084 ( .A(n23798), .Z(n18750) );
  CLKBUF_X1 U12085 ( .A(n23797), .Z(n18751) );
  CLKBUF_X1 U12086 ( .A(n26911), .Z(n18752) );
  CLKBUF_X1 U12087 ( .A(n23804), .Z(n18753) );
  CLKBUF_X1 U12088 ( .A(n23803), .Z(n18754) );
  CLKBUF_X1 U12089 ( .A(n269101), .Z(n18755) );
  CLKBUF_X1 U12090 ( .A(n23810), .Z(n18756) );
  CLKBUF_X1 U12091 ( .A(n23809), .Z(n18757) );
  CLKBUF_X1 U12092 ( .A(n26909), .Z(n18758) );
  CLKBUF_X1 U12093 ( .A(n23816), .Z(n18759) );
  CLKBUF_X1 U12094 ( .A(n23815), .Z(n18760) );
  CLKBUF_X1 U12095 ( .A(n26908), .Z(n18761) );
  CLKBUF_X1 U12096 ( .A(n23822), .Z(n18762) );
  CLKBUF_X1 U12097 ( .A(n23821), .Z(n18763) );
  CLKBUF_X1 U12098 ( .A(n26907), .Z(n18764) );
  CLKBUF_X1 U12099 ( .A(n23827), .Z(n18765) );
  CLKBUF_X1 U12100 ( .A(n23828), .Z(n18766) );
  CLKBUF_X1 U12101 ( .A(n26906), .Z(n18767) );
  CLKBUF_X1 U12102 ( .A(n23834), .Z(n18768) );
  CLKBUF_X1 U12103 ( .A(n23833), .Z(n18769) );
  CLKBUF_X1 U12104 ( .A(n20859), .Z(n18770) );
  CLKBUF_X1 U12105 ( .A(n23840), .Z(n18771) );
  CLKBUF_X1 U12106 ( .A(n23839), .Z(n18772) );
  CLKBUF_X1 U12107 ( .A(n20622), .Z(n18773) );
  CLKBUF_X1 U12108 ( .A(n23846), .Z(n18774) );
  CLKBUF_X1 U12109 ( .A(n23845), .Z(n18775) );
  CLKBUF_X1 U12110 ( .A(n20848), .Z(n18776) );
  CLKBUF_X1 U12111 ( .A(n23852), .Z(n18777) );
  CLKBUF_X1 U12112 ( .A(n23851), .Z(n18778) );
  CLKBUF_X1 U12113 ( .A(n20630), .Z(n18779) );
  CLKBUF_X1 U12114 ( .A(n23858), .Z(n18780) );
  CLKBUF_X1 U12115 ( .A(n23857), .Z(n18781) );
  CLKBUF_X1 U12116 ( .A(n20846), .Z(n18782) );
  CLKBUF_X1 U12117 ( .A(n23864), .Z(n18783) );
  CLKBUF_X1 U12118 ( .A(n23863), .Z(n18784) );
  CLKBUF_X1 U12119 ( .A(n20638), .Z(n18785) );
  CLKBUF_X1 U12120 ( .A(n23870), .Z(n18786) );
  CLKBUF_X1 U12121 ( .A(n23869), .Z(n18787) );
  CLKBUF_X1 U12122 ( .A(n20836), .Z(n18788) );
  CLKBUF_X1 U12123 ( .A(n23876), .Z(n18789) );
  CLKBUF_X1 U12124 ( .A(n23875), .Z(n18790) );
  CLKBUF_X1 U12125 ( .A(n20647), .Z(n18791) );
  CLKBUF_X1 U12126 ( .A(n23882), .Z(n18792) );
  CLKBUF_X1 U12127 ( .A(n23881), .Z(n18793) );
  CLKBUF_X1 U12128 ( .A(n20834), .Z(n18794) );
  CLKBUF_X1 U12129 ( .A(n23888), .Z(n18795) );
  CLKBUF_X1 U12130 ( .A(n23887), .Z(n18796) );
  CLKBUF_X1 U12131 ( .A(n20655), .Z(n18797) );
  CLKBUF_X1 U12132 ( .A(n23894), .Z(n18798) );
  CLKBUF_X1 U12133 ( .A(n23893), .Z(n18799) );
  CLKBUF_X1 U12134 ( .A(n20824), .Z(n18800) );
  CLKBUF_X1 U12135 ( .A(n23900), .Z(n18801) );
  CLKBUF_X1 U12136 ( .A(n23899), .Z(n18802) );
  CLKBUF_X1 U12137 ( .A(n20663), .Z(n18803) );
  CLKBUF_X1 U12138 ( .A(n23906), .Z(n18804) );
  CLKBUF_X1 U12139 ( .A(n23905), .Z(n18805) );
  CLKBUF_X1 U12140 ( .A(n20822), .Z(n18806) );
  CLKBUF_X1 U12141 ( .A(n23912), .Z(n18807) );
  CLKBUF_X1 U12142 ( .A(n23911), .Z(n18808) );
  CLKBUF_X1 U12143 ( .A(n20671), .Z(n18809) );
  CLKBUF_X1 U12144 ( .A(n23918), .Z(n18810) );
  CLKBUF_X1 U12145 ( .A(n23917), .Z(n18811) );
  CLKBUF_X1 U12146 ( .A(n20812), .Z(n18812) );
  CLKBUF_X1 U12147 ( .A(n23924), .Z(n18813) );
  CLKBUF_X1 U12148 ( .A(n23923), .Z(n18814) );
  CLKBUF_X1 U12149 ( .A(n20679), .Z(n18815) );
  CLKBUF_X1 U12150 ( .A(n23930), .Z(n18816) );
  CLKBUF_X1 U12151 ( .A(n23929), .Z(n18817) );
  CLKBUF_X1 U12152 ( .A(n23949), .Z(n18818) );
  CLKBUF_X1 U12153 ( .A(n26610), .Z(n18819) );
  OAI21_X1 U12154 ( .B1(n27295), .B2(n27300), .A(n17998), .ZN(r899_B_4_) );
  CLKBUF_X1 U12155 ( .A(n26614), .Z(n18820) );
  CLKBUF_X1 U12156 ( .A(n26614), .Z(n18821) );
  CLKBUF_X1 U12157 ( .A(n23960), .Z(n18822) );
  CLKBUF_X1 U12158 ( .A(n22694), .Z(n18823) );
  CLKBUF_X1 U12159 ( .A(n26942), .Z(n18824) );
  CLKBUF_X1 U12160 ( .A(n24081), .Z(n18825) );
  CLKBUF_X1 U12161 ( .A(n24081), .Z(n18826) );
  CLKBUF_X1 U12162 ( .A(n24080), .Z(n18827) );
  CLKBUF_X1 U12163 ( .A(n24105), .Z(n18828) );
  CLKBUF_X1 U12164 ( .A(n24106), .Z(n18829) );
  CLKBUF_X1 U12165 ( .A(n25223), .Z(n18830) );
  CLKBUF_X1 U12166 ( .A(n24112), .Z(n18831) );
  CLKBUF_X1 U12167 ( .A(n24111), .Z(n18832) );
  CLKBUF_X1 U12168 ( .A(n25352), .Z(n18833) );
  CLKBUF_X1 U12169 ( .A(n24117), .Z(n18834) );
  CLKBUF_X1 U12170 ( .A(n24118), .Z(n18835) );
  CLKBUF_X1 U12171 ( .A(n25233), .Z(n18836) );
  CLKBUF_X1 U12172 ( .A(n24124), .Z(n18837) );
  CLKBUF_X1 U12173 ( .A(n24123), .Z(n18838) );
  CLKBUF_X1 U12174 ( .A(n25350), .Z(n18839) );
  CLKBUF_X1 U12175 ( .A(n24129), .Z(n18840) );
  CLKBUF_X1 U12176 ( .A(n24130), .Z(n18841) );
  CLKBUF_X1 U12177 ( .A(n25235), .Z(n18842) );
  CLKBUF_X1 U12178 ( .A(n24136), .Z(n18843) );
  CLKBUF_X1 U12179 ( .A(n24135), .Z(n18844) );
  CLKBUF_X1 U12180 ( .A(n21147), .Z(n18845) );
  CLKBUF_X1 U12181 ( .A(n21140), .Z(n18846) );
  CLKBUF_X1 U12182 ( .A(n21173), .Z(n18847) );
  CLKBUF_X1 U12183 ( .A(n21180), .Z(n18848) );
  CLKBUF_X1 U12184 ( .A(n20605), .Z(n18849) );
  CLKBUF_X1 U12185 ( .A(n27803), .Z(n18850) );
  CLKBUF_X1 U12186 ( .A(n20868), .Z(n18851) );
  CLKBUF_X1 U12187 ( .A(n26724), .Z(n18852) );
  CLKBUF_X1 U12188 ( .A(n24825), .Z(n18853) );
  CLKBUF_X1 U12189 ( .A(n26943), .Z(n18854) );
  CLKBUF_X1 U12190 ( .A(n21423), .Z(n18855) );
  CLKBUF_X1 U12191 ( .A(n26944), .Z(n18856) );
  CLKBUF_X1 U12192 ( .A(n24215), .Z(n18857) );
  CLKBUF_X1 U12193 ( .A(n24214), .Z(n18858) );
  CLKBUF_X1 U12194 ( .A(n24215), .Z(n18859) );
  CLKBUF_X1 U12195 ( .A(n24861), .Z(n18860) );
  CLKBUF_X1 U12196 ( .A(n24860), .Z(n18861) );
  CLKBUF_X1 U12197 ( .A(n27113), .Z(n18862) );
  CLKBUF_X1 U12198 ( .A(n24647), .Z(n18863) );
  CLKBUF_X1 U12199 ( .A(n27124), .Z(n18864) );
  CLKBUF_X1 U12200 ( .A(n27123), .Z(n18865) );
  CLKBUF_X1 U12201 ( .A(n27122), .Z(n18866) );
  CLKBUF_X1 U12202 ( .A(n27121), .Z(n18867) );
  CLKBUF_X1 U12203 ( .A(n25248), .Z(n18868) );
  CLKBUF_X1 U12204 ( .A(n25247), .Z(n18869) );
  CLKBUF_X1 U12205 ( .A(n25247), .Z(n18870) );
  CLKBUF_X1 U12206 ( .A(n19068), .Z(n18871) );
  CLKBUF_X1 U12207 ( .A(n25250), .Z(n18872) );
  CLKBUF_X1 U12208 ( .A(n26952), .Z(n18873) );
  CLKBUF_X1 U12209 ( .A(n26951), .Z(n18874) );
  CLKBUF_X1 U12210 ( .A(n26950), .Z(n18875) );
  CLKBUF_X1 U12211 ( .A(n26949), .Z(n18876) );
  CLKBUF_X1 U12212 ( .A(n22691), .Z(n18877) );
  CLKBUF_X1 U12213 ( .A(n22685), .Z(n18878) );
  CLKBUF_X1 U12214 ( .A(n25023), .Z(n18879) );
  INV_X1 U12215 ( .A(n24428), .ZN(n26944) );
  CLKBUF_X1 U12216 ( .A(n27767), .Z(n18880) );
  INV_X1 U12217 ( .A(n26987), .ZN(n27767) );
  INV_X1 U12218 ( .A(n24433), .ZN(n26951) );
  INV_X1 U12219 ( .A(n24433), .ZN(n26949) );
  INV_X1 U12220 ( .A(n24434), .ZN(n26952) );
  CLKBUF_X1 U12221 ( .A(n24603), .Z(n18881) );
  CLKBUF_X1 U12222 ( .A(n24602), .Z(n18882) );
  CLKBUF_X1 U12223 ( .A(n24729), .Z(n18883) );
  CLKBUF_X1 U12224 ( .A(n25192), .Z(n18884) );
  CLKBUF_X1 U12225 ( .A(n25195), .Z(n18885) );
  CLKBUF_X1 U12226 ( .A(n25188), .Z(n18886) );
  CLKBUF_X1 U12227 ( .A(n25189), .Z(n18887) );
  CLKBUF_X1 U12228 ( .A(n19053), .Z(n18888) );
  CLKBUF_X1 U12229 ( .A(n25190), .Z(n18889) );
  CLKBUF_X1 U12230 ( .A(n25191), .Z(n18890) );
  CLKBUF_X1 U12231 ( .A(n19054), .Z(n18891) );
  CLKBUF_X1 U12232 ( .A(n20554), .Z(n18892) );
  CLKBUF_X1 U12233 ( .A(n20553), .Z(n18893) );
  CLKBUF_X1 U12234 ( .A(n24707), .Z(n18894) );
  CLKBUF_X1 U12235 ( .A(n20540), .Z(n18895) );
  CLKBUF_X1 U12236 ( .A(n24744), .Z(n18896) );
  CLKBUF_X1 U12237 ( .A(n20539), .Z(n18897) );
  CLKBUF_X1 U12238 ( .A(n17097), .Z(n18898) );
  CLKBUF_X1 U12239 ( .A(n20542), .Z(n18899) );
  CLKBUF_X1 U12240 ( .A(n27095), .Z(n18900) );
  CLKBUF_X1 U12241 ( .A(n27011), .Z(n18901) );
  CLKBUF_X1 U12242 ( .A(n27026), .Z(n18902) );
  CLKBUF_X1 U12243 ( .A(n24699), .Z(n18903) );
  CLKBUF_X1 U12244 ( .A(n25106), .Z(n18904) );
  CLKBUF_X1 U12245 ( .A(n19029), .Z(n18905) );
  CLKBUF_X1 U12246 ( .A(n25100), .Z(n18906) );
  CLKBUF_X1 U12247 ( .A(n19025), .Z(n18907) );
  CLKBUF_X1 U12248 ( .A(n24617), .Z(n18908) );
  CLKBUF_X1 U12249 ( .A(n24617), .Z(n18909) );
  CLKBUF_X1 U12250 ( .A(n24615), .Z(n18910) );
  CLKBUF_X1 U12251 ( .A(n24630), .Z(n18911) );
  CLKBUF_X1 U12252 ( .A(n24612), .Z(n18912) );
  CLKBUF_X1 U12253 ( .A(n24627), .Z(n18913) );
  CLKBUF_X1 U12254 ( .A(n27058), .Z(n18914) );
  CLKBUF_X1 U12255 ( .A(n27040), .Z(n18915) );
  BUF_X1 U12256 ( .A(n24602), .Z(n26965) );
  CLKBUF_X1 U12257 ( .A(n20903), .Z(n18916) );
  CLKBUF_X1 U12258 ( .A(n20908), .Z(n18917) );
  BUF_X1 U12259 ( .A(n24641), .Z(n27117) );
  BUF_X1 U12260 ( .A(n24641), .Z(n27118) );
  BUF_X1 U12261 ( .A(n24642), .Z(n27120) );
  BUF_X1 U12262 ( .A(n24642), .Z(n27119) );
  BUF_X1 U12263 ( .A(n24650), .Z(n27115) );
  BUF_X1 U12264 ( .A(n24650), .Z(n27116) );
  CLKBUF_X1 U12265 ( .A(n24651), .Z(n18918) );
  CLKBUF_X1 U12266 ( .A(n24651), .Z(n18919) );
  CLKBUF_X1 U12267 ( .A(n24652), .Z(n18920) );
  CLKBUF_X1 U12268 ( .A(n24652), .Z(n18921) );
  CLKBUF_X1 U12269 ( .A(n22955), .Z(n18922) );
  XNOR2_X1 U12270 ( .A(n4569), .B(n553), .ZN(n18923) );
  NAND2_X1 U12271 ( .A1(n27339), .A2(n27338), .ZN(n18924) );
  AND2_X1 U12272 ( .A1(n27297), .A2(n27299), .ZN(n18925) );
  NAND2_X1 U12273 ( .A1(n452), .A2(n24718), .ZN(n18926) );
  NAND2_X1 U12274 ( .A1(n27341), .A2(n27338), .ZN(n18927) );
  OR2_X1 U12275 ( .A1(n53950), .A2(n548), .ZN(n18928) );
  OR2_X1 U12276 ( .A1(n24717), .A2(n456), .ZN(n18929) );
  OR2_X1 U12277 ( .A1(n22953), .A2(n24718), .ZN(n18930) );
  NAND2_X1 U12278 ( .A1(n19175), .A2(n24721), .ZN(n18931) );
  OR2_X1 U12279 ( .A1(n25318), .A2(n4540), .ZN(n18932) );
  OR2_X1 U12280 ( .A1(n26948), .A2(n33000), .ZN(n18933) );
  OR2_X1 U12281 ( .A1(n20794), .A2(n43930), .ZN(n18934) );
  INV_X1 U12282 ( .A(n24697), .ZN(n278001) );
  NAND2_X1 U12283 ( .A1(n26082), .A2(n17265), .ZN(n18935) );
  NAND2_X1 U12284 ( .A1(n26501), .A2(n25314), .ZN(n18936) );
  NAND2_X1 U12285 ( .A1(n27808), .A2(n21517), .ZN(n18937) );
  OR2_X1 U12286 ( .A1(n21502), .A2(n20613), .ZN(n18938) );
  NAND2_X1 U12287 ( .A1(n27819), .A2(n21506), .ZN(n18939) );
  NAND2_X1 U12288 ( .A1(n27818), .A2(n22471), .ZN(n18940) );
  AND3_X1 U12289 ( .A1(n20892), .A2(n25665), .A3(n885), .ZN(n18941) );
  NAND4_X1 U12290 ( .A1(r924_LT_LE), .A2(n27806), .A3(n265301), .A4(n26515), 
        .ZN(n18942) );
  NAND4_X1 U12291 ( .A1(r948_LT_LE), .A2(n26081), .A3(n21869), .A4(n4417), 
        .ZN(n18943) );
  NAND4_X1 U12292 ( .A1(r929_LT_LE), .A2(n260901), .A3(n17114), .A4(n43920), 
        .ZN(n18944) );
  CLKBUF_X1 U12293 ( .A(n24728), .Z(n18945) );
  CLKBUF_X1 U12294 ( .A(n24699), .Z(n18946) );
  CLKBUF_X1 U12295 ( .A(n20543), .Z(n18947) );
  CLKBUF_X1 U12296 ( .A(n17097), .Z(n18948) );
  CLKBUF_X1 U12297 ( .A(n3135), .Z(n18949) );
  CLKBUF_X1 U12298 ( .A(n4170), .Z(n18950) );
  CLKBUF_X1 U12299 ( .A(n24758), .Z(n18951) );
  CLKBUF_X1 U12300 ( .A(n25196), .Z(n18952) );
  CLKBUF_X1 U12301 ( .A(n25193), .Z(n18953) );
  CLKBUF_X1 U12302 ( .A(n20607), .Z(n18954) );
  CLKBUF_X1 U12303 ( .A(n20608), .Z(n18955) );
  CLKBUF_X1 U12304 ( .A(n26961), .Z(n18956) );
  CLKBUF_X1 U12305 ( .A(n26964), .Z(n18957) );
  CLKBUF_X1 U12306 ( .A(n26963), .Z(n18958) );
  CLKBUF_X1 U12307 ( .A(n27781), .Z(n18959) );
  CLKBUF_X1 U12308 ( .A(n24825), .Z(n18960) );
  CLKBUF_X1 U12309 ( .A(n26953), .Z(n18961) );
  CLKBUF_X1 U12310 ( .A(n20627), .Z(n18962) );
  CLKBUF_X1 U12311 ( .A(n24829), .Z(n18963) );
  CLKBUF_X1 U12312 ( .A(n26954), .Z(n18964) );
  CLKBUF_X1 U12313 ( .A(n20643), .Z(n18965) );
  CLKBUF_X1 U12314 ( .A(n24834), .Z(n18966) );
  CLKBUF_X1 U12315 ( .A(n26955), .Z(n18967) );
  CLKBUF_X1 U12316 ( .A(n20651), .Z(n18968) );
  CLKBUF_X1 U12317 ( .A(n24838), .Z(n18969) );
  CLKBUF_X1 U12318 ( .A(n26956), .Z(n18970) );
  CLKBUF_X1 U12319 ( .A(n24842), .Z(n18971) );
  CLKBUF_X1 U12320 ( .A(n26957), .Z(n18972) );
  CLKBUF_X1 U12321 ( .A(n20660), .Z(n18973) );
  CLKBUF_X1 U12322 ( .A(n24846), .Z(n18974) );
  CLKBUF_X1 U12323 ( .A(n26958), .Z(n18975) );
  CLKBUF_X1 U12324 ( .A(n20675), .Z(n18976) );
  CLKBUF_X1 U12325 ( .A(n26959), .Z(n18977) );
  CLKBUF_X1 U12326 ( .A(n20683), .Z(n18978) );
  CLKBUF_X1 U12327 ( .A(n24854), .Z(n18979) );
  CLKBUF_X1 U12328 ( .A(n26960), .Z(n18980) );
  CLKBUF_X1 U12329 ( .A(n24864), .Z(n18981) );
  CLKBUF_X1 U12330 ( .A(n25249), .Z(n18982) );
  CLKBUF_X1 U12331 ( .A(n24864), .Z(n18983) );
  CLKBUF_X1 U12332 ( .A(n26946), .Z(n18984) );
  CLKBUF_X1 U12333 ( .A(n36250), .Z(n18985) );
  CLKBUF_X1 U12334 ( .A(n32110), .Z(n18986) );
  CLKBUF_X1 U12335 ( .A(n26945), .Z(n18987) );
  CLKBUF_X1 U12336 ( .A(n20582), .Z(n18988) );
  CLKBUF_X1 U12337 ( .A(n20578), .Z(n18989) );
  CLKBUF_X1 U12338 ( .A(n24169), .Z(n18990) );
  CLKBUF_X1 U12339 ( .A(n24136), .Z(n18991) );
  CLKBUF_X1 U12340 ( .A(n24124), .Z(n18992) );
  CLKBUF_X1 U12341 ( .A(n24130), .Z(n18993) );
  CLKBUF_X1 U12342 ( .A(n24118), .Z(n18994) );
  CLKBUF_X1 U12343 ( .A(n24123), .Z(n18995) );
  CLKBUF_X1 U12344 ( .A(n24111), .Z(n18996) );
  CLKBUF_X1 U12345 ( .A(n24117), .Z(n18997) );
  CLKBUF_X1 U12346 ( .A(n24105), .Z(n18998) );
  CLKBUF_X1 U12347 ( .A(n24112), .Z(n18999) );
  CLKBUF_X1 U12348 ( .A(n24080), .Z(n19000) );
  CLKBUF_X1 U12349 ( .A(n26975), .Z(n19001) );
  CLKBUF_X1 U12350 ( .A(n20683), .Z(n19002) );
  CLKBUF_X1 U12351 ( .A(n24854), .Z(n19003) );
  CLKBUF_X1 U12352 ( .A(n24850), .Z(n19004) );
  CLKBUF_X1 U12353 ( .A(n20675), .Z(n19005) );
  CLKBUF_X1 U12354 ( .A(n24846), .Z(n19006) );
  CLKBUF_X1 U12355 ( .A(n20667), .Z(n19007) );
  CLKBUF_X1 U12356 ( .A(n20659), .Z(n19008) );
  CLKBUF_X1 U12357 ( .A(n24842), .Z(n19009) );
  CLKBUF_X1 U12358 ( .A(n20651), .Z(n19010) );
  CLKBUF_X1 U12359 ( .A(n24838), .Z(n19011) );
  CLKBUF_X1 U12360 ( .A(n24834), .Z(n19012) );
  CLKBUF_X1 U12361 ( .A(n20643), .Z(n19013) );
  CLKBUF_X1 U12362 ( .A(n24829), .Z(n19014) );
  CLKBUF_X1 U12363 ( .A(n20634), .Z(n19015) );
  CLKBUF_X1 U12364 ( .A(n26997), .Z(n19016) );
  NAND2_X1 U12365 ( .A1(n278101), .A2(n21518), .ZN(n19017) );
  NAND2_X1 U12366 ( .A1(n26499), .A2(n19267), .ZN(n19018) );
  NAND2_X1 U12367 ( .A1(n27814), .A2(n21518), .ZN(n19019) );
  CLKBUF_X1 U12368 ( .A(n27230), .Z(n19020) );
  CLKBUF_X1 U12369 ( .A(n20910), .Z(n19021) );
  CLKBUF_X1 U12370 ( .A(n27175), .Z(n19022) );
  CLKBUF_X1 U12371 ( .A(n27231), .Z(n19023) );
  CLKBUF_X1 U12372 ( .A(n20495), .Z(n19024) );
  CLKBUF_X1 U12373 ( .A(n20914), .Z(n19025) );
  CLKBUF_X1 U12374 ( .A(n27176), .Z(n19026) );
  CLKBUF_X1 U12375 ( .A(n18101), .Z(n19027) );
  CLKBUF_X1 U12376 ( .A(n20497), .Z(n19028) );
  CLKBUF_X1 U12377 ( .A(n20918), .Z(n19029) );
  CLKBUF_X1 U12378 ( .A(n18277), .Z(n19030) );
  CLKBUF_X1 U12379 ( .A(n18102), .Z(n19031) );
  CLKBUF_X1 U12380 ( .A(n20923), .Z(n19032) );
  CLKBUF_X1 U12381 ( .A(n18104), .Z(n19033) );
  CLKBUF_X1 U12382 ( .A(n18106), .Z(n19034) );
  CLKBUF_X1 U12383 ( .A(n18107), .Z(n19035) );
  CLKBUF_X1 U12384 ( .A(n18108), .Z(n19036) );
  CLKBUF_X1 U12385 ( .A(n18109), .Z(n19037) );
  CLKBUF_X1 U12386 ( .A(n18110), .Z(n19038) );
  CLKBUF_X1 U12387 ( .A(n18111), .Z(n19039) );
  CLKBUF_X1 U12388 ( .A(n18112), .Z(n19040) );
  CLKBUF_X1 U12389 ( .A(n18113), .Z(n19041) );
  CLKBUF_X1 U12390 ( .A(n20942), .Z(n19042) );
  CLKBUF_X1 U12391 ( .A(n18114), .Z(n19043) );
  CLKBUF_X1 U12392 ( .A(n18115), .Z(n19044) );
  CLKBUF_X1 U12393 ( .A(n20952), .Z(n19045) );
  CLKBUF_X1 U12394 ( .A(n18116), .Z(n19046) );
  CLKBUF_X1 U12395 ( .A(n18117), .Z(n19047) );
  CLKBUF_X1 U12396 ( .A(n18118), .Z(n19048) );
  CLKBUF_X1 U12397 ( .A(n18119), .Z(n19049) );
  CLKBUF_X1 U12398 ( .A(n18120), .Z(n19050) );
  CLKBUF_X1 U12399 ( .A(n18121), .Z(n19051) );
  CLKBUF_X1 U12400 ( .A(n18123), .Z(n19052) );
  CLKBUF_X1 U12401 ( .A(n20963), .Z(n19053) );
  CLKBUF_X1 U12402 ( .A(n20965), .Z(n19054) );
  CLKBUF_X1 U12403 ( .A(n18127), .Z(n19055) );
  CLKBUF_X1 U12404 ( .A(n18128), .Z(n19056) );
  CLKBUF_X1 U12405 ( .A(n18129), .Z(n19057) );
  CLKBUF_X1 U12406 ( .A(n18130), .Z(n19058) );
  CLKBUF_X1 U12407 ( .A(n18131), .Z(n19059) );
  CLKBUF_X1 U12408 ( .A(n18132), .Z(n19060) );
  CLKBUF_X1 U12409 ( .A(n18133), .Z(n19061) );
  CLKBUF_X1 U12410 ( .A(n18134), .Z(n19062) );
  CLKBUF_X1 U12411 ( .A(n18135), .Z(n19063) );
  CLKBUF_X1 U12412 ( .A(n20998), .Z(n19064) );
  CLKBUF_X1 U12413 ( .A(n18137), .Z(n19065) );
  CLKBUF_X1 U12414 ( .A(n21005), .Z(n19066) );
  CLKBUF_X1 U12415 ( .A(n18139), .Z(n19067) );
  CLKBUF_X1 U12416 ( .A(n18140), .Z(n19068) );
  CLKBUF_X1 U12417 ( .A(n18141), .Z(n19069) );
  INV_X1 U12418 ( .A(n24434), .ZN(n26950) );
  CLKBUF_X1 U12419 ( .A(n18142), .Z(n19070) );
  CLKBUF_X1 U12420 ( .A(n18143), .Z(n19071) );
  CLKBUF_X1 U12421 ( .A(n24179), .Z(n19072) );
  CLKBUF_X1 U12422 ( .A(n18144), .Z(n19073) );
  CLKBUF_X1 U12423 ( .A(n18145), .Z(n19074) );
  CLKBUF_X1 U12424 ( .A(n24174), .Z(n19075) );
  CLKBUF_X1 U12425 ( .A(n18146), .Z(n19076) );
  CLKBUF_X1 U12426 ( .A(n18147), .Z(n19077) );
  CLKBUF_X1 U12427 ( .A(n18148), .Z(n19078) );
  CLKBUF_X1 U12428 ( .A(n18150), .Z(n19079) );
  CLKBUF_X1 U12429 ( .A(n18151), .Z(n19080) );
  CLKBUF_X1 U12430 ( .A(n18152), .Z(n19081) );
  CLKBUF_X1 U12431 ( .A(n21029), .Z(n19082) );
  CLKBUF_X1 U12432 ( .A(n21031), .Z(n19083) );
  CLKBUF_X1 U12433 ( .A(n18153), .Z(n19084) );
  CLKBUF_X1 U12434 ( .A(n21034), .Z(n19085) );
  CLKBUF_X1 U12435 ( .A(n21036), .Z(n19086) );
  CLKBUF_X1 U12436 ( .A(n21038), .Z(n19087) );
  CLKBUF_X1 U12437 ( .A(n18154), .Z(n19088) );
  CLKBUF_X1 U12438 ( .A(n21041), .Z(n19089) );
  CLKBUF_X1 U12439 ( .A(n21043), .Z(n19090) );
  CLKBUF_X1 U12440 ( .A(n21045), .Z(n19091) );
  CLKBUF_X1 U12441 ( .A(n21047), .Z(n19092) );
  CLKBUF_X1 U12442 ( .A(n18155), .Z(n19093) );
  CLKBUF_X1 U12443 ( .A(n18156), .Z(n19094) );
  CLKBUF_X1 U12444 ( .A(n18157), .Z(n19095) );
  CLKBUF_X1 U12445 ( .A(n18158), .Z(n19096) );
  CLKBUF_X1 U12446 ( .A(n18159), .Z(n19097) );
  CLKBUF_X1 U12447 ( .A(n18160), .Z(n19098) );
  CLKBUF_X1 U12448 ( .A(n18161), .Z(n19099) );
  CLKBUF_X1 U12449 ( .A(n18162), .Z(n19100) );
  CLKBUF_X1 U12450 ( .A(n18164), .Z(n19101) );
  CLKBUF_X1 U12451 ( .A(n18165), .Z(n19102) );
  CLKBUF_X1 U12452 ( .A(n22686), .Z(n19103) );
  CLKBUF_X1 U12453 ( .A(n18168), .Z(n19104) );
  CLKBUF_X1 U12454 ( .A(n18169), .Z(n19105) );
  CLKBUF_X1 U12455 ( .A(n18170), .Z(n19106) );
  CLKBUF_X1 U12456 ( .A(n18171), .Z(n19107) );
  CLKBUF_X1 U12457 ( .A(n4571), .Z(n19108) );
  CLKBUF_X1 U12458 ( .A(n54220), .Z(n19109) );
  CLKBUF_X1 U12459 ( .A(n3104), .Z(n19110) );
  CLKBUF_X1 U12460 ( .A(n3072), .Z(n19111) );
  CLKBUF_X1 U12461 ( .A(n3154), .Z(n19112) );
  CLKBUF_X1 U12462 ( .A(n31290), .Z(n19113) );
  CLKBUF_X1 U12463 ( .A(n32040), .Z(n19114) );
  CLKBUF_X1 U12464 ( .A(n3179), .Z(n19115) );
  CLKBUF_X1 U12465 ( .A(n32540), .Z(n19116) );
  CLKBUF_X1 U12466 ( .A(n3229), .Z(n19117) );
  CLKBUF_X1 U12467 ( .A(n33030), .Z(n19118) );
  CLKBUF_X1 U12468 ( .A(n3278), .Z(n19119) );
  CLKBUF_X1 U12469 ( .A(n3347), .Z(n19120) );
  CLKBUF_X1 U12470 ( .A(n3325), .Z(n19121) );
  CLKBUF_X1 U12471 ( .A(n3391), .Z(n19122) );
  CLKBUF_X1 U12472 ( .A(n33690), .Z(n19123) );
  CLKBUF_X1 U12473 ( .A(n3436), .Z(n19124) );
  CLKBUF_X1 U12474 ( .A(n3413), .Z(n19125) );
  CLKBUF_X1 U12475 ( .A(n3485), .Z(n19126) );
  CLKBUF_X1 U12476 ( .A(n34600), .Z(n19127) );
  CLKBUF_X1 U12477 ( .A(n3529), .Z(n19128) );
  CLKBUF_X1 U12478 ( .A(n35070), .Z(n19129) );
  CLKBUF_X1 U12479 ( .A(n3573), .Z(n19130) );
  CLKBUF_X1 U12480 ( .A(n35510), .Z(n19131) );
  CLKBUF_X1 U12481 ( .A(n3618), .Z(n19132) );
  CLKBUF_X1 U12482 ( .A(n35950), .Z(n19133) );
  CLKBUF_X1 U12483 ( .A(n3666), .Z(n19134) );
  CLKBUF_X1 U12484 ( .A(n3642), .Z(n19135) );
  CLKBUF_X1 U12485 ( .A(n37100), .Z(n19136) );
  CLKBUF_X1 U12486 ( .A(n3688), .Z(n19137) );
  CLKBUF_X1 U12487 ( .A(n3754), .Z(n19138) );
  CLKBUF_X1 U12488 ( .A(n3732), .Z(n19139) );
  CLKBUF_X1 U12489 ( .A(n37990), .Z(n19140) );
  CLKBUF_X1 U12490 ( .A(n3776), .Z(n19141) );
  CLKBUF_X1 U12491 ( .A(n38480), .Z(n19142) );
  CLKBUF_X1 U12492 ( .A(n3823), .Z(n19143) );
  CLKBUF_X1 U12493 ( .A(n3892), .Z(n19144) );
  CLKBUF_X1 U12494 ( .A(n3870), .Z(n19145) );
  CLKBUF_X1 U12495 ( .A(n39360), .Z(n19146) );
  CLKBUF_X1 U12496 ( .A(n3914), .Z(n19147) );
  CLKBUF_X1 U12497 ( .A(n3981), .Z(n19148) );
  CLKBUF_X1 U12498 ( .A(n3958), .Z(n19149) );
  CLKBUF_X1 U12499 ( .A(n4031), .Z(n19150) );
  CLKBUF_X1 U12500 ( .A(n4005), .Z(n19151) );
  CLKBUF_X1 U12501 ( .A(n4075), .Z(n19152) );
  CLKBUF_X1 U12502 ( .A(n40530), .Z(n19153) );
  CLKBUF_X1 U12503 ( .A(n4119), .Z(n19154) );
  CLKBUF_X1 U12504 ( .A(n40970), .Z(n19155) );
  CLKBUF_X1 U12505 ( .A(n4164), .Z(n19156) );
  CLKBUF_X1 U12506 ( .A(n41410), .Z(n19157) );
  CLKBUF_X1 U12507 ( .A(n42140), .Z(n19158) );
  CLKBUF_X1 U12508 ( .A(n41880), .Z(n19159) );
  CLKBUF_X1 U12509 ( .A(n4258), .Z(n19160) );
  CLKBUF_X1 U12510 ( .A(n4236), .Z(n19161) );
  CLKBUF_X1 U12511 ( .A(n43020), .Z(n19162) );
  CLKBUF_X1 U12512 ( .A(n4280), .Z(n19163) );
  CLKBUF_X1 U12513 ( .A(n43470), .Z(n19164) );
  CLKBUF_X1 U12514 ( .A(n4324), .Z(n19165) );
  CLKBUF_X1 U12515 ( .A(n4396), .Z(n19166) );
  CLKBUF_X1 U12516 ( .A(n4371), .Z(n19167) );
  CLKBUF_X1 U12517 ( .A(n44450), .Z(n19168) );
  CLKBUF_X1 U12518 ( .A(n4421), .Z(n19169) );
  CLKBUF_X1 U12519 ( .A(n4494), .Z(n19170) );
  CLKBUF_X1 U12520 ( .A(n44700), .Z(n19171) );
  CLKBUF_X1 U12521 ( .A(n4543), .Z(n19172) );
  CLKBUF_X1 U12522 ( .A(n45180), .Z(n19173) );
  CLKBUF_X1 U12523 ( .A(n4419), .Z(n19174) );
  CLKBUF_X1 U12524 ( .A(n21135), .Z(n19175) );
  CLKBUF_X1 U12525 ( .A(n18172), .Z(n19176) );
  CLKBUF_X1 U12526 ( .A(n21138), .Z(n19177) );
  CLKBUF_X1 U12527 ( .A(n21142), .Z(n19178) );
  CLKBUF_X1 U12528 ( .A(n18175), .Z(n19179) );
  CLKBUF_X1 U12529 ( .A(n18177), .Z(n19180) );
  CLKBUF_X1 U12530 ( .A(n18179), .Z(n19181) );
  CLKBUF_X1 U12531 ( .A(n18181), .Z(n19182) );
  CLKBUF_X1 U12532 ( .A(n21338), .Z(n19183) );
  CLKBUF_X1 U12533 ( .A(n18186), .Z(n19184) );
  CLKBUF_X1 U12534 ( .A(n20491), .Z(n19185) );
  CLKBUF_X1 U12535 ( .A(n18189), .Z(n19186) );
  CLKBUF_X1 U12536 ( .A(n18191), .Z(n19187) );
  CLKBUF_X1 U12537 ( .A(n18193), .Z(n19188) );
  CLKBUF_X1 U12538 ( .A(n24616), .Z(n19189) );
  CLKBUF_X1 U12539 ( .A(n18195), .Z(n19190) );
  CLKBUF_X1 U12540 ( .A(n18197), .Z(n19191) );
  CLKBUF_X1 U12541 ( .A(n18199), .Z(n19192) );
  CLKBUF_X1 U12542 ( .A(n21209), .Z(n19193) );
  CLKBUF_X1 U12543 ( .A(n21213), .Z(n19194) );
  CLKBUF_X1 U12544 ( .A(n18203), .Z(n19195) );
  CLKBUF_X1 U12545 ( .A(n18205), .Z(n19196) );
  CLKBUF_X1 U12546 ( .A(n18207), .Z(n19197) );
  CLKBUF_X1 U12547 ( .A(n20483), .Z(n19198) );
  CLKBUF_X1 U12548 ( .A(n18210), .Z(n19199) );
  CLKBUF_X1 U12549 ( .A(n27047), .Z(n19200) );
  CLKBUF_X1 U12550 ( .A(n21234), .Z(n19201) );
  CLKBUF_X1 U12551 ( .A(n20486), .Z(n19202) );
  CLKBUF_X1 U12552 ( .A(n18213), .Z(n19203) );
  CLKBUF_X1 U12553 ( .A(n18215), .Z(n19204) );
  CLKBUF_X1 U12554 ( .A(n18217), .Z(n19205) );
  CLKBUF_X1 U12555 ( .A(n18220), .Z(n19206) );
  CLKBUF_X1 U12556 ( .A(n18222), .Z(n19207) );
  CLKBUF_X1 U12557 ( .A(n20479), .Z(n19208) );
  CLKBUF_X1 U12558 ( .A(n18225), .Z(n19209) );
  CLKBUF_X1 U12559 ( .A(n18228), .Z(n19210) );
  CLKBUF_X1 U12560 ( .A(n18230), .Z(n19211) );
  CLKBUF_X1 U12561 ( .A(n18232), .Z(n19212) );
  BUF_X1 U12562 ( .A(n24603), .Z(n26976) );
  CLKBUF_X1 U12563 ( .A(n21284), .Z(n19213) );
  CLKBUF_X1 U12564 ( .A(n21288), .Z(n19214) );
  CLKBUF_X1 U12565 ( .A(n18236), .Z(n19215) );
  CLKBUF_X1 U12566 ( .A(n18238), .Z(n19216) );
  CLKBUF_X1 U12567 ( .A(n18240), .Z(n19217) );
  CLKBUF_X1 U12568 ( .A(n18242), .Z(n19218) );
  CLKBUF_X1 U12569 ( .A(n18244), .Z(n19219) );
  CLKBUF_X1 U12570 ( .A(n18246), .Z(n19220) );
  CLKBUF_X1 U12571 ( .A(n18248), .Z(n19221) );
  CLKBUF_X1 U12572 ( .A(n18250), .Z(n19222) );
  CLKBUF_X1 U12573 ( .A(n18252), .Z(n19223) );
  CLKBUF_X1 U12574 ( .A(n18254), .Z(n19224) );
  CLKBUF_X1 U12575 ( .A(n18256), .Z(n19225) );
  CLKBUF_X1 U12576 ( .A(n3186), .Z(n19226) );
  CLKBUF_X1 U12577 ( .A(n21328), .Z(n19227) );
  CLKBUF_X1 U12578 ( .A(n18259), .Z(n19228) );
  CLKBUF_X1 U12579 ( .A(n38060), .Z(n19229) );
  CLKBUF_X1 U12580 ( .A(n18261), .Z(n19230) );
  CLKBUF_X1 U12581 ( .A(n18264), .Z(n19231) );
  CLKBUF_X1 U12582 ( .A(n18266), .Z(n19232) );
  CLKBUF_X1 U12583 ( .A(n21352), .Z(n19233) );
  CLKBUF_X1 U12584 ( .A(n18269), .Z(n19234) );
  CLKBUF_X1 U12585 ( .A(n4170), .Z(n19235) );
  CLKBUF_X1 U12586 ( .A(n3135), .Z(n19236) );
  CLKBUF_X1 U12587 ( .A(n21373), .Z(n19237) );
  CLKBUF_X1 U12588 ( .A(n21379), .Z(n19238) );
  CLKBUF_X1 U12589 ( .A(n21383), .Z(n19239) );
  CLKBUF_X1 U12590 ( .A(n18275), .Z(n19240) );
  CLKBUF_X1 U12591 ( .A(n17133), .Z(n19241) );
  CLKBUF_X1 U12592 ( .A(n18278), .Z(n19242) );
  CLKBUF_X1 U12593 ( .A(n18279), .Z(n19243) );
  CLKBUF_X1 U12594 ( .A(n18281), .Z(n19244) );
  CLKBUF_X1 U12595 ( .A(n21421), .Z(n19245) );
  CLKBUF_X1 U12596 ( .A(n21428), .Z(n19246) );
  CLKBUF_X1 U12597 ( .A(n18987), .Z(n19247) );
  CLKBUF_X1 U12598 ( .A(n18061), .Z(n19248) );
  CLKBUF_X1 U12599 ( .A(n18062), .Z(n19249) );
  CLKBUF_X1 U12600 ( .A(n25100), .Z(n19250) );
  CLKBUF_X1 U12601 ( .A(n25106), .Z(n19251) );
  CLKBUF_X1 U12602 ( .A(n18053), .Z(n19252) );
  CLKBUF_X1 U12603 ( .A(n18054), .Z(n19253) );
  CLKBUF_X1 U12604 ( .A(n18057), .Z(n19254) );
  CLKBUF_X1 U12605 ( .A(n18056), .Z(n19255) );
  CLKBUF_X1 U12606 ( .A(n18058), .Z(n19256) );
  CLKBUF_X1 U12607 ( .A(n18060), .Z(n19257) );
  CLKBUF_X1 U12608 ( .A(n18048), .Z(n19258) );
  CLKBUF_X1 U12609 ( .A(n18047), .Z(n19259) );
  CLKBUF_X1 U12610 ( .A(n18050), .Z(n19260) );
  CLKBUF_X1 U12611 ( .A(n18049), .Z(n19261) );
  CLKBUF_X1 U12612 ( .A(n20700), .Z(n19262) );
  CLKBUF_X1 U12613 ( .A(n20704), .Z(n19263) );
  CLKBUF_X1 U12614 ( .A(n18051), .Z(n19264) );
  CLKBUF_X1 U12615 ( .A(n18052), .Z(n19265) );
  CLKBUF_X1 U12616 ( .A(n19752), .Z(n19266) );
  BUF_X1 U12617 ( .A(n24644), .Z(n27122) );
  BUF_X1 U12618 ( .A(n24647), .Z(n27113) );
  BUF_X1 U12619 ( .A(n24648), .Z(n27114) );
  BUF_X1 U12620 ( .A(n24644), .Z(n27121) );
  CLKBUF_X1 U12621 ( .A(n23657), .Z(n19267) );
  CLKBUF_X1 U12622 ( .A(n18705), .Z(n19268) );
  CLKBUF_X1 U12623 ( .A(n18706), .Z(n19269) );
  CLKBUF_X1 U12624 ( .A(n25250), .Z(n19270) );
  CLKBUF_X1 U12625 ( .A(n18721), .Z(n19271) );
  CLKBUF_X1 U12626 ( .A(n18087), .Z(n19272) );
  CLKBUF_X1 U12627 ( .A(n18455), .Z(n19273) );
  CLKBUF_X1 U12628 ( .A(n18456), .Z(n19274) );
  CLKBUF_X1 U12629 ( .A(n18458), .Z(n19275) );
  CLKBUF_X1 U12630 ( .A(n18459), .Z(n19276) );
  CLKBUF_X1 U12631 ( .A(n18460), .Z(n19277) );
  CLKBUF_X1 U12632 ( .A(n18461), .Z(n19278) );
  CLKBUF_X1 U12633 ( .A(n22695), .Z(n19279) );
  CLKBUF_X1 U12634 ( .A(n22699), .Z(n19280) );
  CLKBUF_X1 U12635 ( .A(n18464), .Z(n19281) );
  CLKBUF_X1 U12636 ( .A(n18466), .Z(n19282) );
  CLKBUF_X1 U12637 ( .A(n22709), .Z(n19283) );
  CLKBUF_X1 U12638 ( .A(n18469), .Z(n19284) );
  CLKBUF_X1 U12639 ( .A(n18471), .Z(n19285) );
  CLKBUF_X1 U12640 ( .A(n18473), .Z(n19286) );
  CLKBUF_X1 U12641 ( .A(n18475), .Z(n19287) );
  CLKBUF_X1 U12642 ( .A(n18477), .Z(n19288) );
  CLKBUF_X1 U12643 ( .A(n18478), .Z(n19289) );
  CLKBUF_X1 U12644 ( .A(n18480), .Z(n19290) );
  CLKBUF_X1 U12645 ( .A(n22736), .Z(n19291) );
  CLKBUF_X1 U12646 ( .A(n22741), .Z(n19292) );
  CLKBUF_X1 U12647 ( .A(n22746), .Z(n19293) );
  CLKBUF_X1 U12648 ( .A(n22750), .Z(n19294) );
  CLKBUF_X1 U12649 ( .A(n18483), .Z(n19295) );
  CLKBUF_X1 U12650 ( .A(n18484), .Z(n19296) );
  CLKBUF_X1 U12651 ( .A(n18485), .Z(n19297) );
  CLKBUF_X1 U12652 ( .A(n22778), .Z(n19298) );
  CLKBUF_X1 U12653 ( .A(n22780), .Z(n19299) );
  CLKBUF_X1 U12654 ( .A(n22782), .Z(n19300) );
  CLKBUF_X1 U12655 ( .A(n22784), .Z(n19301) );
  CLKBUF_X1 U12656 ( .A(n22788), .Z(n19302) );
  CLKBUF_X1 U12657 ( .A(n18491), .Z(n19303) );
  CLKBUF_X1 U12658 ( .A(n22807), .Z(n19304) );
  CLKBUF_X1 U12659 ( .A(n22809), .Z(n19305) );
  CLKBUF_X1 U12660 ( .A(n18063), .Z(n19306) );
  CLKBUF_X1 U12661 ( .A(n20716), .Z(n19307) );
  CLKBUF_X1 U12662 ( .A(n18059), .Z(n19308) );
  CLKBUF_X1 U12663 ( .A(n20714), .Z(n19309) );
  CLKBUF_X1 U12664 ( .A(n18055), .Z(n19310) );
  CLKBUF_X1 U12665 ( .A(n20702), .Z(n19311) );
  CLKBUF_X1 U12666 ( .A(n18034), .Z(n19312) );
  CLKBUF_X1 U12667 ( .A(n20555), .Z(n19313) );
  CLKBUF_X1 U12668 ( .A(n22810), .Z(n19314) );
  CLKBUF_X1 U12669 ( .A(n22808), .Z(n19315) );
  CLKBUF_X1 U12670 ( .A(n18002), .Z(n19316) );
  CLKBUF_X1 U12671 ( .A(n18001), .Z(n19317) );
  CLKBUF_X1 U12672 ( .A(n19757), .Z(n19318) );
  OAI21_X1 U12673 ( .B1(n27294), .B2(n27301), .A(n27306), .ZN(r899_B_3_) );
  CLKBUF_X1 U12674 ( .A(n20897), .Z(n19319) );
  CLKBUF_X1 U12675 ( .A(n20898), .Z(n19320) );
  CLKBUF_X1 U12676 ( .A(n22967), .Z(n19321) );
  CLKBUF_X1 U12677 ( .A(n20893), .Z(n19322) );
  CLKBUF_X1 U12678 ( .A(n20894), .Z(n19323) );
  CLKBUF_X1 U12679 ( .A(n22970), .Z(n19324) );
  INV_X1 U12680 ( .A(n28670), .ZN(n19325) );
  INV_X1 U12681 ( .A(n2750), .ZN(n19326) );
  INV_X1 U12682 ( .A(n1859), .ZN(n19327) );
  INV_X1 U12683 ( .A(n2882), .ZN(n19328) );
  INV_X1 U12684 ( .A(n278000), .ZN(n19329) );
  INV_X1 U12685 ( .A(n2765), .ZN(n19330) );
  INV_X1 U12686 ( .A(n2720), .ZN(n19331) );
  INV_X1 U12687 ( .A(n264800), .ZN(n19332) );
  INV_X1 U12688 ( .A(n2633), .ZN(n19333) );
  INV_X1 U12689 ( .A(n2618), .ZN(n19334) );
  INV_X1 U12690 ( .A(n260300), .ZN(n19335) );
  INV_X1 U12691 ( .A(n2552), .ZN(n19336) );
  INV_X1 U12692 ( .A(n2537), .ZN(n19337) );
  INV_X1 U12693 ( .A(n2522), .ZN(n19338) );
  INV_X1 U12694 ( .A(n2507), .ZN(n19339) );
  INV_X1 U12695 ( .A(n2492), .ZN(n19340) );
  INV_X1 U12696 ( .A(n2477), .ZN(n19341) );
  INV_X1 U12697 ( .A(n2426), .ZN(n19342) );
  INV_X1 U12698 ( .A(n2411), .ZN(n19343) );
  INV_X1 U12699 ( .A(n2396), .ZN(n19344) );
  INV_X1 U12700 ( .A(n2381), .ZN(n19345) );
  INV_X1 U12701 ( .A(n2366), .ZN(n19346) );
  INV_X1 U12702 ( .A(n2351), .ZN(n19347) );
  INV_X1 U12703 ( .A(n2336), .ZN(n19348) );
  INV_X1 U12704 ( .A(n2285), .ZN(n19349) );
  INV_X1 U12705 ( .A(n2270), .ZN(n19350) );
  INV_X1 U12706 ( .A(n2255), .ZN(n19351) );
  INV_X1 U12707 ( .A(n2204), .ZN(n19352) );
  INV_X1 U12708 ( .A(n2189), .ZN(n19353) );
  INV_X1 U12709 ( .A(n2174), .ZN(n19354) );
  INV_X1 U12710 ( .A(n2159), .ZN(n19355) );
  INV_X1 U12711 ( .A(n2144), .ZN(n19356) );
  INV_X1 U12712 ( .A(n2129), .ZN(n19357) );
  INV_X1 U12713 ( .A(n2114), .ZN(n19358) );
  INV_X1 U12714 ( .A(n2099), .ZN(n19359) );
  INV_X1 U12715 ( .A(n2000), .ZN(n19360) );
  INV_X1 U12716 ( .A(n1985), .ZN(n19361) );
  INV_X1 U12717 ( .A(n1955), .ZN(n19362) );
  INV_X1 U12718 ( .A(n1919), .ZN(n19363) );
  INV_X1 U12719 ( .A(n1904), .ZN(n19364) );
  INV_X1 U12720 ( .A(n1889), .ZN(n19365) );
  INV_X1 U12721 ( .A(n1874), .ZN(n19366) );
  INV_X1 U12722 ( .A(weight_queue_7__7__0_), .ZN(n19367) );
  INV_X1 U12723 ( .A(n19367), .ZN(n19368) );
  INV_X1 U12724 ( .A(n17137), .ZN(n19369) );
  INV_X1 U12725 ( .A(weight_queue_7__7__1_), .ZN(n19370) );
  INV_X1 U12726 ( .A(n19370), .ZN(n19371) );
  INV_X1 U12727 ( .A(n17138), .ZN(n19372) );
  INV_X1 U12728 ( .A(weight_queue_7__7__2_), .ZN(n19373) );
  INV_X1 U12729 ( .A(n19373), .ZN(n19374) );
  INV_X1 U12730 ( .A(n17139), .ZN(n19375) );
  INV_X1 U12731 ( .A(weight_queue_7__7__3_), .ZN(n19376) );
  INV_X1 U12732 ( .A(n19376), .ZN(n19377) );
  INV_X1 U12733 ( .A(n17140), .ZN(n19378) );
  INV_X1 U12734 ( .A(weight_queue_7__7__4_), .ZN(n19379) );
  INV_X1 U12735 ( .A(n19379), .ZN(n19380) );
  INV_X1 U12736 ( .A(n17141), .ZN(n19381) );
  INV_X1 U12737 ( .A(weight_queue_7__7__5_), .ZN(n19382) );
  INV_X1 U12738 ( .A(n19382), .ZN(n19383) );
  INV_X1 U12739 ( .A(n17142), .ZN(n19384) );
  INV_X1 U12740 ( .A(weight_queue_7__7__6_), .ZN(n19385) );
  INV_X1 U12741 ( .A(n19385), .ZN(n19386) );
  INV_X1 U12742 ( .A(n17143), .ZN(n19387) );
  INV_X1 U12743 ( .A(weight_queue_7__7__7_), .ZN(n19388) );
  INV_X1 U12744 ( .A(n17144), .ZN(n19389) );
  INV_X1 U12745 ( .A(n19388), .ZN(n19390) );
  INV_X1 U12746 ( .A(weight_queue_7__6__0_), .ZN(n19391) );
  INV_X1 U12747 ( .A(n19391), .ZN(n19392) );
  INV_X1 U12748 ( .A(n17145), .ZN(n19393) );
  INV_X1 U12749 ( .A(weight_queue_7__6__1_), .ZN(n19394) );
  INV_X1 U12750 ( .A(n19394), .ZN(n19395) );
  INV_X1 U12751 ( .A(n17146), .ZN(n19396) );
  INV_X1 U12752 ( .A(weight_queue_7__6__2_), .ZN(n19397) );
  INV_X1 U12753 ( .A(n19397), .ZN(n19398) );
  INV_X1 U12754 ( .A(n17147), .ZN(n19399) );
  INV_X1 U12755 ( .A(weight_queue_7__6__3_), .ZN(n19400) );
  INV_X1 U12756 ( .A(n19400), .ZN(n19401) );
  INV_X1 U12757 ( .A(n17148), .ZN(n19402) );
  INV_X1 U12758 ( .A(weight_queue_7__6__4_), .ZN(n19403) );
  INV_X1 U12759 ( .A(n19403), .ZN(n19404) );
  INV_X1 U12760 ( .A(n17149), .ZN(n19405) );
  INV_X1 U12761 ( .A(weight_queue_7__6__5_), .ZN(n19406) );
  INV_X1 U12762 ( .A(n19406), .ZN(n19407) );
  INV_X1 U12763 ( .A(n17150), .ZN(n19408) );
  INV_X1 U12764 ( .A(weight_queue_7__6__6_), .ZN(n19409) );
  INV_X1 U12765 ( .A(n19409), .ZN(n19410) );
  INV_X1 U12766 ( .A(n17151), .ZN(n19411) );
  INV_X1 U12767 ( .A(weight_queue_7__6__7_), .ZN(n19412) );
  INV_X1 U12768 ( .A(n17152), .ZN(n19413) );
  INV_X1 U12769 ( .A(n19412), .ZN(n19414) );
  INV_X1 U12770 ( .A(weight_queue_7__5__0_), .ZN(n19415) );
  INV_X1 U12771 ( .A(n19415), .ZN(n19416) );
  INV_X1 U12772 ( .A(n17153), .ZN(n19417) );
  INV_X1 U12773 ( .A(weight_queue_7__5__1_), .ZN(n19418) );
  INV_X1 U12774 ( .A(n19418), .ZN(n19419) );
  INV_X1 U12775 ( .A(n17154), .ZN(n19420) );
  INV_X1 U12776 ( .A(weight_queue_7__5__2_), .ZN(n19421) );
  INV_X1 U12777 ( .A(n19421), .ZN(n19422) );
  INV_X1 U12778 ( .A(n17155), .ZN(n19423) );
  INV_X1 U12779 ( .A(weight_queue_7__5__3_), .ZN(n19424) );
  INV_X1 U12780 ( .A(n19424), .ZN(n19425) );
  INV_X1 U12781 ( .A(n17156), .ZN(n19426) );
  INV_X1 U12782 ( .A(weight_queue_7__5__4_), .ZN(n19427) );
  INV_X1 U12783 ( .A(n19427), .ZN(n19428) );
  INV_X1 U12784 ( .A(n17157), .ZN(n19429) );
  INV_X1 U12785 ( .A(weight_queue_7__5__5_), .ZN(n19430) );
  INV_X1 U12786 ( .A(n19430), .ZN(n19431) );
  INV_X1 U12787 ( .A(n17158), .ZN(n19432) );
  INV_X1 U12788 ( .A(weight_queue_7__5__6_), .ZN(n19433) );
  INV_X1 U12789 ( .A(n19433), .ZN(n19434) );
  INV_X1 U12790 ( .A(n17159), .ZN(n19435) );
  INV_X1 U12791 ( .A(weight_queue_7__5__7_), .ZN(n19436) );
  INV_X1 U12792 ( .A(n17160), .ZN(n19437) );
  INV_X1 U12793 ( .A(n19436), .ZN(n19438) );
  INV_X1 U12794 ( .A(weight_queue_7__4__0_), .ZN(n19439) );
  INV_X1 U12795 ( .A(n19439), .ZN(n19440) );
  INV_X1 U12796 ( .A(n17161), .ZN(n19441) );
  INV_X1 U12797 ( .A(weight_queue_7__4__1_), .ZN(n19442) );
  INV_X1 U12798 ( .A(n19442), .ZN(n19443) );
  INV_X1 U12799 ( .A(n17162), .ZN(n19444) );
  INV_X1 U12800 ( .A(weight_queue_7__4__2_), .ZN(n19445) );
  INV_X1 U12801 ( .A(n19445), .ZN(n19446) );
  INV_X1 U12802 ( .A(n17163), .ZN(n19447) );
  INV_X1 U12803 ( .A(weight_queue_7__4__3_), .ZN(n19448) );
  INV_X1 U12804 ( .A(n19448), .ZN(n19449) );
  INV_X1 U12805 ( .A(n17164), .ZN(n19450) );
  INV_X1 U12806 ( .A(weight_queue_7__4__4_), .ZN(n19451) );
  INV_X1 U12807 ( .A(n19451), .ZN(n19452) );
  INV_X1 U12808 ( .A(n17165), .ZN(n19453) );
  INV_X1 U12809 ( .A(weight_queue_7__4__5_), .ZN(n19454) );
  INV_X1 U12810 ( .A(n19454), .ZN(n19455) );
  INV_X1 U12811 ( .A(n17166), .ZN(n19456) );
  INV_X1 U12812 ( .A(weight_queue_7__4__6_), .ZN(n19457) );
  INV_X1 U12813 ( .A(n19457), .ZN(n19458) );
  INV_X1 U12814 ( .A(n17167), .ZN(n19459) );
  INV_X1 U12815 ( .A(weight_queue_7__4__7_), .ZN(n19460) );
  INV_X1 U12816 ( .A(n17168), .ZN(n19461) );
  INV_X1 U12817 ( .A(n19460), .ZN(n19462) );
  INV_X1 U12818 ( .A(weight_queue_7__3__0_), .ZN(n19463) );
  INV_X1 U12819 ( .A(n19463), .ZN(n19464) );
  INV_X1 U12820 ( .A(n17169), .ZN(n19465) );
  INV_X1 U12821 ( .A(weight_queue_7__3__1_), .ZN(n19466) );
  INV_X1 U12822 ( .A(n19466), .ZN(n19467) );
  INV_X1 U12823 ( .A(n17170), .ZN(n19468) );
  INV_X1 U12824 ( .A(weight_queue_7__3__2_), .ZN(n19469) );
  INV_X1 U12825 ( .A(n19469), .ZN(n19470) );
  INV_X1 U12826 ( .A(n17171), .ZN(n19471) );
  INV_X1 U12827 ( .A(weight_queue_7__3__3_), .ZN(n19472) );
  INV_X1 U12828 ( .A(n19472), .ZN(n19473) );
  INV_X1 U12829 ( .A(n17172), .ZN(n19474) );
  INV_X1 U12830 ( .A(weight_queue_7__3__4_), .ZN(n19475) );
  INV_X1 U12831 ( .A(n19475), .ZN(n19476) );
  INV_X1 U12832 ( .A(n17173), .ZN(n19477) );
  INV_X1 U12833 ( .A(weight_queue_7__3__5_), .ZN(n19478) );
  INV_X1 U12834 ( .A(n19478), .ZN(n19479) );
  INV_X1 U12835 ( .A(n17174), .ZN(n19480) );
  INV_X1 U12836 ( .A(weight_queue_7__3__6_), .ZN(n19481) );
  INV_X1 U12837 ( .A(n19481), .ZN(n19482) );
  INV_X1 U12838 ( .A(n17175), .ZN(n19483) );
  INV_X1 U12839 ( .A(weight_queue_7__3__7_), .ZN(n19484) );
  INV_X1 U12840 ( .A(n17176), .ZN(n19485) );
  INV_X1 U12841 ( .A(n19484), .ZN(n19486) );
  INV_X1 U12842 ( .A(weight_queue_7__2__0_), .ZN(n19487) );
  INV_X1 U12843 ( .A(n19487), .ZN(n19488) );
  INV_X1 U12844 ( .A(n17177), .ZN(n19489) );
  INV_X1 U12845 ( .A(weight_queue_7__2__1_), .ZN(n19490) );
  INV_X1 U12846 ( .A(n19490), .ZN(n19491) );
  INV_X1 U12847 ( .A(n17178), .ZN(n19492) );
  INV_X1 U12848 ( .A(weight_queue_7__2__2_), .ZN(n19493) );
  INV_X1 U12849 ( .A(n19493), .ZN(n19494) );
  INV_X1 U12850 ( .A(n17179), .ZN(n19495) );
  INV_X1 U12851 ( .A(weight_queue_7__2__3_), .ZN(n19496) );
  INV_X1 U12852 ( .A(n19496), .ZN(n19497) );
  INV_X1 U12853 ( .A(n17180), .ZN(n19498) );
  INV_X1 U12854 ( .A(weight_queue_7__2__4_), .ZN(n19499) );
  INV_X1 U12855 ( .A(n19499), .ZN(n19500) );
  INV_X1 U12856 ( .A(n17181), .ZN(n19501) );
  INV_X1 U12857 ( .A(weight_queue_7__2__5_), .ZN(n19502) );
  INV_X1 U12858 ( .A(n19502), .ZN(n19503) );
  INV_X1 U12859 ( .A(n17182), .ZN(n19504) );
  INV_X1 U12860 ( .A(weight_queue_7__2__6_), .ZN(n19505) );
  INV_X1 U12861 ( .A(n19505), .ZN(n19506) );
  INV_X1 U12862 ( .A(n17183), .ZN(n19507) );
  INV_X1 U12863 ( .A(weight_queue_7__2__7_), .ZN(n19508) );
  INV_X1 U12864 ( .A(n17184), .ZN(n19509) );
  INV_X1 U12865 ( .A(n19508), .ZN(n19510) );
  INV_X1 U12866 ( .A(weight_queue_7__1__0_), .ZN(n19511) );
  INV_X1 U12867 ( .A(n19511), .ZN(n19512) );
  INV_X1 U12868 ( .A(n17185), .ZN(n19513) );
  INV_X1 U12869 ( .A(weight_queue_7__1__1_), .ZN(n19514) );
  INV_X1 U12870 ( .A(n19514), .ZN(n19515) );
  INV_X1 U12871 ( .A(n17186), .ZN(n19516) );
  INV_X1 U12872 ( .A(weight_queue_7__1__2_), .ZN(n19517) );
  INV_X1 U12873 ( .A(n19517), .ZN(n19518) );
  INV_X1 U12874 ( .A(n17187), .ZN(n19519) );
  INV_X1 U12875 ( .A(weight_queue_7__1__3_), .ZN(n19520) );
  INV_X1 U12876 ( .A(n19520), .ZN(n19521) );
  INV_X1 U12877 ( .A(n17188), .ZN(n19522) );
  INV_X1 U12878 ( .A(weight_queue_7__1__4_), .ZN(n19523) );
  INV_X1 U12879 ( .A(n19523), .ZN(n19524) );
  INV_X1 U12880 ( .A(n17189), .ZN(n19525) );
  INV_X1 U12881 ( .A(weight_queue_7__1__5_), .ZN(n19526) );
  INV_X1 U12882 ( .A(n19526), .ZN(n19527) );
  INV_X1 U12883 ( .A(n17190), .ZN(n19528) );
  INV_X1 U12884 ( .A(weight_queue_7__1__6_), .ZN(n19529) );
  INV_X1 U12885 ( .A(n19529), .ZN(n19530) );
  INV_X1 U12886 ( .A(n17191), .ZN(n19531) );
  INV_X1 U12887 ( .A(weight_queue_7__1__7_), .ZN(n19532) );
  INV_X1 U12888 ( .A(n17192), .ZN(n19533) );
  INV_X1 U12889 ( .A(n19532), .ZN(n19534) );
  INV_X1 U12890 ( .A(weight_queue_7__0__0_), .ZN(n19535) );
  INV_X1 U12891 ( .A(n19535), .ZN(n19536) );
  INV_X1 U12892 ( .A(n17193), .ZN(n19537) );
  INV_X1 U12893 ( .A(weight_queue_7__0__1_), .ZN(n19538) );
  INV_X1 U12894 ( .A(n19538), .ZN(n19539) );
  INV_X1 U12895 ( .A(n17194), .ZN(n19540) );
  INV_X1 U12896 ( .A(weight_queue_7__0__2_), .ZN(n19541) );
  INV_X1 U12897 ( .A(n19541), .ZN(n19542) );
  INV_X1 U12898 ( .A(n17195), .ZN(n19543) );
  INV_X1 U12899 ( .A(weight_queue_7__0__3_), .ZN(n19544) );
  INV_X1 U12900 ( .A(n19544), .ZN(n19545) );
  INV_X1 U12901 ( .A(n17196), .ZN(n19546) );
  INV_X1 U12902 ( .A(weight_queue_7__0__4_), .ZN(n19547) );
  INV_X1 U12903 ( .A(n19547), .ZN(n19548) );
  INV_X1 U12904 ( .A(n17197), .ZN(n19549) );
  INV_X1 U12905 ( .A(weight_queue_7__0__5_), .ZN(n19550) );
  INV_X1 U12906 ( .A(n19550), .ZN(n19551) );
  INV_X1 U12907 ( .A(n17198), .ZN(n19552) );
  INV_X1 U12908 ( .A(weight_queue_7__0__6_), .ZN(n19553) );
  INV_X1 U12909 ( .A(n19553), .ZN(n19554) );
  INV_X1 U12910 ( .A(n17199), .ZN(n19555) );
  INV_X1 U12911 ( .A(weight_queue_7__0__7_), .ZN(n19556) );
  INV_X1 U12912 ( .A(n17200), .ZN(n19557) );
  INV_X1 U12913 ( .A(n19556), .ZN(n19558) );
  INV_X1 U12914 ( .A(data_queue_7__7__0_), .ZN(n19559) );
  INV_X1 U12915 ( .A(n19559), .ZN(n19560) );
  INV_X1 U12916 ( .A(n17201), .ZN(n19561) );
  INV_X1 U12917 ( .A(data_queue_7__7__1_), .ZN(n19562) );
  INV_X1 U12918 ( .A(n19562), .ZN(n19563) );
  INV_X1 U12919 ( .A(n17202), .ZN(n19564) );
  INV_X1 U12920 ( .A(data_queue_7__7__2_), .ZN(n19565) );
  INV_X1 U12921 ( .A(n19565), .ZN(n19566) );
  INV_X1 U12922 ( .A(n17203), .ZN(n19567) );
  INV_X1 U12923 ( .A(data_queue_7__7__3_), .ZN(n19568) );
  INV_X1 U12924 ( .A(n19568), .ZN(n19569) );
  INV_X1 U12925 ( .A(n17204), .ZN(n19570) );
  INV_X1 U12926 ( .A(data_queue_7__7__4_), .ZN(n19571) );
  INV_X1 U12927 ( .A(n19571), .ZN(n19572) );
  INV_X1 U12928 ( .A(n17205), .ZN(n19573) );
  INV_X1 U12929 ( .A(data_queue_7__7__5_), .ZN(n19574) );
  INV_X1 U12930 ( .A(n19574), .ZN(n19575) );
  INV_X1 U12931 ( .A(n17206), .ZN(n19576) );
  INV_X1 U12932 ( .A(data_queue_7__7__6_), .ZN(n19577) );
  INV_X1 U12933 ( .A(n19577), .ZN(n19578) );
  INV_X1 U12934 ( .A(n17207), .ZN(n19579) );
  INV_X1 U12935 ( .A(data_queue_7__7__7_), .ZN(n19580) );
  INV_X1 U12936 ( .A(n19580), .ZN(n19581) );
  INV_X1 U12937 ( .A(n17208), .ZN(n19582) );
  INV_X1 U12938 ( .A(data_queue_6__7__0_), .ZN(n19583) );
  INV_X1 U12939 ( .A(n19583), .ZN(n19584) );
  INV_X1 U12940 ( .A(n17209), .ZN(n19585) );
  INV_X1 U12941 ( .A(data_queue_6__7__1_), .ZN(n19586) );
  INV_X1 U12942 ( .A(n19586), .ZN(n19587) );
  INV_X1 U12943 ( .A(n17210), .ZN(n19588) );
  INV_X1 U12944 ( .A(data_queue_6__7__2_), .ZN(n19589) );
  INV_X1 U12945 ( .A(n19589), .ZN(n19590) );
  INV_X1 U12946 ( .A(n17211), .ZN(n19591) );
  INV_X1 U12947 ( .A(data_queue_6__7__3_), .ZN(n19592) );
  INV_X1 U12948 ( .A(n19592), .ZN(n19593) );
  INV_X1 U12949 ( .A(n17212), .ZN(n19594) );
  INV_X1 U12950 ( .A(data_queue_6__7__4_), .ZN(n19595) );
  INV_X1 U12951 ( .A(n19595), .ZN(n19596) );
  INV_X1 U12952 ( .A(n17213), .ZN(n19597) );
  INV_X1 U12953 ( .A(data_queue_6__7__5_), .ZN(n19598) );
  INV_X1 U12954 ( .A(n19598), .ZN(n19599) );
  INV_X1 U12955 ( .A(n17214), .ZN(n19600) );
  INV_X1 U12956 ( .A(data_queue_6__7__6_), .ZN(n19601) );
  INV_X1 U12957 ( .A(n19601), .ZN(n19602) );
  INV_X1 U12958 ( .A(n17215), .ZN(n19603) );
  INV_X1 U12959 ( .A(data_queue_6__7__7_), .ZN(n19604) );
  INV_X1 U12960 ( .A(n19604), .ZN(n19605) );
  INV_X1 U12961 ( .A(n17216), .ZN(n19606) );
  INV_X1 U12962 ( .A(data_queue_5__7__0_), .ZN(n19607) );
  INV_X1 U12963 ( .A(n19607), .ZN(n19608) );
  INV_X1 U12964 ( .A(n17217), .ZN(n19609) );
  INV_X1 U12965 ( .A(data_queue_5__7__1_), .ZN(n19610) );
  INV_X1 U12966 ( .A(n19610), .ZN(n19611) );
  INV_X1 U12967 ( .A(n17218), .ZN(n19612) );
  INV_X1 U12968 ( .A(data_queue_5__7__2_), .ZN(n19613) );
  INV_X1 U12969 ( .A(n19613), .ZN(n19614) );
  INV_X1 U12970 ( .A(n17219), .ZN(n19615) );
  INV_X1 U12971 ( .A(data_queue_5__7__3_), .ZN(n19616) );
  INV_X1 U12972 ( .A(n19616), .ZN(n19617) );
  INV_X1 U12973 ( .A(n17220), .ZN(n19618) );
  INV_X1 U12974 ( .A(data_queue_5__7__4_), .ZN(n19619) );
  INV_X1 U12975 ( .A(n19619), .ZN(n19620) );
  INV_X1 U12976 ( .A(n17221), .ZN(n19621) );
  INV_X1 U12977 ( .A(data_queue_5__7__5_), .ZN(n19622) );
  INV_X1 U12978 ( .A(n19622), .ZN(n19623) );
  INV_X1 U12979 ( .A(n17222), .ZN(n19624) );
  INV_X1 U12980 ( .A(data_queue_5__7__6_), .ZN(n19625) );
  INV_X1 U12981 ( .A(n19625), .ZN(n19626) );
  INV_X1 U12982 ( .A(n17223), .ZN(n19627) );
  INV_X1 U12983 ( .A(data_queue_5__7__7_), .ZN(n19628) );
  INV_X1 U12984 ( .A(n19628), .ZN(n19629) );
  INV_X1 U12985 ( .A(n17224), .ZN(n19630) );
  INV_X1 U12986 ( .A(data_queue_4__7__0_), .ZN(n19631) );
  INV_X1 U12987 ( .A(n19631), .ZN(n19632) );
  INV_X1 U12988 ( .A(n17225), .ZN(n19633) );
  INV_X1 U12989 ( .A(data_queue_4__7__1_), .ZN(n19634) );
  INV_X1 U12990 ( .A(n19634), .ZN(n19635) );
  INV_X1 U12991 ( .A(n17226), .ZN(n19636) );
  INV_X1 U12992 ( .A(data_queue_4__7__2_), .ZN(n19637) );
  INV_X1 U12993 ( .A(n19637), .ZN(n19638) );
  INV_X1 U12994 ( .A(n17227), .ZN(n19639) );
  INV_X1 U12995 ( .A(data_queue_4__7__3_), .ZN(n19640) );
  INV_X1 U12996 ( .A(n19640), .ZN(n19641) );
  INV_X1 U12997 ( .A(n17228), .ZN(n19642) );
  INV_X1 U12998 ( .A(data_queue_4__7__4_), .ZN(n19643) );
  INV_X1 U12999 ( .A(n19643), .ZN(n19644) );
  INV_X1 U13000 ( .A(n17229), .ZN(n19645) );
  INV_X1 U13001 ( .A(data_queue_4__7__5_), .ZN(n19646) );
  INV_X1 U13002 ( .A(n19646), .ZN(n19647) );
  INV_X1 U13003 ( .A(n17230), .ZN(n19648) );
  INV_X1 U13004 ( .A(data_queue_4__7__6_), .ZN(n19649) );
  INV_X1 U13005 ( .A(n19649), .ZN(n19650) );
  INV_X1 U13006 ( .A(n17231), .ZN(n19651) );
  INV_X1 U13007 ( .A(data_queue_4__7__7_), .ZN(n19652) );
  INV_X1 U13008 ( .A(n19652), .ZN(n19653) );
  INV_X1 U13009 ( .A(n17232), .ZN(n19654) );
  INV_X1 U13010 ( .A(data_queue_3__7__0_), .ZN(n19655) );
  INV_X1 U13011 ( .A(n19655), .ZN(n19656) );
  INV_X1 U13012 ( .A(n17233), .ZN(n19657) );
  INV_X1 U13013 ( .A(data_queue_3__7__1_), .ZN(n19658) );
  INV_X1 U13014 ( .A(n19658), .ZN(n19659) );
  INV_X1 U13015 ( .A(n17234), .ZN(n19660) );
  INV_X1 U13016 ( .A(data_queue_3__7__2_), .ZN(n19661) );
  INV_X1 U13017 ( .A(n19661), .ZN(n19662) );
  INV_X1 U13018 ( .A(n17235), .ZN(n19663) );
  INV_X1 U13019 ( .A(data_queue_3__7__3_), .ZN(n19664) );
  INV_X1 U13020 ( .A(n19664), .ZN(n19665) );
  INV_X1 U13021 ( .A(n17236), .ZN(n19666) );
  INV_X1 U13022 ( .A(data_queue_3__7__4_), .ZN(n19667) );
  INV_X1 U13023 ( .A(n19667), .ZN(n19668) );
  INV_X1 U13024 ( .A(n17237), .ZN(n19669) );
  INV_X1 U13025 ( .A(data_queue_3__7__5_), .ZN(n19670) );
  INV_X1 U13026 ( .A(n19670), .ZN(n19671) );
  INV_X1 U13027 ( .A(n17238), .ZN(n19672) );
  INV_X1 U13028 ( .A(data_queue_3__7__6_), .ZN(n19673) );
  INV_X1 U13029 ( .A(n19673), .ZN(n19674) );
  INV_X1 U13030 ( .A(n17239), .ZN(n19675) );
  INV_X1 U13031 ( .A(data_queue_3__7__7_), .ZN(n19676) );
  INV_X1 U13032 ( .A(n19676), .ZN(n19677) );
  INV_X1 U13033 ( .A(n17240), .ZN(n19678) );
  INV_X1 U13034 ( .A(data_queue_2__7__0_), .ZN(n19679) );
  INV_X1 U13035 ( .A(n19679), .ZN(n19680) );
  INV_X1 U13036 ( .A(n17241), .ZN(n19681) );
  INV_X1 U13037 ( .A(data_queue_2__7__1_), .ZN(n19682) );
  INV_X1 U13038 ( .A(n19682), .ZN(n19683) );
  INV_X1 U13039 ( .A(n17242), .ZN(n19684) );
  INV_X1 U13040 ( .A(data_queue_2__7__2_), .ZN(n19685) );
  INV_X1 U13041 ( .A(n19685), .ZN(n19686) );
  INV_X1 U13042 ( .A(n17243), .ZN(n19687) );
  INV_X1 U13043 ( .A(data_queue_2__7__3_), .ZN(n19688) );
  INV_X1 U13044 ( .A(n19688), .ZN(n19689) );
  INV_X1 U13045 ( .A(n17244), .ZN(n19690) );
  INV_X1 U13046 ( .A(data_queue_2__7__4_), .ZN(n19691) );
  INV_X1 U13047 ( .A(n19691), .ZN(n19692) );
  INV_X1 U13048 ( .A(n17245), .ZN(n19693) );
  INV_X1 U13049 ( .A(data_queue_2__7__5_), .ZN(n19694) );
  INV_X1 U13050 ( .A(n19694), .ZN(n19695) );
  INV_X1 U13051 ( .A(n17246), .ZN(n19696) );
  INV_X1 U13052 ( .A(data_queue_2__7__6_), .ZN(n19697) );
  INV_X1 U13053 ( .A(n19697), .ZN(n19698) );
  INV_X1 U13054 ( .A(n17247), .ZN(n19699) );
  INV_X1 U13055 ( .A(data_queue_2__7__7_), .ZN(n19700) );
  INV_X1 U13056 ( .A(n19700), .ZN(n19701) );
  INV_X1 U13057 ( .A(n17248), .ZN(n19702) );
  INV_X1 U13058 ( .A(data_queue_1__7__0_), .ZN(n19703) );
  INV_X1 U13059 ( .A(n19703), .ZN(n19704) );
  INV_X1 U13060 ( .A(n17249), .ZN(n19705) );
  INV_X1 U13061 ( .A(data_queue_1__7__1_), .ZN(n19706) );
  INV_X1 U13062 ( .A(n19706), .ZN(n19707) );
  INV_X1 U13063 ( .A(n17250), .ZN(n19708) );
  INV_X1 U13064 ( .A(data_queue_1__7__2_), .ZN(n19709) );
  INV_X1 U13065 ( .A(n19709), .ZN(n19710) );
  INV_X1 U13066 ( .A(n17251), .ZN(n19711) );
  INV_X1 U13067 ( .A(data_queue_1__7__3_), .ZN(n19712) );
  INV_X1 U13068 ( .A(n19712), .ZN(n19713) );
  INV_X1 U13069 ( .A(n17252), .ZN(n19714) );
  INV_X1 U13070 ( .A(data_queue_1__7__4_), .ZN(n19715) );
  INV_X1 U13071 ( .A(n19715), .ZN(n19716) );
  INV_X1 U13072 ( .A(n17253), .ZN(n19717) );
  INV_X1 U13073 ( .A(data_queue_1__7__5_), .ZN(n19718) );
  INV_X1 U13074 ( .A(n19718), .ZN(n19719) );
  INV_X1 U13075 ( .A(n17254), .ZN(n19720) );
  INV_X1 U13076 ( .A(data_queue_1__7__6_), .ZN(n19721) );
  INV_X1 U13077 ( .A(n19721), .ZN(n19722) );
  INV_X1 U13078 ( .A(n17255), .ZN(n19723) );
  INV_X1 U13079 ( .A(data_queue_1__7__7_), .ZN(n19724) );
  INV_X1 U13080 ( .A(n19724), .ZN(n19725) );
  INV_X1 U13081 ( .A(n17256), .ZN(n19726) );
  INV_X1 U13082 ( .A(data_queue_0__7__0_), .ZN(n19727) );
  INV_X1 U13083 ( .A(n19727), .ZN(n19728) );
  INV_X1 U13084 ( .A(n17257), .ZN(n19729) );
  INV_X1 U13085 ( .A(data_queue_0__7__1_), .ZN(n19730) );
  INV_X1 U13086 ( .A(n19730), .ZN(n19731) );
  INV_X1 U13087 ( .A(n17258), .ZN(n19732) );
  INV_X1 U13088 ( .A(data_queue_0__7__2_), .ZN(n19733) );
  INV_X1 U13089 ( .A(n19733), .ZN(n19734) );
  INV_X1 U13090 ( .A(n17259), .ZN(n19735) );
  INV_X1 U13091 ( .A(data_queue_0__7__3_), .ZN(n19736) );
  INV_X1 U13092 ( .A(n19736), .ZN(n19737) );
  INV_X1 U13093 ( .A(n17260), .ZN(n19738) );
  INV_X1 U13094 ( .A(data_queue_0__7__4_), .ZN(n19739) );
  INV_X1 U13095 ( .A(n19739), .ZN(n19740) );
  INV_X1 U13096 ( .A(n17261), .ZN(n19741) );
  INV_X1 U13097 ( .A(data_queue_0__7__5_), .ZN(n19742) );
  INV_X1 U13098 ( .A(n19742), .ZN(n19743) );
  INV_X1 U13099 ( .A(n17262), .ZN(n19744) );
  INV_X1 U13100 ( .A(data_queue_0__7__6_), .ZN(n19745) );
  INV_X1 U13101 ( .A(n19745), .ZN(n19746) );
  INV_X1 U13102 ( .A(n17263), .ZN(n19747) );
  INV_X1 U13103 ( .A(data_queue_0__7__7_), .ZN(n19748) );
  INV_X1 U13104 ( .A(n19748), .ZN(n19749) );
  INV_X1 U13105 ( .A(n17264), .ZN(n19750) );
  INV_X1 U13106 ( .A(n17267), .ZN(n19751) );
  INV_X1 U13107 ( .A(n17267), .ZN(n19752) );
  INV_X1 U13108 ( .A(n54230), .ZN(n19753) );
  INV_X1 U13109 ( .A(n19753), .ZN(n19754) );
  INV_X1 U13110 ( .A(n19753), .ZN(n19755) );
  INV_X1 U13111 ( .A(n17269), .ZN(n19756) );
  INV_X1 U13112 ( .A(n17269), .ZN(n19757) );
  INV_X1 U13113 ( .A(matrix_mul_2D_7__7__20_), .ZN(n19758) );
  INV_X1 U13114 ( .A(n19758), .ZN(n19759) );
  INV_X1 U13115 ( .A(matrix_mul_2D_7__7__19_), .ZN(n19760) );
  INV_X1 U13116 ( .A(n19760), .ZN(n19761) );
  INV_X1 U13117 ( .A(matrix_mul_2D_7__7__18_), .ZN(n19762) );
  INV_X1 U13118 ( .A(n19762), .ZN(n19763) );
  INV_X1 U13119 ( .A(matrix_mul_2D_7__7__17_), .ZN(n19764) );
  INV_X1 U13120 ( .A(n19764), .ZN(n19765) );
  INV_X1 U13121 ( .A(matrix_mul_2D_7__7__16_), .ZN(n19766) );
  INV_X1 U13122 ( .A(n19766), .ZN(n19767) );
  INV_X1 U13123 ( .A(matrix_mul_2D_7__7__15_), .ZN(n19768) );
  INV_X1 U13124 ( .A(n19768), .ZN(n19769) );
  INV_X1 U13125 ( .A(matrix_mul_2D_7__6__20_), .ZN(n19770) );
  INV_X1 U13126 ( .A(n19770), .ZN(n19771) );
  INV_X1 U13127 ( .A(matrix_mul_2D_7__6__19_), .ZN(n19772) );
  INV_X1 U13128 ( .A(n19772), .ZN(n19773) );
  INV_X1 U13129 ( .A(matrix_mul_2D_7__6__18_), .ZN(n19774) );
  INV_X1 U13130 ( .A(n19774), .ZN(n19775) );
  INV_X1 U13131 ( .A(matrix_mul_2D_7__6__17_), .ZN(n19776) );
  INV_X1 U13132 ( .A(n19776), .ZN(n19777) );
  INV_X1 U13133 ( .A(matrix_mul_2D_7__6__16_), .ZN(n19778) );
  INV_X1 U13134 ( .A(n19778), .ZN(n19779) );
  INV_X1 U13135 ( .A(matrix_mul_2D_7__6__15_), .ZN(n19780) );
  INV_X1 U13136 ( .A(n19780), .ZN(n19781) );
  INV_X1 U13137 ( .A(matrix_mul_2D_7__5__20_), .ZN(n19782) );
  INV_X1 U13138 ( .A(n19782), .ZN(n19783) );
  INV_X1 U13139 ( .A(matrix_mul_2D_7__5__19_), .ZN(n19784) );
  INV_X1 U13140 ( .A(n19784), .ZN(n19785) );
  INV_X1 U13141 ( .A(matrix_mul_2D_7__5__18_), .ZN(n19786) );
  INV_X1 U13142 ( .A(n19786), .ZN(n19787) );
  INV_X1 U13143 ( .A(matrix_mul_2D_7__5__17_), .ZN(n19788) );
  INV_X1 U13144 ( .A(n19788), .ZN(n19789) );
  INV_X1 U13145 ( .A(matrix_mul_2D_7__5__16_), .ZN(n19790) );
  INV_X1 U13146 ( .A(n19790), .ZN(n19791) );
  INV_X1 U13147 ( .A(matrix_mul_2D_7__5__15_), .ZN(n19792) );
  INV_X1 U13148 ( .A(n19792), .ZN(n19793) );
  INV_X1 U13149 ( .A(matrix_mul_2D_7__4__20_), .ZN(n19794) );
  INV_X1 U13150 ( .A(n19794), .ZN(n19795) );
  INV_X1 U13151 ( .A(matrix_mul_2D_7__4__19_), .ZN(n19796) );
  INV_X1 U13152 ( .A(n19796), .ZN(n19797) );
  INV_X1 U13153 ( .A(matrix_mul_2D_7__4__18_), .ZN(n19798) );
  INV_X1 U13154 ( .A(n19798), .ZN(n19799) );
  INV_X1 U13155 ( .A(matrix_mul_2D_7__4__17_), .ZN(n19800) );
  INV_X1 U13156 ( .A(n19800), .ZN(n19801) );
  INV_X1 U13157 ( .A(matrix_mul_2D_7__4__16_), .ZN(n19802) );
  INV_X1 U13158 ( .A(n19802), .ZN(n19803) );
  INV_X1 U13159 ( .A(matrix_mul_2D_7__4__15_), .ZN(n19804) );
  INV_X1 U13160 ( .A(n19804), .ZN(n19805) );
  INV_X1 U13161 ( .A(matrix_mul_2D_7__3__20_), .ZN(n19806) );
  INV_X1 U13162 ( .A(n19806), .ZN(n19807) );
  INV_X1 U13163 ( .A(matrix_mul_2D_7__3__19_), .ZN(n19808) );
  INV_X1 U13164 ( .A(n19808), .ZN(n19809) );
  INV_X1 U13165 ( .A(matrix_mul_2D_7__3__18_), .ZN(n19810) );
  INV_X1 U13166 ( .A(n19810), .ZN(n19811) );
  INV_X1 U13167 ( .A(matrix_mul_2D_7__3__17_), .ZN(n19812) );
  INV_X1 U13168 ( .A(n19812), .ZN(n19813) );
  INV_X1 U13169 ( .A(matrix_mul_2D_7__3__16_), .ZN(n19814) );
  INV_X1 U13170 ( .A(n19814), .ZN(n19815) );
  INV_X1 U13171 ( .A(matrix_mul_2D_7__3__15_), .ZN(n19816) );
  INV_X1 U13172 ( .A(n19816), .ZN(n19817) );
  INV_X1 U13173 ( .A(matrix_mul_2D_7__2__20_), .ZN(n19818) );
  INV_X1 U13174 ( .A(n19818), .ZN(n19819) );
  INV_X1 U13175 ( .A(matrix_mul_2D_7__2__19_), .ZN(n19820) );
  INV_X1 U13176 ( .A(n19820), .ZN(n19821) );
  INV_X1 U13177 ( .A(matrix_mul_2D_7__2__18_), .ZN(n19822) );
  INV_X1 U13178 ( .A(n19822), .ZN(n19823) );
  INV_X1 U13179 ( .A(matrix_mul_2D_7__2__17_), .ZN(n19824) );
  INV_X1 U13180 ( .A(n19824), .ZN(n19825) );
  INV_X1 U13181 ( .A(matrix_mul_2D_7__2__16_), .ZN(n19826) );
  INV_X1 U13182 ( .A(n19826), .ZN(n19827) );
  INV_X1 U13183 ( .A(matrix_mul_2D_7__2__15_), .ZN(n19828) );
  INV_X1 U13184 ( .A(n19828), .ZN(n19829) );
  INV_X1 U13185 ( .A(matrix_mul_2D_7__1__20_), .ZN(n19830) );
  INV_X1 U13186 ( .A(n19830), .ZN(n19831) );
  INV_X1 U13187 ( .A(matrix_mul_2D_7__1__19_), .ZN(n19832) );
  INV_X1 U13188 ( .A(n19832), .ZN(n19833) );
  INV_X1 U13189 ( .A(matrix_mul_2D_7__1__18_), .ZN(n19834) );
  INV_X1 U13190 ( .A(n19834), .ZN(n19835) );
  INV_X1 U13191 ( .A(matrix_mul_2D_7__1__17_), .ZN(n19836) );
  INV_X1 U13192 ( .A(n19836), .ZN(n19837) );
  INV_X1 U13193 ( .A(matrix_mul_2D_7__1__16_), .ZN(n19838) );
  INV_X1 U13194 ( .A(n19838), .ZN(n19839) );
  INV_X1 U13195 ( .A(matrix_mul_2D_7__1__15_), .ZN(n19840) );
  INV_X1 U13196 ( .A(n19840), .ZN(n19841) );
  INV_X1 U13197 ( .A(matrix_mul_2D_7__0__20_), .ZN(n19842) );
  INV_X1 U13198 ( .A(n19842), .ZN(n19843) );
  INV_X1 U13199 ( .A(matrix_mul_2D_7__0__19_), .ZN(n19844) );
  INV_X1 U13200 ( .A(n19844), .ZN(n19845) );
  INV_X1 U13201 ( .A(matrix_mul_2D_7__0__18_), .ZN(n19846) );
  INV_X1 U13202 ( .A(n19846), .ZN(n19847) );
  INV_X1 U13203 ( .A(matrix_mul_2D_7__0__17_), .ZN(n19848) );
  INV_X1 U13204 ( .A(n19848), .ZN(n19849) );
  INV_X1 U13205 ( .A(matrix_mul_2D_7__0__16_), .ZN(n19850) );
  INV_X1 U13206 ( .A(n19850), .ZN(n19851) );
  INV_X1 U13207 ( .A(matrix_mul_2D_7__0__15_), .ZN(n19852) );
  INV_X1 U13208 ( .A(n19852), .ZN(n19853) );
  INV_X1 U13209 ( .A(matrix_mul_2D_6__7__20_), .ZN(n19854) );
  INV_X1 U13210 ( .A(n19854), .ZN(n19855) );
  INV_X1 U13211 ( .A(matrix_mul_2D_6__7__19_), .ZN(n19856) );
  INV_X1 U13212 ( .A(n19856), .ZN(n19857) );
  INV_X1 U13213 ( .A(matrix_mul_2D_6__7__18_), .ZN(n19858) );
  INV_X1 U13214 ( .A(n19858), .ZN(n19859) );
  INV_X1 U13215 ( .A(matrix_mul_2D_6__7__17_), .ZN(n19860) );
  INV_X1 U13216 ( .A(n19860), .ZN(n19861) );
  INV_X1 U13217 ( .A(matrix_mul_2D_6__7__16_), .ZN(n19862) );
  INV_X1 U13218 ( .A(n19862), .ZN(n19863) );
  INV_X1 U13219 ( .A(matrix_mul_2D_6__7__15_), .ZN(n19864) );
  INV_X1 U13220 ( .A(n19864), .ZN(n19865) );
  INV_X1 U13221 ( .A(matrix_mul_2D_6__6__20_), .ZN(n19866) );
  INV_X1 U13222 ( .A(n19866), .ZN(n19867) );
  INV_X1 U13223 ( .A(matrix_mul_2D_6__6__19_), .ZN(n19868) );
  INV_X1 U13224 ( .A(n19868), .ZN(n19869) );
  INV_X1 U13225 ( .A(matrix_mul_2D_6__6__18_), .ZN(n19870) );
  INV_X1 U13226 ( .A(n19870), .ZN(n19871) );
  INV_X1 U13227 ( .A(matrix_mul_2D_6__6__17_), .ZN(n19872) );
  INV_X1 U13228 ( .A(n19872), .ZN(n19873) );
  INV_X1 U13229 ( .A(matrix_mul_2D_6__6__16_), .ZN(n19874) );
  INV_X1 U13230 ( .A(n19874), .ZN(n19875) );
  INV_X1 U13231 ( .A(matrix_mul_2D_6__6__15_), .ZN(n19876) );
  INV_X1 U13232 ( .A(n19876), .ZN(n19877) );
  INV_X1 U13233 ( .A(matrix_mul_2D_6__5__20_), .ZN(n19878) );
  INV_X1 U13234 ( .A(n19878), .ZN(n19879) );
  INV_X1 U13235 ( .A(matrix_mul_2D_6__5__19_), .ZN(n19880) );
  INV_X1 U13236 ( .A(n19880), .ZN(n19881) );
  INV_X1 U13237 ( .A(matrix_mul_2D_6__5__18_), .ZN(n19882) );
  INV_X1 U13238 ( .A(n19882), .ZN(n19883) );
  INV_X1 U13239 ( .A(matrix_mul_2D_6__5__17_), .ZN(n19884) );
  INV_X1 U13240 ( .A(n19884), .ZN(n19885) );
  INV_X1 U13241 ( .A(matrix_mul_2D_6__5__16_), .ZN(n19886) );
  INV_X1 U13242 ( .A(n19886), .ZN(n19887) );
  INV_X1 U13243 ( .A(matrix_mul_2D_6__5__15_), .ZN(n19888) );
  INV_X1 U13244 ( .A(n19888), .ZN(n19889) );
  INV_X1 U13245 ( .A(matrix_mul_2D_6__4__20_), .ZN(n19890) );
  INV_X1 U13246 ( .A(n19890), .ZN(n19891) );
  INV_X1 U13247 ( .A(matrix_mul_2D_6__4__19_), .ZN(n19892) );
  INV_X1 U13248 ( .A(n19892), .ZN(n19893) );
  INV_X1 U13249 ( .A(matrix_mul_2D_6__4__18_), .ZN(n19894) );
  INV_X1 U13250 ( .A(n19894), .ZN(n19895) );
  INV_X1 U13251 ( .A(matrix_mul_2D_6__4__17_), .ZN(n19896) );
  INV_X1 U13252 ( .A(n19896), .ZN(n19897) );
  INV_X1 U13253 ( .A(matrix_mul_2D_6__4__16_), .ZN(n19898) );
  INV_X1 U13254 ( .A(n19898), .ZN(n19899) );
  INV_X1 U13255 ( .A(matrix_mul_2D_6__4__15_), .ZN(n19900) );
  INV_X1 U13256 ( .A(n19900), .ZN(n19901) );
  INV_X1 U13257 ( .A(matrix_mul_2D_6__3__20_), .ZN(n19902) );
  INV_X1 U13258 ( .A(n19902), .ZN(n19903) );
  INV_X1 U13259 ( .A(matrix_mul_2D_6__3__19_), .ZN(n19904) );
  INV_X1 U13260 ( .A(n19904), .ZN(n19905) );
  INV_X1 U13261 ( .A(matrix_mul_2D_6__3__18_), .ZN(n19906) );
  INV_X1 U13262 ( .A(n19906), .ZN(n19907) );
  INV_X1 U13263 ( .A(matrix_mul_2D_6__3__17_), .ZN(n19908) );
  INV_X1 U13264 ( .A(n19908), .ZN(n19909) );
  INV_X1 U13265 ( .A(matrix_mul_2D_6__3__16_), .ZN(n19910) );
  INV_X1 U13266 ( .A(n19910), .ZN(n19911) );
  INV_X1 U13267 ( .A(matrix_mul_2D_6__3__15_), .ZN(n19912) );
  INV_X1 U13268 ( .A(n19912), .ZN(n19913) );
  INV_X1 U13269 ( .A(matrix_mul_2D_6__2__20_), .ZN(n19914) );
  INV_X1 U13270 ( .A(n19914), .ZN(n19915) );
  INV_X1 U13271 ( .A(matrix_mul_2D_6__2__19_), .ZN(n19916) );
  INV_X1 U13272 ( .A(n19916), .ZN(n19917) );
  INV_X1 U13273 ( .A(matrix_mul_2D_6__2__18_), .ZN(n19918) );
  INV_X1 U13274 ( .A(n19918), .ZN(n19919) );
  INV_X1 U13275 ( .A(matrix_mul_2D_6__2__17_), .ZN(n19920) );
  INV_X1 U13276 ( .A(n19920), .ZN(n19921) );
  INV_X1 U13277 ( .A(matrix_mul_2D_6__2__16_), .ZN(n19922) );
  INV_X1 U13278 ( .A(n19922), .ZN(n19923) );
  INV_X1 U13279 ( .A(matrix_mul_2D_6__2__15_), .ZN(n19924) );
  INV_X1 U13280 ( .A(n19924), .ZN(n19925) );
  INV_X1 U13281 ( .A(matrix_mul_2D_6__1__20_), .ZN(n19926) );
  INV_X1 U13282 ( .A(n19926), .ZN(n19927) );
  INV_X1 U13283 ( .A(matrix_mul_2D_6__1__19_), .ZN(n19928) );
  INV_X1 U13284 ( .A(n19928), .ZN(n19929) );
  INV_X1 U13285 ( .A(matrix_mul_2D_6__1__18_), .ZN(n19930) );
  INV_X1 U13286 ( .A(n19930), .ZN(n19931) );
  INV_X1 U13287 ( .A(matrix_mul_2D_6__1__17_), .ZN(n19932) );
  INV_X1 U13288 ( .A(n19932), .ZN(n19933) );
  INV_X1 U13289 ( .A(matrix_mul_2D_6__1__16_), .ZN(n19934) );
  INV_X1 U13290 ( .A(n19934), .ZN(n19935) );
  INV_X1 U13291 ( .A(matrix_mul_2D_6__1__15_), .ZN(n19936) );
  INV_X1 U13292 ( .A(n19936), .ZN(n19937) );
  INV_X1 U13293 ( .A(matrix_mul_2D_6__0__20_), .ZN(n19938) );
  INV_X1 U13294 ( .A(n19938), .ZN(n19939) );
  INV_X1 U13295 ( .A(matrix_mul_2D_6__0__19_), .ZN(n19940) );
  INV_X1 U13296 ( .A(n19940), .ZN(n19941) );
  INV_X1 U13297 ( .A(matrix_mul_2D_6__0__18_), .ZN(n19942) );
  INV_X1 U13298 ( .A(n19942), .ZN(n19943) );
  INV_X1 U13299 ( .A(matrix_mul_2D_6__0__17_), .ZN(n19944) );
  INV_X1 U13300 ( .A(n19944), .ZN(n19945) );
  INV_X1 U13301 ( .A(matrix_mul_2D_6__0__16_), .ZN(n19946) );
  INV_X1 U13302 ( .A(n19946), .ZN(n19947) );
  INV_X1 U13303 ( .A(matrix_mul_2D_6__0__15_), .ZN(n19948) );
  INV_X1 U13304 ( .A(n19948), .ZN(n19949) );
  INV_X1 U13305 ( .A(matrix_mul_2D_5__7__20_), .ZN(n19950) );
  INV_X1 U13306 ( .A(n19950), .ZN(n19951) );
  INV_X1 U13307 ( .A(matrix_mul_2D_5__7__19_), .ZN(n19952) );
  INV_X1 U13308 ( .A(n19952), .ZN(n19953) );
  INV_X1 U13309 ( .A(matrix_mul_2D_5__7__18_), .ZN(n19954) );
  INV_X1 U13310 ( .A(n19954), .ZN(n19955) );
  INV_X1 U13311 ( .A(matrix_mul_2D_5__7__17_), .ZN(n19956) );
  INV_X1 U13312 ( .A(n19956), .ZN(n19957) );
  INV_X1 U13313 ( .A(matrix_mul_2D_5__7__16_), .ZN(n19958) );
  INV_X1 U13314 ( .A(n19958), .ZN(n19959) );
  INV_X1 U13315 ( .A(matrix_mul_2D_5__7__15_), .ZN(n19960) );
  INV_X1 U13316 ( .A(n19960), .ZN(n19961) );
  INV_X1 U13317 ( .A(matrix_mul_2D_5__6__20_), .ZN(n19962) );
  INV_X1 U13318 ( .A(n19962), .ZN(n19963) );
  INV_X1 U13319 ( .A(matrix_mul_2D_5__6__19_), .ZN(n19964) );
  INV_X1 U13320 ( .A(n19964), .ZN(n19965) );
  INV_X1 U13321 ( .A(matrix_mul_2D_5__6__18_), .ZN(n19966) );
  INV_X1 U13322 ( .A(n19966), .ZN(n19967) );
  INV_X1 U13323 ( .A(matrix_mul_2D_5__6__17_), .ZN(n19968) );
  INV_X1 U13324 ( .A(n19968), .ZN(n19969) );
  INV_X1 U13325 ( .A(matrix_mul_2D_5__6__16_), .ZN(n19970) );
  INV_X1 U13326 ( .A(n19970), .ZN(n19971) );
  INV_X1 U13327 ( .A(matrix_mul_2D_5__6__15_), .ZN(n19972) );
  INV_X1 U13328 ( .A(n19972), .ZN(n19973) );
  INV_X1 U13329 ( .A(matrix_mul_2D_5__5__20_), .ZN(n19974) );
  INV_X1 U13330 ( .A(n19974), .ZN(n19975) );
  INV_X1 U13331 ( .A(matrix_mul_2D_5__5__19_), .ZN(n19976) );
  INV_X1 U13332 ( .A(n19976), .ZN(n19977) );
  INV_X1 U13333 ( .A(matrix_mul_2D_5__5__18_), .ZN(n19978) );
  INV_X1 U13334 ( .A(n19978), .ZN(n19979) );
  INV_X1 U13335 ( .A(matrix_mul_2D_5__5__17_), .ZN(n19980) );
  INV_X1 U13336 ( .A(n19980), .ZN(n19981) );
  INV_X1 U13337 ( .A(matrix_mul_2D_5__5__16_), .ZN(n19982) );
  INV_X1 U13338 ( .A(n19982), .ZN(n19983) );
  INV_X1 U13339 ( .A(matrix_mul_2D_5__5__15_), .ZN(n19984) );
  INV_X1 U13340 ( .A(n19984), .ZN(n19985) );
  INV_X1 U13341 ( .A(matrix_mul_2D_5__4__20_), .ZN(n19986) );
  INV_X1 U13342 ( .A(n19986), .ZN(n19987) );
  INV_X1 U13343 ( .A(matrix_mul_2D_5__4__19_), .ZN(n19988) );
  INV_X1 U13344 ( .A(n19988), .ZN(n19989) );
  INV_X1 U13345 ( .A(matrix_mul_2D_5__4__18_), .ZN(n19990) );
  INV_X1 U13346 ( .A(n19990), .ZN(n19991) );
  INV_X1 U13347 ( .A(matrix_mul_2D_5__4__17_), .ZN(n19992) );
  INV_X1 U13348 ( .A(n19992), .ZN(n19993) );
  INV_X1 U13349 ( .A(matrix_mul_2D_5__4__16_), .ZN(n19994) );
  INV_X1 U13350 ( .A(n19994), .ZN(n19995) );
  INV_X1 U13351 ( .A(matrix_mul_2D_5__4__15_), .ZN(n19996) );
  INV_X1 U13352 ( .A(n19996), .ZN(n19997) );
  INV_X1 U13353 ( .A(matrix_mul_2D_5__3__20_), .ZN(n19998) );
  INV_X1 U13354 ( .A(n19998), .ZN(n19999) );
  INV_X1 U13355 ( .A(matrix_mul_2D_5__3__19_), .ZN(n20000) );
  INV_X1 U13356 ( .A(n20000), .ZN(n20001) );
  INV_X1 U13357 ( .A(matrix_mul_2D_5__3__18_), .ZN(n20002) );
  INV_X1 U13358 ( .A(n20002), .ZN(n20003) );
  INV_X1 U13359 ( .A(matrix_mul_2D_5__3__17_), .ZN(n20004) );
  INV_X1 U13360 ( .A(n20004), .ZN(n20005) );
  INV_X1 U13361 ( .A(matrix_mul_2D_5__3__16_), .ZN(n20006) );
  INV_X1 U13362 ( .A(n20006), .ZN(n20007) );
  INV_X1 U13363 ( .A(matrix_mul_2D_5__3__15_), .ZN(n20008) );
  INV_X1 U13364 ( .A(n20008), .ZN(n20009) );
  INV_X1 U13365 ( .A(matrix_mul_2D_5__2__20_), .ZN(n20010) );
  INV_X1 U13366 ( .A(n20010), .ZN(n20011) );
  INV_X1 U13367 ( .A(matrix_mul_2D_5__2__19_), .ZN(n20012) );
  INV_X1 U13368 ( .A(n20012), .ZN(n20013) );
  INV_X1 U13369 ( .A(matrix_mul_2D_5__2__18_), .ZN(n20014) );
  INV_X1 U13370 ( .A(n20014), .ZN(n20015) );
  INV_X1 U13371 ( .A(matrix_mul_2D_5__2__17_), .ZN(n20016) );
  INV_X1 U13372 ( .A(n20016), .ZN(n20017) );
  INV_X1 U13373 ( .A(matrix_mul_2D_5__2__16_), .ZN(n20018) );
  INV_X1 U13374 ( .A(n20018), .ZN(n20019) );
  INV_X1 U13375 ( .A(matrix_mul_2D_5__2__15_), .ZN(n20020) );
  INV_X1 U13376 ( .A(n20020), .ZN(n20021) );
  INV_X1 U13377 ( .A(matrix_mul_2D_5__1__20_), .ZN(n20022) );
  INV_X1 U13378 ( .A(n20022), .ZN(n20023) );
  INV_X1 U13379 ( .A(matrix_mul_2D_5__1__19_), .ZN(n20024) );
  INV_X1 U13380 ( .A(n20024), .ZN(n20025) );
  INV_X1 U13381 ( .A(matrix_mul_2D_5__1__18_), .ZN(n20026) );
  INV_X1 U13382 ( .A(n20026), .ZN(n20027) );
  INV_X1 U13383 ( .A(matrix_mul_2D_5__1__17_), .ZN(n20028) );
  INV_X1 U13384 ( .A(n20028), .ZN(n20029) );
  INV_X1 U13385 ( .A(matrix_mul_2D_5__1__16_), .ZN(n20030) );
  INV_X1 U13386 ( .A(n20030), .ZN(n20031) );
  INV_X1 U13387 ( .A(matrix_mul_2D_5__1__15_), .ZN(n20032) );
  INV_X1 U13388 ( .A(n20032), .ZN(n20033) );
  INV_X1 U13389 ( .A(matrix_mul_2D_5__0__20_), .ZN(n20034) );
  INV_X1 U13390 ( .A(n20034), .ZN(n20035) );
  INV_X1 U13391 ( .A(matrix_mul_2D_5__0__19_), .ZN(n20036) );
  INV_X1 U13392 ( .A(n20036), .ZN(n20037) );
  INV_X1 U13393 ( .A(matrix_mul_2D_5__0__18_), .ZN(n20038) );
  INV_X1 U13394 ( .A(n20038), .ZN(n20039) );
  INV_X1 U13395 ( .A(matrix_mul_2D_5__0__17_), .ZN(n20040) );
  INV_X1 U13396 ( .A(n20040), .ZN(n20041) );
  INV_X1 U13397 ( .A(matrix_mul_2D_5__0__16_), .ZN(n20042) );
  INV_X1 U13398 ( .A(n20042), .ZN(n20043) );
  INV_X1 U13399 ( .A(matrix_mul_2D_5__0__15_), .ZN(n20044) );
  INV_X1 U13400 ( .A(n20044), .ZN(n20045) );
  INV_X1 U13401 ( .A(matrix_mul_2D_4__7__20_), .ZN(n20046) );
  INV_X1 U13402 ( .A(n20046), .ZN(n20047) );
  INV_X1 U13403 ( .A(matrix_mul_2D_4__7__19_), .ZN(n20048) );
  INV_X1 U13404 ( .A(n20048), .ZN(n20049) );
  INV_X1 U13405 ( .A(matrix_mul_2D_4__7__18_), .ZN(n20050) );
  INV_X1 U13406 ( .A(n20050), .ZN(n20051) );
  INV_X1 U13407 ( .A(matrix_mul_2D_4__7__17_), .ZN(n20052) );
  INV_X1 U13408 ( .A(n20052), .ZN(n20053) );
  INV_X1 U13409 ( .A(matrix_mul_2D_4__7__16_), .ZN(n20054) );
  INV_X1 U13410 ( .A(n20054), .ZN(n20055) );
  INV_X1 U13411 ( .A(matrix_mul_2D_4__7__15_), .ZN(n20056) );
  INV_X1 U13412 ( .A(n20056), .ZN(n20057) );
  INV_X1 U13413 ( .A(matrix_mul_2D_4__6__20_), .ZN(n20058) );
  INV_X1 U13414 ( .A(n20058), .ZN(n20059) );
  INV_X1 U13415 ( .A(matrix_mul_2D_4__6__19_), .ZN(n20060) );
  INV_X1 U13416 ( .A(n20060), .ZN(n20061) );
  INV_X1 U13417 ( .A(matrix_mul_2D_4__6__18_), .ZN(n20062) );
  INV_X1 U13418 ( .A(n20062), .ZN(n20063) );
  INV_X1 U13419 ( .A(matrix_mul_2D_4__6__17_), .ZN(n20064) );
  INV_X1 U13420 ( .A(n20064), .ZN(n20065) );
  INV_X1 U13421 ( .A(matrix_mul_2D_4__6__16_), .ZN(n20066) );
  INV_X1 U13422 ( .A(n20066), .ZN(n20067) );
  INV_X1 U13423 ( .A(matrix_mul_2D_4__6__15_), .ZN(n20068) );
  INV_X1 U13424 ( .A(n20068), .ZN(n20069) );
  INV_X1 U13425 ( .A(matrix_mul_2D_4__5__20_), .ZN(n20070) );
  INV_X1 U13426 ( .A(n20070), .ZN(n20071) );
  INV_X1 U13427 ( .A(matrix_mul_2D_4__5__19_), .ZN(n20072) );
  INV_X1 U13428 ( .A(n20072), .ZN(n20073) );
  INV_X1 U13429 ( .A(matrix_mul_2D_4__5__18_), .ZN(n20074) );
  INV_X1 U13430 ( .A(n20074), .ZN(n20075) );
  INV_X1 U13431 ( .A(matrix_mul_2D_4__5__17_), .ZN(n20076) );
  INV_X1 U13432 ( .A(n20076), .ZN(n20077) );
  INV_X1 U13433 ( .A(matrix_mul_2D_4__5__16_), .ZN(n20078) );
  INV_X1 U13434 ( .A(n20078), .ZN(n20079) );
  INV_X1 U13435 ( .A(matrix_mul_2D_4__5__15_), .ZN(n20080) );
  INV_X1 U13436 ( .A(n20080), .ZN(n20081) );
  INV_X1 U13437 ( .A(matrix_mul_2D_4__4__20_), .ZN(n20082) );
  INV_X1 U13438 ( .A(n20082), .ZN(n20083) );
  INV_X1 U13439 ( .A(matrix_mul_2D_4__4__19_), .ZN(n20084) );
  INV_X1 U13440 ( .A(n20084), .ZN(n20085) );
  INV_X1 U13441 ( .A(matrix_mul_2D_4__4__18_), .ZN(n20086) );
  INV_X1 U13442 ( .A(n20086), .ZN(n20087) );
  INV_X1 U13443 ( .A(matrix_mul_2D_4__4__17_), .ZN(n20088) );
  INV_X1 U13444 ( .A(n20088), .ZN(n20089) );
  INV_X1 U13445 ( .A(matrix_mul_2D_4__4__16_), .ZN(n20090) );
  INV_X1 U13446 ( .A(n20090), .ZN(n20091) );
  INV_X1 U13447 ( .A(matrix_mul_2D_4__4__15_), .ZN(n20092) );
  INV_X1 U13448 ( .A(n20092), .ZN(n20093) );
  INV_X1 U13449 ( .A(matrix_mul_2D_4__3__20_), .ZN(n20094) );
  INV_X1 U13450 ( .A(n20094), .ZN(n20095) );
  INV_X1 U13451 ( .A(matrix_mul_2D_4__3__19_), .ZN(n20096) );
  INV_X1 U13452 ( .A(n20096), .ZN(n20097) );
  INV_X1 U13453 ( .A(matrix_mul_2D_4__3__18_), .ZN(n20098) );
  INV_X1 U13454 ( .A(n20098), .ZN(n20099) );
  INV_X1 U13455 ( .A(matrix_mul_2D_4__3__17_), .ZN(n20100) );
  INV_X1 U13456 ( .A(n20100), .ZN(n20101) );
  INV_X1 U13457 ( .A(matrix_mul_2D_4__3__16_), .ZN(n20102) );
  INV_X1 U13458 ( .A(n20102), .ZN(n20103) );
  INV_X1 U13459 ( .A(matrix_mul_2D_4__3__15_), .ZN(n20104) );
  INV_X1 U13460 ( .A(n20104), .ZN(n20105) );
  INV_X1 U13461 ( .A(matrix_mul_2D_4__2__20_), .ZN(n20106) );
  INV_X1 U13462 ( .A(n20106), .ZN(n20107) );
  INV_X1 U13463 ( .A(matrix_mul_2D_4__2__19_), .ZN(n20108) );
  INV_X1 U13464 ( .A(n20108), .ZN(n20109) );
  INV_X1 U13465 ( .A(matrix_mul_2D_4__2__18_), .ZN(n20110) );
  INV_X1 U13466 ( .A(n20110), .ZN(n20111) );
  INV_X1 U13467 ( .A(matrix_mul_2D_4__2__17_), .ZN(n20112) );
  INV_X1 U13468 ( .A(n20112), .ZN(n20113) );
  INV_X1 U13469 ( .A(matrix_mul_2D_4__2__16_), .ZN(n20114) );
  INV_X1 U13470 ( .A(n20114), .ZN(n20115) );
  INV_X1 U13471 ( .A(matrix_mul_2D_4__2__15_), .ZN(n20116) );
  INV_X1 U13472 ( .A(n20116), .ZN(n20117) );
  INV_X1 U13473 ( .A(matrix_mul_2D_4__1__20_), .ZN(n20118) );
  INV_X1 U13474 ( .A(n20118), .ZN(n20119) );
  INV_X1 U13475 ( .A(matrix_mul_2D_4__1__19_), .ZN(n20120) );
  INV_X1 U13476 ( .A(n20120), .ZN(n20121) );
  INV_X1 U13477 ( .A(matrix_mul_2D_4__1__18_), .ZN(n20122) );
  INV_X1 U13478 ( .A(n20122), .ZN(n20123) );
  INV_X1 U13479 ( .A(matrix_mul_2D_4__1__17_), .ZN(n20124) );
  INV_X1 U13480 ( .A(n20124), .ZN(n20125) );
  INV_X1 U13481 ( .A(matrix_mul_2D_4__1__16_), .ZN(n20126) );
  INV_X1 U13482 ( .A(n20126), .ZN(n20127) );
  INV_X1 U13483 ( .A(matrix_mul_2D_4__1__15_), .ZN(n20128) );
  INV_X1 U13484 ( .A(n20128), .ZN(n20129) );
  INV_X1 U13485 ( .A(matrix_mul_2D_4__0__20_), .ZN(n20130) );
  INV_X1 U13486 ( .A(n20130), .ZN(n20131) );
  INV_X1 U13487 ( .A(matrix_mul_2D_4__0__19_), .ZN(n20132) );
  INV_X1 U13488 ( .A(n20132), .ZN(n20133) );
  INV_X1 U13489 ( .A(matrix_mul_2D_4__0__18_), .ZN(n20134) );
  INV_X1 U13490 ( .A(n20134), .ZN(n20135) );
  INV_X1 U13491 ( .A(matrix_mul_2D_4__0__17_), .ZN(n20136) );
  INV_X1 U13492 ( .A(n20136), .ZN(n20137) );
  INV_X1 U13493 ( .A(matrix_mul_2D_4__0__16_), .ZN(n20138) );
  INV_X1 U13494 ( .A(n20138), .ZN(n20139) );
  INV_X1 U13495 ( .A(matrix_mul_2D_4__0__15_), .ZN(n20140) );
  INV_X1 U13496 ( .A(n20140), .ZN(n20141) );
  INV_X1 U13497 ( .A(matrix_mul_2D_3__7__20_), .ZN(n20142) );
  INV_X1 U13498 ( .A(n20142), .ZN(n20143) );
  INV_X1 U13499 ( .A(matrix_mul_2D_3__7__19_), .ZN(n20144) );
  INV_X1 U13500 ( .A(n20144), .ZN(n20145) );
  INV_X1 U13501 ( .A(matrix_mul_2D_3__7__18_), .ZN(n20146) );
  INV_X1 U13502 ( .A(n20146), .ZN(n20147) );
  INV_X1 U13503 ( .A(matrix_mul_2D_3__7__17_), .ZN(n20148) );
  INV_X1 U13504 ( .A(n20148), .ZN(n20149) );
  INV_X1 U13505 ( .A(matrix_mul_2D_3__7__16_), .ZN(n20150) );
  INV_X1 U13506 ( .A(n20150), .ZN(n20151) );
  INV_X1 U13507 ( .A(matrix_mul_2D_3__7__15_), .ZN(n20152) );
  INV_X1 U13508 ( .A(n20152), .ZN(n20153) );
  INV_X1 U13509 ( .A(matrix_mul_2D_3__6__20_), .ZN(n20154) );
  INV_X1 U13510 ( .A(n20154), .ZN(n20155) );
  INV_X1 U13511 ( .A(matrix_mul_2D_3__6__19_), .ZN(n20156) );
  INV_X1 U13512 ( .A(n20156), .ZN(n20157) );
  INV_X1 U13513 ( .A(matrix_mul_2D_3__6__18_), .ZN(n20158) );
  INV_X1 U13514 ( .A(n20158), .ZN(n20159) );
  INV_X1 U13515 ( .A(matrix_mul_2D_3__6__17_), .ZN(n20160) );
  INV_X1 U13516 ( .A(n20160), .ZN(n20161) );
  INV_X1 U13517 ( .A(matrix_mul_2D_3__6__16_), .ZN(n20162) );
  INV_X1 U13518 ( .A(n20162), .ZN(n20163) );
  INV_X1 U13519 ( .A(matrix_mul_2D_3__6__15_), .ZN(n20164) );
  INV_X1 U13520 ( .A(n20164), .ZN(n20165) );
  INV_X1 U13521 ( .A(matrix_mul_2D_3__5__20_), .ZN(n20166) );
  INV_X1 U13522 ( .A(n20166), .ZN(n20167) );
  INV_X1 U13523 ( .A(matrix_mul_2D_3__5__19_), .ZN(n20168) );
  INV_X1 U13524 ( .A(n20168), .ZN(n20169) );
  INV_X1 U13525 ( .A(matrix_mul_2D_3__5__18_), .ZN(n20170) );
  INV_X1 U13526 ( .A(n20170), .ZN(n20171) );
  INV_X1 U13527 ( .A(matrix_mul_2D_3__5__17_), .ZN(n20172) );
  INV_X1 U13528 ( .A(n20172), .ZN(n20173) );
  INV_X1 U13529 ( .A(matrix_mul_2D_3__5__16_), .ZN(n20174) );
  INV_X1 U13530 ( .A(n20174), .ZN(n20175) );
  INV_X1 U13531 ( .A(matrix_mul_2D_3__5__15_), .ZN(n20176) );
  INV_X1 U13532 ( .A(n20176), .ZN(n20177) );
  INV_X1 U13533 ( .A(matrix_mul_2D_3__4__20_), .ZN(n20178) );
  INV_X1 U13534 ( .A(n20178), .ZN(n20179) );
  INV_X1 U13535 ( .A(matrix_mul_2D_3__4__19_), .ZN(n20180) );
  INV_X1 U13536 ( .A(n20180), .ZN(n20181) );
  INV_X1 U13537 ( .A(matrix_mul_2D_3__4__18_), .ZN(n20182) );
  INV_X1 U13538 ( .A(n20182), .ZN(n20183) );
  INV_X1 U13539 ( .A(matrix_mul_2D_3__4__17_), .ZN(n20184) );
  INV_X1 U13540 ( .A(n20184), .ZN(n20185) );
  INV_X1 U13541 ( .A(matrix_mul_2D_3__4__16_), .ZN(n20186) );
  INV_X1 U13542 ( .A(n20186), .ZN(n20187) );
  INV_X1 U13543 ( .A(matrix_mul_2D_3__4__15_), .ZN(n20188) );
  INV_X1 U13544 ( .A(n20188), .ZN(n20189) );
  INV_X1 U13545 ( .A(matrix_mul_2D_3__3__20_), .ZN(n20190) );
  INV_X1 U13546 ( .A(n20190), .ZN(n20191) );
  INV_X1 U13547 ( .A(matrix_mul_2D_3__3__19_), .ZN(n20192) );
  INV_X1 U13548 ( .A(n20192), .ZN(n20193) );
  INV_X1 U13549 ( .A(matrix_mul_2D_3__3__18_), .ZN(n20194) );
  INV_X1 U13550 ( .A(n20194), .ZN(n20195) );
  INV_X1 U13551 ( .A(matrix_mul_2D_3__3__17_), .ZN(n20196) );
  INV_X1 U13552 ( .A(n20196), .ZN(n20197) );
  INV_X1 U13553 ( .A(matrix_mul_2D_3__3__16_), .ZN(n20198) );
  INV_X1 U13554 ( .A(n20198), .ZN(n20199) );
  INV_X1 U13555 ( .A(matrix_mul_2D_3__3__15_), .ZN(n20200) );
  INV_X1 U13556 ( .A(n20200), .ZN(n20201) );
  INV_X1 U13557 ( .A(matrix_mul_2D_3__2__20_), .ZN(n20202) );
  INV_X1 U13558 ( .A(n20202), .ZN(n20203) );
  INV_X1 U13559 ( .A(matrix_mul_2D_3__2__19_), .ZN(n20204) );
  INV_X1 U13560 ( .A(n20204), .ZN(n20205) );
  INV_X1 U13561 ( .A(matrix_mul_2D_3__2__18_), .ZN(n20206) );
  INV_X1 U13562 ( .A(n20206), .ZN(n20207) );
  INV_X1 U13563 ( .A(matrix_mul_2D_3__2__17_), .ZN(n20208) );
  INV_X1 U13564 ( .A(n20208), .ZN(n20209) );
  INV_X1 U13565 ( .A(matrix_mul_2D_3__2__16_), .ZN(n20210) );
  INV_X1 U13566 ( .A(n20210), .ZN(n20211) );
  INV_X1 U13567 ( .A(matrix_mul_2D_3__2__15_), .ZN(n20212) );
  INV_X1 U13568 ( .A(n20212), .ZN(n20213) );
  INV_X1 U13569 ( .A(matrix_mul_2D_3__1__20_), .ZN(n20214) );
  INV_X1 U13570 ( .A(n20214), .ZN(n20215) );
  INV_X1 U13571 ( .A(matrix_mul_2D_3__1__19_), .ZN(n20216) );
  INV_X1 U13572 ( .A(n20216), .ZN(n20217) );
  INV_X1 U13573 ( .A(matrix_mul_2D_3__1__18_), .ZN(n20218) );
  INV_X1 U13574 ( .A(n20218), .ZN(n20219) );
  INV_X1 U13575 ( .A(matrix_mul_2D_3__1__17_), .ZN(n20220) );
  INV_X1 U13576 ( .A(n20220), .ZN(n20221) );
  INV_X1 U13577 ( .A(matrix_mul_2D_3__1__16_), .ZN(n20222) );
  INV_X1 U13578 ( .A(n20222), .ZN(n20223) );
  INV_X1 U13579 ( .A(matrix_mul_2D_3__1__15_), .ZN(n20224) );
  INV_X1 U13580 ( .A(n20224), .ZN(n20225) );
  INV_X1 U13581 ( .A(matrix_mul_2D_3__0__20_), .ZN(n20226) );
  INV_X1 U13582 ( .A(n20226), .ZN(n20227) );
  INV_X1 U13583 ( .A(matrix_mul_2D_3__0__19_), .ZN(n20228) );
  INV_X1 U13584 ( .A(n20228), .ZN(n20229) );
  INV_X1 U13585 ( .A(matrix_mul_2D_3__0__18_), .ZN(n20230) );
  INV_X1 U13586 ( .A(n20230), .ZN(n20231) );
  INV_X1 U13587 ( .A(matrix_mul_2D_3__0__17_), .ZN(n20232) );
  INV_X1 U13588 ( .A(n20232), .ZN(n20233) );
  INV_X1 U13589 ( .A(matrix_mul_2D_3__0__16_), .ZN(n20234) );
  INV_X1 U13590 ( .A(n20234), .ZN(n20235) );
  INV_X1 U13591 ( .A(matrix_mul_2D_3__0__15_), .ZN(n20236) );
  INV_X1 U13592 ( .A(n20236), .ZN(n20237) );
  INV_X1 U13593 ( .A(matrix_mul_2D_2__7__20_), .ZN(n20238) );
  INV_X1 U13594 ( .A(n20238), .ZN(n20239) );
  INV_X1 U13595 ( .A(matrix_mul_2D_2__7__19_), .ZN(n20240) );
  INV_X1 U13596 ( .A(n20240), .ZN(n20241) );
  INV_X1 U13597 ( .A(matrix_mul_2D_2__7__18_), .ZN(n20242) );
  INV_X1 U13598 ( .A(n20242), .ZN(n20243) );
  INV_X1 U13599 ( .A(matrix_mul_2D_2__7__17_), .ZN(n20244) );
  INV_X1 U13600 ( .A(n20244), .ZN(n20245) );
  INV_X1 U13601 ( .A(matrix_mul_2D_2__7__16_), .ZN(n20246) );
  INV_X1 U13602 ( .A(n20246), .ZN(n20247) );
  INV_X1 U13603 ( .A(matrix_mul_2D_2__7__15_), .ZN(n20248) );
  INV_X1 U13604 ( .A(n20248), .ZN(n20249) );
  INV_X1 U13605 ( .A(matrix_mul_2D_2__6__20_), .ZN(n20250) );
  INV_X1 U13606 ( .A(n20250), .ZN(n20251) );
  INV_X1 U13607 ( .A(matrix_mul_2D_2__6__19_), .ZN(n20252) );
  INV_X1 U13608 ( .A(n20252), .ZN(n20253) );
  INV_X1 U13609 ( .A(matrix_mul_2D_2__6__18_), .ZN(n20254) );
  INV_X1 U13610 ( .A(n20254), .ZN(n20255) );
  INV_X1 U13611 ( .A(matrix_mul_2D_2__6__17_), .ZN(n20256) );
  INV_X1 U13612 ( .A(n20256), .ZN(n20257) );
  INV_X1 U13613 ( .A(matrix_mul_2D_2__6__16_), .ZN(n20258) );
  INV_X1 U13614 ( .A(n20258), .ZN(n20259) );
  INV_X1 U13615 ( .A(matrix_mul_2D_2__6__15_), .ZN(n20260) );
  INV_X1 U13616 ( .A(n20260), .ZN(n20261) );
  INV_X1 U13617 ( .A(matrix_mul_2D_2__5__20_), .ZN(n20262) );
  INV_X1 U13618 ( .A(n20262), .ZN(n20263) );
  INV_X1 U13619 ( .A(matrix_mul_2D_2__5__19_), .ZN(n20264) );
  INV_X1 U13620 ( .A(n20264), .ZN(n20265) );
  INV_X1 U13621 ( .A(matrix_mul_2D_2__5__18_), .ZN(n20266) );
  INV_X1 U13622 ( .A(n20266), .ZN(n20267) );
  INV_X1 U13623 ( .A(matrix_mul_2D_2__5__17_), .ZN(n20268) );
  INV_X1 U13624 ( .A(n20268), .ZN(n20269) );
  INV_X1 U13625 ( .A(matrix_mul_2D_2__5__16_), .ZN(n20270) );
  INV_X1 U13626 ( .A(n20270), .ZN(n20271) );
  INV_X1 U13627 ( .A(matrix_mul_2D_2__5__15_), .ZN(n20272) );
  INV_X1 U13628 ( .A(n20272), .ZN(n20273) );
  INV_X1 U13629 ( .A(matrix_mul_2D_2__4__20_), .ZN(n20274) );
  INV_X1 U13630 ( .A(n20274), .ZN(n20275) );
  INV_X1 U13631 ( .A(matrix_mul_2D_2__4__19_), .ZN(n20276) );
  INV_X1 U13632 ( .A(n20276), .ZN(n20277) );
  INV_X1 U13633 ( .A(matrix_mul_2D_2__4__18_), .ZN(n20278) );
  INV_X1 U13634 ( .A(n20278), .ZN(n20279) );
  INV_X1 U13635 ( .A(matrix_mul_2D_2__4__17_), .ZN(n20280) );
  INV_X1 U13636 ( .A(n20280), .ZN(n20281) );
  INV_X1 U13637 ( .A(matrix_mul_2D_2__4__16_), .ZN(n20282) );
  INV_X1 U13638 ( .A(n20282), .ZN(n20283) );
  INV_X1 U13639 ( .A(matrix_mul_2D_2__4__15_), .ZN(n20284) );
  INV_X1 U13640 ( .A(n20284), .ZN(n20285) );
  INV_X1 U13641 ( .A(matrix_mul_2D_2__3__20_), .ZN(n20286) );
  INV_X1 U13642 ( .A(n20286), .ZN(n20287) );
  INV_X1 U13643 ( .A(matrix_mul_2D_2__3__19_), .ZN(n20288) );
  INV_X1 U13644 ( .A(n20288), .ZN(n20289) );
  INV_X1 U13645 ( .A(matrix_mul_2D_2__3__18_), .ZN(n20290) );
  INV_X1 U13646 ( .A(n20290), .ZN(n20291) );
  INV_X1 U13647 ( .A(matrix_mul_2D_2__3__17_), .ZN(n20292) );
  INV_X1 U13648 ( .A(n20292), .ZN(n20293) );
  INV_X1 U13649 ( .A(matrix_mul_2D_2__3__16_), .ZN(n20294) );
  INV_X1 U13650 ( .A(n20294), .ZN(n20295) );
  INV_X1 U13651 ( .A(matrix_mul_2D_2__3__15_), .ZN(n20296) );
  INV_X1 U13652 ( .A(n20296), .ZN(n20297) );
  INV_X1 U13653 ( .A(matrix_mul_2D_2__2__20_), .ZN(n20298) );
  INV_X1 U13654 ( .A(n20298), .ZN(n20299) );
  INV_X1 U13655 ( .A(matrix_mul_2D_2__2__19_), .ZN(n20300) );
  INV_X1 U13656 ( .A(n20300), .ZN(n20301) );
  INV_X1 U13657 ( .A(matrix_mul_2D_2__2__18_), .ZN(n20302) );
  INV_X1 U13658 ( .A(n20302), .ZN(n20303) );
  INV_X1 U13659 ( .A(matrix_mul_2D_2__2__17_), .ZN(n20304) );
  INV_X1 U13660 ( .A(n20304), .ZN(n20305) );
  INV_X1 U13661 ( .A(matrix_mul_2D_2__2__16_), .ZN(n20306) );
  INV_X1 U13662 ( .A(n20306), .ZN(n20307) );
  INV_X1 U13663 ( .A(matrix_mul_2D_2__2__15_), .ZN(n20308) );
  INV_X1 U13664 ( .A(n20308), .ZN(n20309) );
  INV_X1 U13665 ( .A(matrix_mul_2D_2__1__20_), .ZN(n20310) );
  INV_X1 U13666 ( .A(n20310), .ZN(n20311) );
  INV_X1 U13667 ( .A(matrix_mul_2D_2__1__19_), .ZN(n20312) );
  INV_X1 U13668 ( .A(n20312), .ZN(n20313) );
  INV_X1 U13669 ( .A(matrix_mul_2D_2__1__18_), .ZN(n20314) );
  INV_X1 U13670 ( .A(n20314), .ZN(n20315) );
  INV_X1 U13671 ( .A(matrix_mul_2D_2__1__17_), .ZN(n20316) );
  INV_X1 U13672 ( .A(n20316), .ZN(n20317) );
  INV_X1 U13673 ( .A(matrix_mul_2D_2__1__16_), .ZN(n20318) );
  INV_X1 U13674 ( .A(n20318), .ZN(n20319) );
  INV_X1 U13675 ( .A(matrix_mul_2D_2__1__15_), .ZN(n20320) );
  INV_X1 U13676 ( .A(n20320), .ZN(n20321) );
  INV_X1 U13677 ( .A(matrix_mul_2D_2__0__20_), .ZN(n20322) );
  INV_X1 U13678 ( .A(n20322), .ZN(n20323) );
  INV_X1 U13679 ( .A(matrix_mul_2D_2__0__19_), .ZN(n20324) );
  INV_X1 U13680 ( .A(n20324), .ZN(n20325) );
  INV_X1 U13681 ( .A(matrix_mul_2D_2__0__18_), .ZN(n20326) );
  INV_X1 U13682 ( .A(n20326), .ZN(n20327) );
  INV_X1 U13683 ( .A(matrix_mul_2D_2__0__17_), .ZN(n20328) );
  INV_X1 U13684 ( .A(n20328), .ZN(n20329) );
  INV_X1 U13685 ( .A(matrix_mul_2D_2__0__16_), .ZN(n20330) );
  INV_X1 U13686 ( .A(n20330), .ZN(n20331) );
  INV_X1 U13687 ( .A(matrix_mul_2D_2__0__15_), .ZN(n20332) );
  INV_X1 U13688 ( .A(n20332), .ZN(n20333) );
  INV_X1 U13689 ( .A(matrix_mul_2D_1__7__20_), .ZN(n20334) );
  INV_X1 U13690 ( .A(n20334), .ZN(n20335) );
  INV_X1 U13691 ( .A(matrix_mul_2D_1__7__19_), .ZN(n20336) );
  INV_X1 U13692 ( .A(n20336), .ZN(n20337) );
  INV_X1 U13693 ( .A(matrix_mul_2D_1__7__18_), .ZN(n20338) );
  INV_X1 U13694 ( .A(n20338), .ZN(n20339) );
  INV_X1 U13695 ( .A(matrix_mul_2D_1__7__17_), .ZN(n20340) );
  INV_X1 U13696 ( .A(n20340), .ZN(n20341) );
  INV_X1 U13697 ( .A(matrix_mul_2D_1__7__16_), .ZN(n20342) );
  INV_X1 U13698 ( .A(n20342), .ZN(n20343) );
  INV_X1 U13699 ( .A(matrix_mul_2D_1__7__15_), .ZN(n20344) );
  INV_X1 U13700 ( .A(n20344), .ZN(n20345) );
  INV_X1 U13701 ( .A(matrix_mul_2D_1__6__20_), .ZN(n20346) );
  INV_X1 U13702 ( .A(n20346), .ZN(n20347) );
  INV_X1 U13703 ( .A(matrix_mul_2D_1__6__19_), .ZN(n20348) );
  INV_X1 U13704 ( .A(n20348), .ZN(n20349) );
  INV_X1 U13705 ( .A(matrix_mul_2D_1__6__18_), .ZN(n20350) );
  INV_X1 U13706 ( .A(n20350), .ZN(n20351) );
  INV_X1 U13707 ( .A(matrix_mul_2D_1__6__17_), .ZN(n20352) );
  INV_X1 U13708 ( .A(n20352), .ZN(n20353) );
  INV_X1 U13709 ( .A(matrix_mul_2D_1__6__16_), .ZN(n20354) );
  INV_X1 U13710 ( .A(n20354), .ZN(n20355) );
  INV_X1 U13711 ( .A(matrix_mul_2D_1__6__15_), .ZN(n20356) );
  INV_X1 U13712 ( .A(n20356), .ZN(n20357) );
  INV_X1 U13713 ( .A(matrix_mul_2D_1__1__20_), .ZN(n20358) );
  INV_X1 U13714 ( .A(n20358), .ZN(n20359) );
  INV_X1 U13715 ( .A(matrix_mul_2D_1__1__19_), .ZN(n20360) );
  INV_X1 U13716 ( .A(n20360), .ZN(n20361) );
  INV_X1 U13717 ( .A(matrix_mul_2D_1__1__18_), .ZN(n20362) );
  INV_X1 U13718 ( .A(n20362), .ZN(n20363) );
  INV_X1 U13719 ( .A(matrix_mul_2D_1__1__17_), .ZN(n20364) );
  INV_X1 U13720 ( .A(n20364), .ZN(n20365) );
  INV_X1 U13721 ( .A(matrix_mul_2D_1__1__16_), .ZN(n20366) );
  INV_X1 U13722 ( .A(n20366), .ZN(n20367) );
  INV_X1 U13723 ( .A(matrix_mul_2D_1__1__15_), .ZN(n20368) );
  INV_X1 U13724 ( .A(n20368), .ZN(n20369) );
  INV_X1 U13725 ( .A(matrix_mul_2D_1__0__20_), .ZN(n20370) );
  INV_X1 U13726 ( .A(n20370), .ZN(n20371) );
  INV_X1 U13727 ( .A(matrix_mul_2D_1__0__19_), .ZN(n20372) );
  INV_X1 U13728 ( .A(n20372), .ZN(n20373) );
  INV_X1 U13729 ( .A(matrix_mul_2D_1__0__18_), .ZN(n20374) );
  INV_X1 U13730 ( .A(n20374), .ZN(n20375) );
  INV_X1 U13731 ( .A(matrix_mul_2D_1__0__17_), .ZN(n20376) );
  INV_X1 U13732 ( .A(n20376), .ZN(n20377) );
  INV_X1 U13733 ( .A(matrix_mul_2D_1__0__16_), .ZN(n20378) );
  INV_X1 U13734 ( .A(n20378), .ZN(n20379) );
  INV_X1 U13735 ( .A(matrix_mul_2D_1__0__15_), .ZN(n20380) );
  INV_X1 U13736 ( .A(n20380), .ZN(n20381) );
  INV_X1 U13737 ( .A(matrix_mul_2D_0__7__20_), .ZN(n20382) );
  INV_X1 U13738 ( .A(n20382), .ZN(n20383) );
  INV_X1 U13739 ( .A(matrix_mul_2D_0__7__19_), .ZN(n20384) );
  INV_X1 U13740 ( .A(n20384), .ZN(n20385) );
  INV_X1 U13741 ( .A(matrix_mul_2D_0__7__18_), .ZN(n20386) );
  INV_X1 U13742 ( .A(n20386), .ZN(n20387) );
  INV_X1 U13743 ( .A(matrix_mul_2D_0__7__17_), .ZN(n20388) );
  INV_X1 U13744 ( .A(n20388), .ZN(n20389) );
  INV_X1 U13745 ( .A(matrix_mul_2D_0__7__16_), .ZN(n20390) );
  INV_X1 U13746 ( .A(n20390), .ZN(n20391) );
  INV_X1 U13747 ( .A(matrix_mul_2D_0__7__15_), .ZN(n20392) );
  INV_X1 U13748 ( .A(n20392), .ZN(n20393) );
  INV_X1 U13749 ( .A(matrix_mul_2D_0__6__20_), .ZN(n20394) );
  INV_X1 U13750 ( .A(n20394), .ZN(n20395) );
  INV_X1 U13751 ( .A(matrix_mul_2D_0__6__19_), .ZN(n20396) );
  INV_X1 U13752 ( .A(n20396), .ZN(n20397) );
  INV_X1 U13753 ( .A(matrix_mul_2D_0__6__18_), .ZN(n20398) );
  INV_X1 U13754 ( .A(n20398), .ZN(n20399) );
  INV_X1 U13755 ( .A(matrix_mul_2D_0__6__17_), .ZN(n20400) );
  INV_X1 U13756 ( .A(n20400), .ZN(n20401) );
  INV_X1 U13757 ( .A(matrix_mul_2D_0__6__16_), .ZN(n20402) );
  INV_X1 U13758 ( .A(n20402), .ZN(n20403) );
  INV_X1 U13759 ( .A(matrix_mul_2D_0__6__15_), .ZN(n20404) );
  INV_X1 U13760 ( .A(n20404), .ZN(n20405) );
  INV_X1 U13761 ( .A(matrix_mul_2D_0__5__20_), .ZN(n20406) );
  INV_X1 U13762 ( .A(n20406), .ZN(n20407) );
  INV_X1 U13763 ( .A(matrix_mul_2D_0__5__19_), .ZN(n20408) );
  INV_X1 U13764 ( .A(n20408), .ZN(n20409) );
  INV_X1 U13765 ( .A(matrix_mul_2D_0__5__18_), .ZN(n20410) );
  INV_X1 U13766 ( .A(n20410), .ZN(n20411) );
  INV_X1 U13767 ( .A(matrix_mul_2D_0__5__17_), .ZN(n20412) );
  INV_X1 U13768 ( .A(n20412), .ZN(n20413) );
  INV_X1 U13769 ( .A(matrix_mul_2D_0__5__16_), .ZN(n20414) );
  INV_X1 U13770 ( .A(n20414), .ZN(n20415) );
  INV_X1 U13771 ( .A(matrix_mul_2D_0__5__15_), .ZN(n20416) );
  INV_X1 U13772 ( .A(n20416), .ZN(n20417) );
  INV_X1 U13773 ( .A(matrix_mul_2D_0__4__20_), .ZN(n20418) );
  INV_X1 U13774 ( .A(n20418), .ZN(n20419) );
  INV_X1 U13775 ( .A(matrix_mul_2D_0__4__19_), .ZN(n20420) );
  INV_X1 U13776 ( .A(n20420), .ZN(n20421) );
  INV_X1 U13777 ( .A(matrix_mul_2D_0__4__18_), .ZN(n20422) );
  INV_X1 U13778 ( .A(n20422), .ZN(n20423) );
  INV_X1 U13779 ( .A(matrix_mul_2D_0__4__17_), .ZN(n20424) );
  INV_X1 U13780 ( .A(n20424), .ZN(n20425) );
  INV_X1 U13781 ( .A(matrix_mul_2D_0__4__16_), .ZN(n20426) );
  INV_X1 U13782 ( .A(n20426), .ZN(n20427) );
  INV_X1 U13783 ( .A(matrix_mul_2D_0__4__15_), .ZN(n20428) );
  INV_X1 U13784 ( .A(n20428), .ZN(n20429) );
  INV_X1 U13785 ( .A(matrix_mul_2D_0__3__20_), .ZN(n20430) );
  INV_X1 U13786 ( .A(n20430), .ZN(n20431) );
  INV_X1 U13787 ( .A(matrix_mul_2D_0__3__19_), .ZN(n20432) );
  INV_X1 U13788 ( .A(n20432), .ZN(n20433) );
  INV_X1 U13789 ( .A(matrix_mul_2D_0__3__18_), .ZN(n20434) );
  INV_X1 U13790 ( .A(n20434), .ZN(n20435) );
  INV_X1 U13791 ( .A(matrix_mul_2D_0__3__17_), .ZN(n20436) );
  INV_X1 U13792 ( .A(n20436), .ZN(n20437) );
  INV_X1 U13793 ( .A(matrix_mul_2D_0__3__16_), .ZN(n20438) );
  INV_X1 U13794 ( .A(n20438), .ZN(n20439) );
  INV_X1 U13795 ( .A(matrix_mul_2D_0__3__15_), .ZN(n20440) );
  INV_X1 U13796 ( .A(n20440), .ZN(n20441) );
  INV_X1 U13797 ( .A(matrix_mul_2D_0__2__20_), .ZN(n20442) );
  INV_X1 U13798 ( .A(n20442), .ZN(n20443) );
  INV_X1 U13799 ( .A(matrix_mul_2D_0__2__19_), .ZN(n20444) );
  INV_X1 U13800 ( .A(n20444), .ZN(n20445) );
  INV_X1 U13801 ( .A(matrix_mul_2D_0__2__18_), .ZN(n20446) );
  INV_X1 U13802 ( .A(n20446), .ZN(n20447) );
  INV_X1 U13803 ( .A(matrix_mul_2D_0__2__17_), .ZN(n20448) );
  INV_X1 U13804 ( .A(n20448), .ZN(n20449) );
  INV_X1 U13805 ( .A(matrix_mul_2D_0__2__16_), .ZN(n20450) );
  INV_X1 U13806 ( .A(n20450), .ZN(n20451) );
  INV_X1 U13807 ( .A(matrix_mul_2D_0__2__15_), .ZN(n20452) );
  INV_X1 U13808 ( .A(n20452), .ZN(n20453) );
  INV_X1 U13809 ( .A(matrix_mul_2D_0__1__20_), .ZN(n20454) );
  INV_X1 U13810 ( .A(n20454), .ZN(n20455) );
  INV_X1 U13811 ( .A(matrix_mul_2D_0__1__19_), .ZN(n20456) );
  INV_X1 U13812 ( .A(n20456), .ZN(n20457) );
  INV_X1 U13813 ( .A(matrix_mul_2D_0__1__18_), .ZN(n20458) );
  INV_X1 U13814 ( .A(n20458), .ZN(n20459) );
  INV_X1 U13815 ( .A(matrix_mul_2D_0__1__17_), .ZN(n20460) );
  INV_X1 U13816 ( .A(n20460), .ZN(n20461) );
  INV_X1 U13817 ( .A(matrix_mul_2D_0__1__16_), .ZN(n20462) );
  INV_X1 U13818 ( .A(n20462), .ZN(n20463) );
  INV_X1 U13819 ( .A(matrix_mul_2D_0__1__15_), .ZN(n20464) );
  INV_X1 U13820 ( .A(n20464), .ZN(n20465) );
  INV_X1 U13821 ( .A(matrix_mul_2D_0__0__20_), .ZN(n20466) );
  INV_X1 U13822 ( .A(n20466), .ZN(n20467) );
  INV_X1 U13823 ( .A(matrix_mul_2D_0__0__19_), .ZN(n20468) );
  INV_X1 U13824 ( .A(n20468), .ZN(n20469) );
  INV_X1 U13825 ( .A(matrix_mul_2D_0__0__18_), .ZN(n20470) );
  INV_X1 U13826 ( .A(n20470), .ZN(n20471) );
  INV_X1 U13827 ( .A(matrix_mul_2D_0__0__17_), .ZN(n20472) );
  INV_X1 U13828 ( .A(n20472), .ZN(n20473) );
  INV_X1 U13829 ( .A(matrix_mul_2D_0__0__16_), .ZN(n20474) );
  INV_X1 U13830 ( .A(n20474), .ZN(n20475) );
  INV_X1 U13831 ( .A(matrix_mul_2D_0__0__15_), .ZN(n20476) );
  INV_X1 U13832 ( .A(n20476), .ZN(n20477) );
  INV_X1 U13833 ( .A(n4989), .ZN(n20478) );
  INV_X1 U13834 ( .A(n20478), .ZN(n20479) );
  INV_X1 U13835 ( .A(n20478), .ZN(n20480) );
  INV_X1 U13836 ( .A(n20961), .ZN(n20481) );
  INV_X1 U13837 ( .A(n4990), .ZN(n20482) );
  INV_X1 U13838 ( .A(n20482), .ZN(n20483) );
  INV_X1 U13839 ( .A(n20482), .ZN(n20484) );
  INV_X1 U13840 ( .A(n4985), .ZN(n20485) );
  INV_X1 U13841 ( .A(n20485), .ZN(n20486) );
  INV_X1 U13842 ( .A(n20485), .ZN(n20487) );
  INV_X1 U13843 ( .A(n17991), .ZN(n20488) );
  INV_X1 U13844 ( .A(n17991), .ZN(n20489) );
  INV_X1 U13845 ( .A(n47890), .ZN(n20490) );
  INV_X1 U13846 ( .A(n20490), .ZN(n20491) );
  INV_X1 U13847 ( .A(n20490), .ZN(n20492) );
  INV_X1 U13848 ( .A(n17993), .ZN(n20493) );
  INV_X1 U13849 ( .A(n17993), .ZN(n20494) );
  BUF_X1 U13850 ( .A(n3098), .Z(n27110) );
  INV_X1 U13851 ( .A(n17994), .ZN(n20495) );
  INV_X1 U13852 ( .A(n17994), .ZN(n20496) );
  INV_X1 U13853 ( .A(n17995), .ZN(n20497) );
  INV_X1 U13854 ( .A(n17995), .ZN(n20498) );
  INV_X1 U13855 ( .A(n23389), .ZN(n20499) );
  INV_X1 U13856 ( .A(n20499), .ZN(n20500) );
  INV_X1 U13857 ( .A(n20499), .ZN(n20501) );
  INV_X1 U13858 ( .A(n23411), .ZN(n20502) );
  INV_X1 U13859 ( .A(n20502), .ZN(n20503) );
  INV_X1 U13860 ( .A(n20502), .ZN(n20504) );
  INV_X1 U13861 ( .A(n18000), .ZN(n20505) );
  INV_X1 U13862 ( .A(n18000), .ZN(n20506) );
  INV_X1 U13863 ( .A(n18001), .ZN(n20507) );
  INV_X1 U13864 ( .A(n20906), .ZN(n20508) );
  INV_X1 U13865 ( .A(n20508), .ZN(n20509) );
  INV_X1 U13866 ( .A(n20508), .ZN(n20510) );
  INV_X1 U13867 ( .A(n18002), .ZN(n20511) );
  INV_X1 U13868 ( .A(n20901), .ZN(n20512) );
  INV_X1 U13869 ( .A(n20512), .ZN(n20513) );
  INV_X1 U13870 ( .A(n20512), .ZN(n20514) );
  INV_X1 U13871 ( .A(n27275), .ZN(n20515) );
  INV_X1 U13872 ( .A(n20515), .ZN(n20516) );
  INV_X1 U13873 ( .A(n20515), .ZN(n20517) );
  INV_X1 U13874 ( .A(n18003), .ZN(n20518) );
  INV_X1 U13875 ( .A(n18003), .ZN(n20519) );
  INV_X1 U13876 ( .A(n27127), .ZN(n20520) );
  INV_X1 U13877 ( .A(n20520), .ZN(n20521) );
  INV_X1 U13878 ( .A(n20520), .ZN(n20522) );
  INV_X1 U13879 ( .A(n18004), .ZN(n20523) );
  INV_X1 U13880 ( .A(n18004), .ZN(n20524) );
  INV_X1 U13881 ( .A(n18005), .ZN(n20525) );
  INV_X1 U13882 ( .A(n18005), .ZN(n20526) );
  INV_X1 U13883 ( .A(n27127), .ZN(n20527) );
  INV_X1 U13884 ( .A(n20527), .ZN(n20528) );
  INV_X1 U13885 ( .A(n20527), .ZN(n20529) );
  INV_X1 U13886 ( .A(n27275), .ZN(n20530) );
  INV_X1 U13887 ( .A(n20530), .ZN(n20531) );
  INV_X1 U13888 ( .A(n20530), .ZN(n20532) );
  INV_X1 U13889 ( .A(n27126), .ZN(n20533) );
  INV_X1 U13890 ( .A(n20533), .ZN(n20534) );
  INV_X1 U13891 ( .A(n20533), .ZN(n20535) );
  INV_X1 U13892 ( .A(n27274), .ZN(n20536) );
  INV_X1 U13893 ( .A(n20536), .ZN(n20537) );
  INV_X1 U13894 ( .A(n20536), .ZN(n20538) );
  INV_X1 U13895 ( .A(n18006), .ZN(n20539) );
  INV_X1 U13896 ( .A(n18006), .ZN(n20540) );
  INV_X1 U13897 ( .A(n27219), .ZN(n20541) );
  INV_X1 U13898 ( .A(n20541), .ZN(n20542) );
  INV_X1 U13899 ( .A(n20541), .ZN(n20543) );
  INV_X1 U13900 ( .A(n18007), .ZN(n20544) );
  INV_X1 U13901 ( .A(n18007), .ZN(n20545) );
  INV_X1 U13902 ( .A(n18008), .ZN(n20546) );
  INV_X1 U13903 ( .A(n18008), .ZN(n20547) );
  INV_X1 U13904 ( .A(n18009), .ZN(n20548) );
  INV_X1 U13905 ( .A(n18009), .ZN(n20549) );
  INV_X1 U13906 ( .A(n18010), .ZN(n20550) );
  INV_X1 U13907 ( .A(n18010), .ZN(n20551) );
  INV_X1 U13908 ( .A(n24757), .ZN(n20552) );
  INV_X1 U13909 ( .A(n20552), .ZN(n20553) );
  INV_X1 U13910 ( .A(n20552), .ZN(n20554) );
  INV_X1 U13911 ( .A(n27197), .ZN(n20555) );
  INV_X1 U13912 ( .A(n20555), .ZN(n20556) );
  INV_X1 U13913 ( .A(n18949), .ZN(n20557) );
  INV_X1 U13914 ( .A(n20557), .ZN(n20558) );
  INV_X1 U13915 ( .A(n20557), .ZN(n20559) );
  INV_X1 U13916 ( .A(n18011), .ZN(n20560) );
  INV_X1 U13917 ( .A(n18011), .ZN(n20561) );
  INV_X1 U13918 ( .A(n18950), .ZN(n20562) );
  INV_X1 U13919 ( .A(n20562), .ZN(n20563) );
  INV_X1 U13920 ( .A(n20562), .ZN(n20564) );
  INV_X1 U13921 ( .A(n18012), .ZN(n20565) );
  INV_X1 U13922 ( .A(n18012), .ZN(n20566) );
  INV_X1 U13923 ( .A(n18013), .ZN(n20567) );
  INV_X1 U13924 ( .A(n18013), .ZN(n20568) );
  INV_X1 U13925 ( .A(n24768), .ZN(n20569) );
  INV_X1 U13926 ( .A(n20569), .ZN(n20570) );
  INV_X1 U13927 ( .A(n20569), .ZN(n20571) );
  INV_X1 U13928 ( .A(n18014), .ZN(n20572) );
  INV_X1 U13929 ( .A(n18014), .ZN(n20573) );
  INV_X1 U13930 ( .A(n24773), .ZN(n20574) );
  INV_X1 U13931 ( .A(n20574), .ZN(n20575) );
  INV_X1 U13932 ( .A(n20574), .ZN(n20576) );
  INV_X1 U13933 ( .A(n27209), .ZN(n20577) );
  INV_X1 U13934 ( .A(n20577), .ZN(n20578) );
  INV_X1 U13935 ( .A(n20577), .ZN(n20579) );
  INV_X1 U13936 ( .A(n18015), .ZN(n20580) );
  INV_X1 U13937 ( .A(n18015), .ZN(n20581) );
  INV_X1 U13938 ( .A(n18016), .ZN(n20582) );
  INV_X1 U13939 ( .A(n18016), .ZN(n20583) );
  CLKBUF_X1 U13940 ( .A(n24782), .Z(n20584) );
  INV_X1 U13941 ( .A(n18017), .ZN(n20585) );
  INV_X1 U13942 ( .A(n18017), .ZN(n20586) );
  INV_X1 U13943 ( .A(n18018), .ZN(n20587) );
  INV_X1 U13944 ( .A(n18018), .ZN(n20588) );
  INV_X1 U13945 ( .A(n18019), .ZN(n20589) );
  INV_X1 U13946 ( .A(n18019), .ZN(n20590) );
  INV_X1 U13947 ( .A(n18020), .ZN(n20591) );
  INV_X1 U13948 ( .A(n18020), .ZN(n20592) );
  INV_X1 U13949 ( .A(n18021), .ZN(n20593) );
  INV_X1 U13950 ( .A(n18021), .ZN(n20594) );
  INV_X1 U13951 ( .A(n18022), .ZN(n20595) );
  INV_X1 U13952 ( .A(n18022), .ZN(n20596) );
  INV_X1 U13953 ( .A(n18023), .ZN(n20597) );
  INV_X1 U13954 ( .A(n18023), .ZN(n20598) );
  INV_X1 U13955 ( .A(n18024), .ZN(n20599) );
  INV_X1 U13956 ( .A(n18024), .ZN(n20600) );
  INV_X1 U13957 ( .A(n18025), .ZN(n20601) );
  INV_X1 U13958 ( .A(n18025), .ZN(n20602) );
  INV_X1 U13959 ( .A(n18026), .ZN(n20603) );
  INV_X1 U13960 ( .A(n18026), .ZN(n20604) );
  INV_X1 U13961 ( .A(n18027), .ZN(n20605) );
  INV_X1 U13962 ( .A(n18027), .ZN(n20606) );
  INV_X1 U13963 ( .A(n18028), .ZN(n20607) );
  INV_X1 U13964 ( .A(n18028), .ZN(n20608) );
  INV_X1 U13965 ( .A(n20608), .ZN(n20609) );
  INV_X1 U13966 ( .A(n18955), .ZN(n20610) );
  INV_X1 U13967 ( .A(n18029), .ZN(n20611) );
  INV_X1 U13968 ( .A(n18029), .ZN(n20612) );
  INV_X1 U13969 ( .A(n18030), .ZN(n20613) );
  INV_X1 U13970 ( .A(n18030), .ZN(n20614) );
  INV_X1 U13971 ( .A(n18031), .ZN(n20615) );
  INV_X1 U13972 ( .A(n18031), .ZN(n20616) );
  INV_X1 U13973 ( .A(n18032), .ZN(n20617) );
  INV_X1 U13974 ( .A(n18032), .ZN(n20618) );
  INV_X1 U13975 ( .A(n18033), .ZN(n20619) );
  INV_X1 U13976 ( .A(n18033), .ZN(n20620) );
  INV_X1 U13977 ( .A(n18034), .ZN(n20621) );
  INV_X1 U13978 ( .A(n451), .ZN(n20622) );
  INV_X1 U13979 ( .A(n451), .ZN(n20623) );
  INV_X1 U13980 ( .A(n450), .ZN(n20624) );
  INV_X1 U13981 ( .A(n450), .ZN(n20625) );
  INV_X1 U13982 ( .A(n18035), .ZN(n20626) );
  INV_X1 U13983 ( .A(n18035), .ZN(n20627) );
  INV_X1 U13984 ( .A(n449), .ZN(n20628) );
  INV_X1 U13985 ( .A(n449), .ZN(n20629) );
  INV_X1 U13986 ( .A(n448), .ZN(n20630) );
  INV_X1 U13987 ( .A(n448), .ZN(n20631) );
  INV_X1 U13988 ( .A(n447), .ZN(n20632) );
  INV_X1 U13989 ( .A(n447), .ZN(n20633) );
  INV_X1 U13990 ( .A(n18036), .ZN(n20634) );
  INV_X1 U13991 ( .A(n18036), .ZN(n20635) );
  INV_X1 U13992 ( .A(n446), .ZN(n20636) );
  INV_X1 U13993 ( .A(n446), .ZN(n20637) );
  INV_X1 U13994 ( .A(n445), .ZN(n20638) );
  INV_X1 U13995 ( .A(n445), .ZN(n20639) );
  INV_X1 U13996 ( .A(n24832), .ZN(n20640) );
  INV_X1 U13997 ( .A(n20640), .ZN(n20641) );
  INV_X1 U13998 ( .A(n20640), .ZN(n20642) );
  INV_X1 U13999 ( .A(n18037), .ZN(n20643) );
  INV_X1 U14000 ( .A(n18037), .ZN(n20644) );
  INV_X1 U14001 ( .A(n444), .ZN(n20645) );
  INV_X1 U14002 ( .A(n444), .ZN(n20646) );
  INV_X1 U14003 ( .A(n443), .ZN(n20647) );
  INV_X1 U14004 ( .A(n443), .ZN(n20648) );
  INV_X1 U14005 ( .A(n442), .ZN(n20649) );
  INV_X1 U14006 ( .A(n442), .ZN(n20650) );
  INV_X1 U14007 ( .A(n18038), .ZN(n20651) );
  INV_X1 U14008 ( .A(n18038), .ZN(n20652) );
  INV_X1 U14009 ( .A(n441), .ZN(n20653) );
  INV_X1 U14010 ( .A(n441), .ZN(n20654) );
  INV_X1 U14011 ( .A(n440), .ZN(n20655) );
  INV_X1 U14012 ( .A(n440), .ZN(n20656) );
  INV_X1 U14013 ( .A(n439), .ZN(n20657) );
  INV_X1 U14014 ( .A(n439), .ZN(n20658) );
  INV_X1 U14015 ( .A(n18039), .ZN(n20659) );
  INV_X1 U14016 ( .A(n18039), .ZN(n20660) );
  INV_X1 U14017 ( .A(n438), .ZN(n20661) );
  INV_X1 U14018 ( .A(n438), .ZN(n20662) );
  INV_X1 U14019 ( .A(n437), .ZN(n20663) );
  INV_X1 U14020 ( .A(n437), .ZN(n20664) );
  INV_X1 U14021 ( .A(n436), .ZN(n20665) );
  INV_X1 U14022 ( .A(n436), .ZN(n20666) );
  INV_X1 U14023 ( .A(n18040), .ZN(n20667) );
  INV_X1 U14024 ( .A(n18040), .ZN(n20668) );
  INV_X1 U14025 ( .A(n435), .ZN(n20669) );
  INV_X1 U14026 ( .A(n435), .ZN(n20670) );
  INV_X1 U14027 ( .A(n434), .ZN(n20671) );
  INV_X1 U14028 ( .A(n434), .ZN(n20672) );
  INV_X1 U14029 ( .A(n433), .ZN(n20673) );
  INV_X1 U14030 ( .A(n433), .ZN(n20674) );
  INV_X1 U14031 ( .A(n18041), .ZN(n20675) );
  INV_X1 U14032 ( .A(n18041), .ZN(n20676) );
  INV_X1 U14033 ( .A(n432), .ZN(n20677) );
  INV_X1 U14034 ( .A(n432), .ZN(n20678) );
  INV_X1 U14035 ( .A(n431), .ZN(n20679) );
  INV_X1 U14036 ( .A(n431), .ZN(n20680) );
  INV_X1 U14037 ( .A(n430), .ZN(n20681) );
  INV_X1 U14038 ( .A(n430), .ZN(n20682) );
  INV_X1 U14039 ( .A(n18042), .ZN(n20683) );
  INV_X1 U14040 ( .A(n18042), .ZN(n20684) );
  INV_X1 U14041 ( .A(n429), .ZN(n20685) );
  INV_X1 U14042 ( .A(n429), .ZN(n20686) );
  INV_X1 U14043 ( .A(n18043), .ZN(n20687) );
  INV_X1 U14044 ( .A(n18043), .ZN(n20688) );
  INV_X1 U14045 ( .A(n18044), .ZN(n20689) );
  INV_X1 U14046 ( .A(n18044), .ZN(n20690) );
  INV_X1 U14047 ( .A(n18045), .ZN(n20691) );
  INV_X1 U14048 ( .A(n18045), .ZN(n20692) );
  INV_X1 U14049 ( .A(n18046), .ZN(n20693) );
  INV_X1 U14050 ( .A(n18046), .ZN(n20694) );
  INV_X1 U14051 ( .A(n27123), .ZN(n20695) );
  BUF_X1 U14052 ( .A(n24645), .Z(n27123) );
  BUF_X1 U14053 ( .A(n24645), .Z(n27124) );
  INV_X1 U14054 ( .A(n18047), .ZN(n20696) );
  INV_X1 U14055 ( .A(n18048), .ZN(n20697) );
  INV_X1 U14056 ( .A(n18049), .ZN(n20698) );
  INV_X1 U14057 ( .A(n18050), .ZN(n20699) );
  INV_X1 U14058 ( .A(n24874), .ZN(n20700) );
  INV_X1 U14059 ( .A(n20700), .ZN(n20701) );
  INV_X1 U14060 ( .A(n26806), .ZN(n20702) );
  INV_X1 U14061 ( .A(n20702), .ZN(n20703) );
  INV_X1 U14062 ( .A(n24879), .ZN(n20704) );
  INV_X1 U14063 ( .A(n20704), .ZN(n20705) );
  INV_X1 U14064 ( .A(n18051), .ZN(n20706) );
  INV_X1 U14065 ( .A(n18052), .ZN(n20707) );
  INV_X1 U14066 ( .A(n18053), .ZN(n20708) );
  INV_X1 U14067 ( .A(n18054), .ZN(n20709) );
  INV_X1 U14068 ( .A(n18055), .ZN(n20710) );
  INV_X1 U14069 ( .A(n18056), .ZN(n20711) );
  INV_X1 U14070 ( .A(n18057), .ZN(n20712) );
  INV_X1 U14071 ( .A(n18058), .ZN(n20713) );
  INV_X1 U14072 ( .A(n18985), .ZN(n20714) );
  INV_X1 U14073 ( .A(n20714), .ZN(n20715) );
  INV_X1 U14074 ( .A(n18986), .ZN(n20716) );
  INV_X1 U14075 ( .A(n20716), .ZN(n20717) );
  INV_X1 U14076 ( .A(n18059), .ZN(n20718) );
  INV_X1 U14077 ( .A(n18060), .ZN(n20719) );
  INV_X1 U14078 ( .A(n18061), .ZN(n20720) );
  INV_X1 U14079 ( .A(n18062), .ZN(n20721) );
  INV_X1 U14080 ( .A(n18063), .ZN(n20722) );
  INV_X1 U14081 ( .A(n18064), .ZN(n20723) );
  INV_X1 U14082 ( .A(n18064), .ZN(n20724) );
  INV_X1 U14083 ( .A(n18065), .ZN(n20725) );
  INV_X1 U14084 ( .A(n18065), .ZN(n20726) );
  INV_X1 U14085 ( .A(n18066), .ZN(n20727) );
  INV_X1 U14086 ( .A(n18066), .ZN(n20728) );
  INV_X1 U14087 ( .A(n18067), .ZN(n20729) );
  INV_X1 U14088 ( .A(n18067), .ZN(n20730) );
  INV_X1 U14089 ( .A(n18068), .ZN(n20731) );
  INV_X1 U14090 ( .A(n18069), .ZN(n20732) );
  INV_X1 U14091 ( .A(n18069), .ZN(n20733) );
  INV_X1 U14092 ( .A(n17089), .ZN(n20734) );
  INV_X1 U14093 ( .A(n20734), .ZN(n20735) );
  INV_X1 U14094 ( .A(n20734), .ZN(n20736) );
  INV_X1 U14095 ( .A(n17089), .ZN(n20737) );
  INV_X1 U14096 ( .A(n20737), .ZN(n20738) );
  INV_X1 U14097 ( .A(n20737), .ZN(n20739) );
  INV_X1 U14098 ( .A(n18070), .ZN(n20740) );
  INV_X1 U14099 ( .A(n18070), .ZN(n20741) );
  INV_X1 U14100 ( .A(n18071), .ZN(n20742) );
  INV_X1 U14101 ( .A(n18071), .ZN(n20743) );
  INV_X1 U14102 ( .A(n18072), .ZN(n20744) );
  INV_X1 U14103 ( .A(n18072), .ZN(n20745) );
  INV_X1 U14104 ( .A(n18073), .ZN(n20746) );
  INV_X1 U14105 ( .A(n18073), .ZN(n20747) );
  INV_X1 U14106 ( .A(n18074), .ZN(n20748) );
  INV_X1 U14107 ( .A(n18074), .ZN(n20749) );
  INV_X1 U14108 ( .A(n428), .ZN(n20750) );
  INV_X1 U14109 ( .A(n428), .ZN(n20751) );
  INV_X1 U14110 ( .A(n18075), .ZN(n20752) );
  INV_X1 U14111 ( .A(n18075), .ZN(n20753) );
  INV_X1 U14112 ( .A(n427), .ZN(n20754) );
  INV_X1 U14113 ( .A(n427), .ZN(n20755) );
  INV_X1 U14114 ( .A(n426), .ZN(n20756) );
  INV_X1 U14115 ( .A(n426), .ZN(n20757) );
  INV_X1 U14116 ( .A(n425), .ZN(n20758) );
  INV_X1 U14117 ( .A(n425), .ZN(n20759) );
  INV_X1 U14118 ( .A(n424), .ZN(n20760) );
  INV_X1 U14119 ( .A(n424), .ZN(n20761) );
  INV_X1 U14120 ( .A(n423), .ZN(n20762) );
  INV_X1 U14121 ( .A(n423), .ZN(n20763) );
  INV_X1 U14122 ( .A(n422), .ZN(n20764) );
  INV_X1 U14123 ( .A(n422), .ZN(n20765) );
  INV_X1 U14124 ( .A(n421), .ZN(n20766) );
  INV_X1 U14125 ( .A(n421), .ZN(n20767) );
  INV_X1 U14126 ( .A(n420), .ZN(n20768) );
  INV_X1 U14127 ( .A(n420), .ZN(n20769) );
  INV_X1 U14128 ( .A(n419), .ZN(n20770) );
  INV_X1 U14129 ( .A(n419), .ZN(n20771) );
  INV_X1 U14130 ( .A(n418), .ZN(n20772) );
  INV_X1 U14131 ( .A(n418), .ZN(n20773) );
  INV_X1 U14132 ( .A(n24984), .ZN(n20774) );
  INV_X1 U14133 ( .A(n20883), .ZN(n20775) );
  INV_X1 U14134 ( .A(n25060), .ZN(n20776) );
  INV_X1 U14135 ( .A(n20776), .ZN(n20777) );
  INV_X1 U14136 ( .A(n20776), .ZN(n20778) );
  INV_X1 U14137 ( .A(n27796), .ZN(n20779) );
  INV_X1 U14138 ( .A(n20779), .ZN(n20780) );
  INV_X1 U14139 ( .A(n20779), .ZN(n20781) );
  INV_X1 U14140 ( .A(n25083), .ZN(n20782) );
  INV_X1 U14141 ( .A(n20782), .ZN(n20783) );
  INV_X1 U14142 ( .A(n20782), .ZN(n20784) );
  INV_X1 U14143 ( .A(n18076), .ZN(n20785) );
  INV_X1 U14144 ( .A(n18076), .ZN(n20786) );
  INV_X1 U14145 ( .A(n18077), .ZN(n20787) );
  INV_X1 U14146 ( .A(n18077), .ZN(n20788) );
  INV_X1 U14147 ( .A(n18078), .ZN(n20789) );
  INV_X1 U14148 ( .A(n18078), .ZN(n20790) );
  CLKBUF_X1 U14149 ( .A(n24993), .Z(n20791) );
  INV_X1 U14150 ( .A(n18079), .ZN(n20792) );
  INV_X1 U14151 ( .A(n18079), .ZN(n20793) );
  INV_X1 U14152 ( .A(n18080), .ZN(n20794) );
  INV_X1 U14153 ( .A(n18080), .ZN(n20795) );
  INV_X1 U14154 ( .A(n18081), .ZN(n20796) );
  INV_X1 U14155 ( .A(n18081), .ZN(n20797) );
  CLKBUF_X1 U14156 ( .A(n25001), .Z(n20798) );
  INV_X1 U14157 ( .A(n18082), .ZN(n20799) );
  INV_X1 U14158 ( .A(n18082), .ZN(n20800) );
  INV_X1 U14159 ( .A(n18083), .ZN(n20801) );
  INV_X1 U14160 ( .A(n18083), .ZN(n20802) );
  INV_X1 U14161 ( .A(n18084), .ZN(n20803) );
  INV_X1 U14162 ( .A(n18084), .ZN(n20804) );
  INV_X1 U14163 ( .A(n18085), .ZN(n20805) );
  INV_X1 U14164 ( .A(n18085), .ZN(n20806) );
  INV_X1 U14165 ( .A(n18086), .ZN(n20807) );
  INV_X1 U14166 ( .A(n18086), .ZN(n20808) );
  INV_X1 U14167 ( .A(n18087), .ZN(n20809) );
  INV_X1 U14168 ( .A(n18088), .ZN(n20810) );
  INV_X1 U14169 ( .A(n18088), .ZN(n20811) );
  INV_X1 U14170 ( .A(n417), .ZN(n20812) );
  INV_X1 U14171 ( .A(n417), .ZN(n20813) );
  INV_X1 U14172 ( .A(n18089), .ZN(n20814) );
  INV_X1 U14173 ( .A(n18089), .ZN(n20815) );
  INV_X1 U14174 ( .A(n416), .ZN(n20816) );
  INV_X1 U14175 ( .A(n416), .ZN(n20817) );
  INV_X1 U14176 ( .A(n415), .ZN(n20818) );
  INV_X1 U14177 ( .A(n415), .ZN(n20819) );
  INV_X1 U14178 ( .A(n414), .ZN(n20820) );
  INV_X1 U14179 ( .A(n414), .ZN(n20821) );
  INV_X1 U14180 ( .A(n413), .ZN(n20822) );
  INV_X1 U14181 ( .A(n413), .ZN(n20823) );
  INV_X1 U14182 ( .A(n412), .ZN(n20824) );
  INV_X1 U14183 ( .A(n412), .ZN(n20825) );
  INV_X1 U14184 ( .A(n411), .ZN(n20826) );
  INV_X1 U14185 ( .A(n411), .ZN(n20827) );
  INV_X1 U14186 ( .A(n410), .ZN(n20828) );
  INV_X1 U14187 ( .A(n410), .ZN(n20829) );
  INV_X1 U14188 ( .A(n409), .ZN(n20830) );
  INV_X1 U14189 ( .A(n409), .ZN(n20831) );
  INV_X1 U14190 ( .A(n408), .ZN(n20832) );
  INV_X1 U14191 ( .A(n408), .ZN(n20833) );
  INV_X1 U14192 ( .A(n407), .ZN(n20834) );
  INV_X1 U14193 ( .A(n407), .ZN(n20835) );
  INV_X1 U14194 ( .A(n406), .ZN(n20836) );
  INV_X1 U14195 ( .A(n406), .ZN(n20837) );
  INV_X1 U14196 ( .A(n405), .ZN(n20838) );
  INV_X1 U14197 ( .A(n405), .ZN(n20839) );
  INV_X1 U14198 ( .A(n404), .ZN(n20840) );
  INV_X1 U14199 ( .A(n404), .ZN(n20841) );
  INV_X1 U14200 ( .A(n403), .ZN(n20842) );
  INV_X1 U14201 ( .A(n403), .ZN(n20843) );
  INV_X1 U14202 ( .A(n402), .ZN(n20844) );
  INV_X1 U14203 ( .A(n402), .ZN(n20845) );
  INV_X1 U14204 ( .A(n401), .ZN(n20846) );
  INV_X1 U14205 ( .A(n401), .ZN(n20847) );
  INV_X1 U14206 ( .A(n400), .ZN(n20848) );
  INV_X1 U14207 ( .A(n400), .ZN(n20849) );
  INV_X1 U14208 ( .A(n399), .ZN(n20850) );
  INV_X1 U14209 ( .A(n399), .ZN(n20851) );
  INV_X1 U14210 ( .A(n398), .ZN(n20852) );
  INV_X1 U14211 ( .A(n398), .ZN(n20853) );
  INV_X1 U14212 ( .A(n397), .ZN(n20854) );
  INV_X1 U14213 ( .A(n397), .ZN(n20855) );
  INV_X1 U14214 ( .A(n25060), .ZN(n20856) );
  INV_X1 U14215 ( .A(n20856), .ZN(n20857) );
  INV_X1 U14216 ( .A(n20856), .ZN(n20858) );
  INV_X1 U14217 ( .A(n396), .ZN(n20859) );
  INV_X1 U14218 ( .A(n396), .ZN(n20860) );
  INV_X1 U14219 ( .A(n18090), .ZN(n20861) );
  INV_X1 U14220 ( .A(n18090), .ZN(n20862) );
  INV_X1 U14221 ( .A(n26584), .ZN(n20863) );
  INV_X1 U14222 ( .A(n20863), .ZN(n20864) );
  INV_X1 U14223 ( .A(n20863), .ZN(n20865) );
  INV_X1 U14224 ( .A(n18091), .ZN(n20866) );
  INV_X1 U14225 ( .A(n18091), .ZN(n20867) );
  INV_X1 U14226 ( .A(n18092), .ZN(n20868) );
  INV_X1 U14227 ( .A(n18092), .ZN(n20869) );
  INV_X1 U14228 ( .A(n18093), .ZN(n20870) );
  INV_X1 U14229 ( .A(n18093), .ZN(n20871) );
  INV_X1 U14230 ( .A(n18094), .ZN(n20872) );
  INV_X1 U14231 ( .A(n18094), .ZN(n20873) );
  INV_X1 U14232 ( .A(n18095), .ZN(n20874) );
  INV_X1 U14233 ( .A(n18095), .ZN(n20875) );
  INV_X1 U14234 ( .A(n18096), .ZN(n20876) );
  INV_X1 U14235 ( .A(n18096), .ZN(n20877) );
  INV_X1 U14236 ( .A(n25079), .ZN(n20878) );
  INV_X1 U14237 ( .A(n18097), .ZN(n20879) );
  INV_X1 U14238 ( .A(n18097), .ZN(n20880) );
  INV_X1 U14239 ( .A(n259701), .ZN(n20881) );
  INV_X1 U14240 ( .A(n20881), .ZN(n20882) );
  INV_X1 U14241 ( .A(n20881), .ZN(n20883) );
  INV_X1 U14242 ( .A(n27293), .ZN(n20884) );
  INV_X1 U14243 ( .A(n20884), .ZN(n20885) );
  INV_X1 U14244 ( .A(n20884), .ZN(n20886) );
  INV_X1 U14245 ( .A(n19016), .ZN(n20887) );
  INV_X1 U14246 ( .A(n20887), .ZN(n20888) );
  INV_X1 U14247 ( .A(n20887), .ZN(n20889) );
  INV_X1 U14248 ( .A(n54240), .ZN(n20890) );
  INV_X1 U14249 ( .A(n20890), .ZN(n20891) );
  INV_X1 U14250 ( .A(n20890), .ZN(n20892) );
  INV_X1 U14251 ( .A(n25085), .ZN(n20893) );
  INV_X1 U14252 ( .A(n20893), .ZN(n20894) );
  INV_X1 U14253 ( .A(n18098), .ZN(n20895) );
  INV_X1 U14254 ( .A(n18098), .ZN(n20896) );
  INV_X1 U14255 ( .A(n25088), .ZN(n20897) );
  INV_X1 U14256 ( .A(n20897), .ZN(n20898) );
  INV_X1 U14257 ( .A(n43460), .ZN(n20899) );
  INV_X1 U14258 ( .A(n20899), .ZN(n20900) );
  INV_X1 U14259 ( .A(n20899), .ZN(n20901) );
  INV_X1 U14260 ( .A(n18099), .ZN(n20902) );
  INV_X1 U14261 ( .A(n18099), .ZN(n20903) );
  INV_X1 U14262 ( .A(n3103), .ZN(n20904) );
  INV_X1 U14263 ( .A(n20904), .ZN(n20905) );
  INV_X1 U14264 ( .A(n20904), .ZN(n20906) );
  INV_X1 U14265 ( .A(n18100), .ZN(n20907) );
  INV_X1 U14266 ( .A(n18100), .ZN(n20908) );
  INV_X1 U14267 ( .A(n27230), .ZN(n20909) );
  INV_X1 U14268 ( .A(n25092), .ZN(n20910) );
  INV_X1 U14269 ( .A(n20910), .ZN(n20911) );
  INV_X1 U14270 ( .A(n27175), .ZN(n20912) );
  INV_X1 U14271 ( .A(n27231), .ZN(n20913) );
  INV_X1 U14272 ( .A(n19024), .ZN(n20914) );
  INV_X1 U14273 ( .A(n20914), .ZN(n20915) );
  INV_X1 U14274 ( .A(n27176), .ZN(n20916) );
  INV_X1 U14275 ( .A(n18101), .ZN(n20917) );
  INV_X1 U14276 ( .A(n19028), .ZN(n20918) );
  INV_X1 U14277 ( .A(n20918), .ZN(n20919) );
  INV_X1 U14278 ( .A(n18102), .ZN(n20920) );
  INV_X1 U14279 ( .A(n18103), .ZN(n20921) );
  INV_X1 U14280 ( .A(n18103), .ZN(n20922) );
  INV_X1 U14281 ( .A(n21399), .ZN(n20923) );
  INV_X1 U14282 ( .A(n20923), .ZN(n20924) );
  INV_X1 U14283 ( .A(n18104), .ZN(n20925) );
  INV_X1 U14284 ( .A(n18105), .ZN(n20926) );
  INV_X1 U14285 ( .A(n18105), .ZN(n20927) );
  INV_X1 U14286 ( .A(n18106), .ZN(n20928) );
  INV_X1 U14287 ( .A(n18107), .ZN(n20929) );
  INV_X1 U14288 ( .A(n18108), .ZN(n20930) );
  INV_X1 U14289 ( .A(n18109), .ZN(n20931) );
  INV_X1 U14290 ( .A(n18110), .ZN(n20932) );
  INV_X1 U14291 ( .A(n18111), .ZN(n20933) );
  INV_X1 U14292 ( .A(n18112), .ZN(n20934) );
  INV_X1 U14293 ( .A(n25133), .ZN(n20935) );
  INV_X1 U14294 ( .A(n20935), .ZN(n20936) );
  INV_X1 U14295 ( .A(n20935), .ZN(n20937) );
  INV_X1 U14296 ( .A(n25133), .ZN(n20938) );
  INV_X1 U14297 ( .A(n20938), .ZN(n20939) );
  INV_X1 U14298 ( .A(n20938), .ZN(n20940) );
  INV_X1 U14299 ( .A(n18113), .ZN(n20941) );
  INV_X1 U14300 ( .A(n25142), .ZN(n20942) );
  INV_X1 U14301 ( .A(n20942), .ZN(n20943) );
  INV_X1 U14302 ( .A(n18114), .ZN(n20944) );
  INV_X1 U14303 ( .A(n25151), .ZN(n20945) );
  INV_X1 U14304 ( .A(n20945), .ZN(n20946) );
  INV_X1 U14305 ( .A(n20945), .ZN(n20947) );
  INV_X1 U14306 ( .A(n25151), .ZN(n20948) );
  INV_X1 U14307 ( .A(n20948), .ZN(n20949) );
  INV_X1 U14308 ( .A(n20948), .ZN(n20950) );
  INV_X1 U14309 ( .A(n17136), .ZN(n20951) );
  INV_X1 U14310 ( .A(n25160), .ZN(n20952) );
  INV_X1 U14311 ( .A(n20952), .ZN(n20953) );
  INV_X1 U14312 ( .A(n18116), .ZN(n20954) );
  INV_X1 U14313 ( .A(n18117), .ZN(n20955) );
  INV_X1 U14314 ( .A(n18118), .ZN(n20956) );
  INV_X1 U14315 ( .A(n18119), .ZN(n20957) );
  INV_X1 U14316 ( .A(n18120), .ZN(n20958) );
  INV_X1 U14317 ( .A(n18121), .ZN(n20959) );
  INV_X1 U14318 ( .A(n18122), .ZN(n20960) );
  INV_X1 U14319 ( .A(n18122), .ZN(n20961) );
  INV_X1 U14320 ( .A(n18123), .ZN(n20962) );
  INV_X1 U14321 ( .A(n20968), .ZN(n20963) );
  INV_X1 U14322 ( .A(n20963), .ZN(n20964) );
  INV_X1 U14323 ( .A(n20970), .ZN(n20965) );
  INV_X1 U14324 ( .A(n20965), .ZN(n20966) );
  INV_X1 U14325 ( .A(n27188), .ZN(n20967) );
  INV_X1 U14326 ( .A(n25075), .ZN(n20968) );
  INV_X1 U14327 ( .A(n27244), .ZN(n20969) );
  INV_X1 U14328 ( .A(n25081), .ZN(n20970) );
  INV_X1 U14329 ( .A(n23089), .ZN(n20971) );
  INV_X1 U14330 ( .A(n20971), .ZN(n20972) );
  INV_X1 U14331 ( .A(n20971), .ZN(n20973) );
  INV_X1 U14332 ( .A(n18124), .ZN(n20974) );
  INV_X1 U14333 ( .A(n18124), .ZN(n20975) );
  INV_X1 U14334 ( .A(n23090), .ZN(n20976) );
  INV_X1 U14335 ( .A(n20976), .ZN(n20977) );
  INV_X1 U14336 ( .A(n20976), .ZN(n20978) );
  INV_X1 U14337 ( .A(n25207), .ZN(n20979) );
  INV_X1 U14338 ( .A(n20979), .ZN(n20980) );
  INV_X1 U14339 ( .A(n20979), .ZN(n20981) );
  INV_X1 U14340 ( .A(n18125), .ZN(n20982) );
  INV_X1 U14341 ( .A(n18125), .ZN(n20983) );
  INV_X1 U14342 ( .A(n18126), .ZN(n20984) );
  INV_X1 U14343 ( .A(n18126), .ZN(n20985) );
  INV_X1 U14344 ( .A(n18127), .ZN(n20986) );
  INV_X1 U14345 ( .A(n25219), .ZN(n20987) );
  INV_X1 U14346 ( .A(n20987), .ZN(n20988) );
  INV_X1 U14347 ( .A(n20987), .ZN(n20989) );
  INV_X1 U14348 ( .A(n18128), .ZN(n20990) );
  INV_X1 U14349 ( .A(n18129), .ZN(n20991) );
  INV_X1 U14350 ( .A(n18130), .ZN(n20992) );
  INV_X1 U14351 ( .A(n18131), .ZN(n20993) );
  INV_X1 U14352 ( .A(n18132), .ZN(n20994) );
  INV_X1 U14353 ( .A(n18133), .ZN(n20995) );
  INV_X1 U14354 ( .A(n18134), .ZN(n20996) );
  INV_X1 U14355 ( .A(n18135), .ZN(n20997) );
  INV_X1 U14356 ( .A(n24654), .ZN(n20998) );
  INV_X1 U14357 ( .A(n20998), .ZN(n20999) );
  INV_X1 U14358 ( .A(n18136), .ZN(n21000) );
  INV_X1 U14359 ( .A(n18136), .ZN(n21001) );
  INV_X1 U14360 ( .A(n18137), .ZN(n21002) );
  INV_X1 U14361 ( .A(n18138), .ZN(n21003) );
  INV_X1 U14362 ( .A(n18138), .ZN(n21004) );
  INV_X1 U14363 ( .A(n27803), .ZN(n21005) );
  INV_X1 U14364 ( .A(n21005), .ZN(n21006) );
  INV_X1 U14365 ( .A(n18139), .ZN(n21007) );
  INV_X1 U14366 ( .A(n18140), .ZN(n21008) );
  INV_X1 U14367 ( .A(n25252), .ZN(n21009) );
  INV_X1 U14368 ( .A(n21009), .ZN(n21010) );
  INV_X1 U14369 ( .A(n21009), .ZN(n21011) );
  INV_X1 U14370 ( .A(n18141), .ZN(n21012) );
  INV_X1 U14371 ( .A(n25285), .ZN(n21013) );
  INV_X1 U14372 ( .A(n21013), .ZN(n21014) );
  INV_X1 U14373 ( .A(n21013), .ZN(n21015) );
  INV_X1 U14374 ( .A(n18142), .ZN(n21016) );
  INV_X1 U14375 ( .A(n18143), .ZN(n21017) );
  INV_X1 U14376 ( .A(n18144), .ZN(n21018) );
  INV_X1 U14377 ( .A(n18145), .ZN(n21019) );
  INV_X1 U14378 ( .A(n18146), .ZN(n21020) );
  INV_X1 U14379 ( .A(n18147), .ZN(n21021) );
  INV_X1 U14380 ( .A(n27792), .ZN(n21022) );
  INV_X1 U14381 ( .A(n21022), .ZN(n21023) );
  INV_X1 U14382 ( .A(n21022), .ZN(n21024) );
  INV_X1 U14383 ( .A(n18148), .ZN(n21025) );
  INV_X1 U14384 ( .A(n18150), .ZN(n21026) );
  INV_X1 U14385 ( .A(n18151), .ZN(n21027) );
  INV_X1 U14386 ( .A(n18152), .ZN(n21028) );
  INV_X1 U14387 ( .A(n26712), .ZN(n21029) );
  INV_X1 U14388 ( .A(n21029), .ZN(n21030) );
  INV_X1 U14389 ( .A(n26708), .ZN(n21031) );
  INV_X1 U14390 ( .A(n21031), .ZN(n21032) );
  INV_X1 U14391 ( .A(n18153), .ZN(n21033) );
  INV_X1 U14392 ( .A(n26702), .ZN(n21034) );
  INV_X1 U14393 ( .A(n21034), .ZN(n21035) );
  INV_X1 U14394 ( .A(n26705), .ZN(n21036) );
  INV_X1 U14395 ( .A(n21036), .ZN(n21037) );
  INV_X1 U14396 ( .A(n25332), .ZN(n21038) );
  INV_X1 U14397 ( .A(n21038), .ZN(n21039) );
  INV_X1 U14398 ( .A(n18154), .ZN(n21040) );
  INV_X1 U14399 ( .A(n25337), .ZN(n21041) );
  INV_X1 U14400 ( .A(n21041), .ZN(n21042) );
  INV_X1 U14401 ( .A(n25340), .ZN(n21043) );
  INV_X1 U14402 ( .A(n21043), .ZN(n21044) );
  INV_X1 U14403 ( .A(n25343), .ZN(n21045) );
  INV_X1 U14404 ( .A(n21045), .ZN(n21046) );
  INV_X1 U14405 ( .A(n25092), .ZN(n21047) );
  INV_X1 U14406 ( .A(n21047), .ZN(n21048) );
  INV_X1 U14407 ( .A(n18155), .ZN(n21049) );
  INV_X1 U14408 ( .A(n18156), .ZN(n21050) );
  INV_X1 U14409 ( .A(n18157), .ZN(n21051) );
  INV_X1 U14410 ( .A(n18158), .ZN(n21052) );
  INV_X1 U14411 ( .A(n18159), .ZN(n21053) );
  INV_X1 U14412 ( .A(n18160), .ZN(n21054) );
  INV_X1 U14413 ( .A(n18161), .ZN(n21055) );
  INV_X1 U14414 ( .A(n22692), .ZN(n21056) );
  INV_X1 U14415 ( .A(n22692), .ZN(n21057) );
  INV_X1 U14416 ( .A(n18163), .ZN(n21058) );
  INV_X1 U14417 ( .A(n18163), .ZN(n21059) );
  INV_X1 U14418 ( .A(n18164), .ZN(n21060) );
  INV_X1 U14419 ( .A(n18165), .ZN(n21061) );
  INV_X1 U14420 ( .A(n18166), .ZN(n21062) );
  INV_X1 U14421 ( .A(n18166), .ZN(n21063) );
  INV_X1 U14422 ( .A(n27260), .ZN(n21064) );
  INV_X1 U14423 ( .A(n18167), .ZN(n21065) );
  INV_X1 U14424 ( .A(n18167), .ZN(n21066) );
  INV_X1 U14425 ( .A(n18168), .ZN(n21067) );
  INV_X1 U14426 ( .A(n18169), .ZN(n21068) );
  INV_X1 U14427 ( .A(n18170), .ZN(n21069) );
  INV_X1 U14428 ( .A(n18171), .ZN(n21070) );
  INV_X1 U14429 ( .A(n3104), .ZN(n21071) );
  INV_X1 U14430 ( .A(n3072), .ZN(n21072) );
  INV_X1 U14431 ( .A(n3154), .ZN(n21073) );
  INV_X1 U14432 ( .A(n31290), .ZN(n21074) );
  INV_X1 U14433 ( .A(n32040), .ZN(n21075) );
  INV_X1 U14434 ( .A(n3179), .ZN(n21076) );
  INV_X1 U14435 ( .A(n32540), .ZN(n21077) );
  INV_X1 U14436 ( .A(n3229), .ZN(n21078) );
  INV_X1 U14437 ( .A(n33030), .ZN(n21079) );
  INV_X1 U14438 ( .A(n3278), .ZN(n21080) );
  INV_X1 U14439 ( .A(n3347), .ZN(n21081) );
  INV_X1 U14440 ( .A(n3325), .ZN(n21082) );
  INV_X1 U14441 ( .A(n3391), .ZN(n21083) );
  INV_X1 U14442 ( .A(n33690), .ZN(n21084) );
  INV_X1 U14443 ( .A(n3436), .ZN(n21085) );
  INV_X1 U14444 ( .A(n3413), .ZN(n21086) );
  INV_X1 U14445 ( .A(n3485), .ZN(n21087) );
  INV_X1 U14446 ( .A(n34600), .ZN(n21088) );
  INV_X1 U14447 ( .A(n3529), .ZN(n21089) );
  INV_X1 U14448 ( .A(n35070), .ZN(n21090) );
  INV_X1 U14449 ( .A(n3573), .ZN(n21091) );
  INV_X1 U14450 ( .A(n35510), .ZN(n21092) );
  INV_X1 U14451 ( .A(n3618), .ZN(n21093) );
  INV_X1 U14452 ( .A(n35950), .ZN(n21094) );
  INV_X1 U14453 ( .A(n3666), .ZN(n21095) );
  INV_X1 U14454 ( .A(n3642), .ZN(n21096) );
  INV_X1 U14455 ( .A(n37100), .ZN(n21097) );
  INV_X1 U14456 ( .A(n3688), .ZN(n21098) );
  INV_X1 U14457 ( .A(n3754), .ZN(n21099) );
  INV_X1 U14458 ( .A(n3732), .ZN(n21100) );
  INV_X1 U14459 ( .A(n37990), .ZN(n21101) );
  INV_X1 U14460 ( .A(n3776), .ZN(n21102) );
  INV_X1 U14461 ( .A(n38480), .ZN(n21103) );
  INV_X1 U14462 ( .A(n3823), .ZN(n21104) );
  INV_X1 U14463 ( .A(n3892), .ZN(n21105) );
  INV_X1 U14464 ( .A(n3870), .ZN(n21106) );
  INV_X1 U14465 ( .A(n39360), .ZN(n21107) );
  INV_X1 U14466 ( .A(n3914), .ZN(n21108) );
  INV_X1 U14467 ( .A(n3981), .ZN(n21109) );
  INV_X1 U14468 ( .A(n3958), .ZN(n21110) );
  INV_X1 U14469 ( .A(n4031), .ZN(n21111) );
  INV_X1 U14470 ( .A(n4005), .ZN(n21112) );
  INV_X1 U14471 ( .A(n4075), .ZN(n21113) );
  INV_X1 U14472 ( .A(n4119), .ZN(n21114) );
  INV_X1 U14473 ( .A(n40970), .ZN(n21115) );
  INV_X1 U14474 ( .A(n4164), .ZN(n21116) );
  INV_X1 U14475 ( .A(n41410), .ZN(n21117) );
  INV_X1 U14476 ( .A(n42140), .ZN(n21118) );
  INV_X1 U14477 ( .A(n41880), .ZN(n21119) );
  INV_X1 U14478 ( .A(n4258), .ZN(n21120) );
  INV_X1 U14479 ( .A(n4236), .ZN(n21121) );
  INV_X1 U14480 ( .A(n43020), .ZN(n21122) );
  INV_X1 U14481 ( .A(n4280), .ZN(n21123) );
  INV_X1 U14482 ( .A(n43470), .ZN(n21124) );
  INV_X1 U14483 ( .A(n4324), .ZN(n21125) );
  INV_X1 U14484 ( .A(n4396), .ZN(n21126) );
  INV_X1 U14485 ( .A(n4371), .ZN(n21127) );
  INV_X1 U14486 ( .A(n44450), .ZN(n21128) );
  INV_X1 U14487 ( .A(n4421), .ZN(n21129) );
  INV_X1 U14488 ( .A(n4494), .ZN(n21130) );
  INV_X1 U14489 ( .A(n44700), .ZN(n21131) );
  INV_X1 U14490 ( .A(n4543), .ZN(n21132) );
  INV_X1 U14491 ( .A(n45180), .ZN(n21133) );
  INV_X1 U14492 ( .A(n4419), .ZN(n21134) );
  INV_X1 U14493 ( .A(n25510), .ZN(n21135) );
  INV_X1 U14494 ( .A(n21135), .ZN(n21136) );
  INV_X1 U14495 ( .A(n18172), .ZN(n21137) );
  INV_X1 U14496 ( .A(n25515), .ZN(n21138) );
  INV_X1 U14497 ( .A(n21138), .ZN(n21139) );
  INV_X1 U14498 ( .A(n18173), .ZN(n21140) );
  INV_X1 U14499 ( .A(n18173), .ZN(n21141) );
  INV_X1 U14500 ( .A(n4029), .ZN(n21142) );
  INV_X1 U14501 ( .A(n21142), .ZN(n21143) );
  INV_X1 U14502 ( .A(n25519), .ZN(n21144) );
  INV_X1 U14503 ( .A(n21144), .ZN(n21145) );
  INV_X1 U14504 ( .A(n21144), .ZN(n21146) );
  INV_X1 U14505 ( .A(n18174), .ZN(n21147) );
  INV_X1 U14506 ( .A(n18174), .ZN(n21148) );
  INV_X1 U14507 ( .A(n18175), .ZN(n21149) );
  INV_X1 U14508 ( .A(n18176), .ZN(n21150) );
  INV_X1 U14509 ( .A(n18176), .ZN(n21151) );
  INV_X1 U14510 ( .A(n18177), .ZN(n21152) );
  INV_X1 U14511 ( .A(n18178), .ZN(n21153) );
  INV_X1 U14512 ( .A(n18178), .ZN(n21154) );
  INV_X1 U14513 ( .A(n18179), .ZN(n21155) );
  INV_X1 U14514 ( .A(n18180), .ZN(n21156) );
  INV_X1 U14515 ( .A(n18180), .ZN(n21157) );
  INV_X1 U14516 ( .A(n18181), .ZN(n21158) );
  INV_X1 U14517 ( .A(n18182), .ZN(n21159) );
  INV_X1 U14518 ( .A(n18182), .ZN(n21160) );
  INV_X1 U14519 ( .A(n25528), .ZN(n21161) );
  INV_X1 U14520 ( .A(n21161), .ZN(n21162) );
  INV_X1 U14521 ( .A(n21161), .ZN(n21163) );
  INV_X1 U14522 ( .A(n25340), .ZN(n21164) );
  INV_X1 U14523 ( .A(n21162), .ZN(n21165) );
  INV_X1 U14524 ( .A(n27158), .ZN(n21166) );
  INV_X1 U14525 ( .A(n18183), .ZN(n21167) );
  INV_X1 U14526 ( .A(n18183), .ZN(n21168) );
  INV_X1 U14527 ( .A(n18184), .ZN(n21169) );
  INV_X1 U14528 ( .A(n18184), .ZN(n21170) );
  INV_X1 U14529 ( .A(n18185), .ZN(n21171) );
  INV_X1 U14530 ( .A(n18185), .ZN(n21172) );
  CLKBUF_X1 U14531 ( .A(n17082), .Z(n21173) );
  INV_X1 U14532 ( .A(n25535), .ZN(n21174) );
  INV_X1 U14533 ( .A(n21174), .ZN(n21175) );
  INV_X1 U14534 ( .A(n21174), .ZN(n21176) );
  INV_X1 U14535 ( .A(n18186), .ZN(n21177) );
  INV_X1 U14536 ( .A(n18187), .ZN(n21178) );
  INV_X1 U14537 ( .A(n18187), .ZN(n21179) );
  CLKBUF_X1 U14538 ( .A(n25634), .Z(n21180) );
  INV_X1 U14539 ( .A(n25538), .ZN(n21181) );
  INV_X1 U14540 ( .A(n21181), .ZN(n21182) );
  INV_X1 U14541 ( .A(n21181), .ZN(n21183) );
  INV_X1 U14542 ( .A(n20491), .ZN(n21184) );
  INV_X1 U14543 ( .A(n18188), .ZN(n21185) );
  INV_X1 U14544 ( .A(n18188), .ZN(n21186) );
  INV_X1 U14545 ( .A(n25540), .ZN(n21187) );
  INV_X1 U14546 ( .A(n21187), .ZN(n21188) );
  INV_X1 U14547 ( .A(n25540), .ZN(n21189) );
  INV_X1 U14548 ( .A(n21188), .ZN(n21190) );
  INV_X1 U14549 ( .A(n18189), .ZN(n21191) );
  INV_X1 U14550 ( .A(n18190), .ZN(n21192) );
  INV_X1 U14551 ( .A(n18190), .ZN(n21193) );
  INV_X1 U14552 ( .A(n18191), .ZN(n21194) );
  INV_X1 U14553 ( .A(n18192), .ZN(n21195) );
  INV_X1 U14554 ( .A(n18192), .ZN(n21196) );
  INV_X1 U14555 ( .A(n18193), .ZN(n21197) );
  INV_X1 U14556 ( .A(n18194), .ZN(n21198) );
  INV_X1 U14557 ( .A(n18194), .ZN(n21199) );
  INV_X1 U14558 ( .A(n18195), .ZN(n21200) );
  INV_X1 U14559 ( .A(n18196), .ZN(n21201) );
  INV_X1 U14560 ( .A(n18196), .ZN(n21202) );
  INV_X1 U14561 ( .A(n18197), .ZN(n21203) );
  INV_X1 U14562 ( .A(n18198), .ZN(n21204) );
  INV_X1 U14563 ( .A(n18198), .ZN(n21205) );
  INV_X1 U14564 ( .A(n18199), .ZN(n21206) );
  INV_X1 U14565 ( .A(n18200), .ZN(n21207) );
  INV_X1 U14566 ( .A(n18200), .ZN(n21208) );
  INV_X1 U14567 ( .A(n24630), .ZN(n21209) );
  INV_X1 U14568 ( .A(n21209), .ZN(n21210) );
  INV_X1 U14569 ( .A(n18201), .ZN(n21211) );
  INV_X1 U14570 ( .A(n18201), .ZN(n21212) );
  INV_X1 U14571 ( .A(n24615), .ZN(n21213) );
  INV_X1 U14572 ( .A(n21213), .ZN(n21214) );
  INV_X1 U14573 ( .A(n18202), .ZN(n21215) );
  INV_X1 U14574 ( .A(n18202), .ZN(n21216) );
  INV_X1 U14575 ( .A(n18203), .ZN(n21217) );
  INV_X1 U14576 ( .A(n18204), .ZN(n21218) );
  INV_X1 U14577 ( .A(n18204), .ZN(n21219) );
  INV_X1 U14578 ( .A(n18205), .ZN(n21220) );
  INV_X1 U14579 ( .A(n18206), .ZN(n21221) );
  INV_X1 U14580 ( .A(n18206), .ZN(n21222) );
  INV_X1 U14581 ( .A(n18207), .ZN(n21223) );
  INV_X1 U14582 ( .A(n18208), .ZN(n21224) );
  INV_X1 U14583 ( .A(n18208), .ZN(n21225) );
  INV_X1 U14584 ( .A(n20483), .ZN(n21226) );
  INV_X1 U14585 ( .A(n18209), .ZN(n21227) );
  INV_X1 U14586 ( .A(n18209), .ZN(n21228) );
  INV_X1 U14587 ( .A(n18210), .ZN(n21229) );
  INV_X1 U14588 ( .A(n21229), .ZN(n21230) );
  INV_X1 U14589 ( .A(n4986), .ZN(n21231) );
  INV_X1 U14590 ( .A(n18211), .ZN(n21232) );
  INV_X1 U14591 ( .A(n18211), .ZN(n21233) );
  INV_X1 U14592 ( .A(n25569), .ZN(n21234) );
  INV_X1 U14593 ( .A(n21234), .ZN(n21235) );
  INV_X1 U14594 ( .A(n25569), .ZN(n21236) );
  INV_X1 U14595 ( .A(n21235), .ZN(n21237) );
  INV_X1 U14596 ( .A(n20486), .ZN(n21238) );
  INV_X1 U14597 ( .A(n18212), .ZN(n21239) );
  INV_X1 U14598 ( .A(n18212), .ZN(n21240) );
  INV_X1 U14599 ( .A(n25572), .ZN(n21241) );
  INV_X1 U14600 ( .A(n21241), .ZN(n21242) );
  INV_X1 U14601 ( .A(n25572), .ZN(n21243) );
  INV_X1 U14602 ( .A(n21242), .ZN(n21244) );
  INV_X1 U14603 ( .A(n18213), .ZN(n21245) );
  INV_X1 U14604 ( .A(n18214), .ZN(n21246) );
  INV_X1 U14605 ( .A(n18214), .ZN(n21247) );
  INV_X1 U14606 ( .A(n18215), .ZN(n21248) );
  INV_X1 U14607 ( .A(n21248), .ZN(n21249) );
  INV_X1 U14608 ( .A(n18216), .ZN(n21250) );
  INV_X1 U14609 ( .A(n18216), .ZN(n21251) );
  INV_X1 U14610 ( .A(n18217), .ZN(n21252) );
  INV_X1 U14611 ( .A(n18218), .ZN(n21253) );
  INV_X1 U14612 ( .A(n18218), .ZN(n21254) );
  INV_X1 U14613 ( .A(n18219), .ZN(n21255) );
  INV_X1 U14614 ( .A(n18219), .ZN(n21256) );
  INV_X1 U14615 ( .A(n18220), .ZN(n21257) );
  INV_X1 U14616 ( .A(n18221), .ZN(n21258) );
  INV_X1 U14617 ( .A(n18221), .ZN(n21259) );
  INV_X1 U14618 ( .A(n18222), .ZN(n21260) );
  INV_X1 U14619 ( .A(n18223), .ZN(n21261) );
  INV_X1 U14620 ( .A(n18223), .ZN(n21262) );
  INV_X1 U14621 ( .A(n20479), .ZN(n21263) );
  INV_X1 U14622 ( .A(n18224), .ZN(n21264) );
  INV_X1 U14623 ( .A(n18224), .ZN(n21265) );
  INV_X1 U14624 ( .A(n18225), .ZN(n21266) );
  INV_X1 U14625 ( .A(n21266), .ZN(n21267) );
  INV_X1 U14626 ( .A(n18226), .ZN(n21268) );
  INV_X1 U14627 ( .A(n18226), .ZN(n21269) );
  INV_X1 U14628 ( .A(n18227), .ZN(n21270) );
  INV_X1 U14629 ( .A(n18227), .ZN(n21271) );
  INV_X1 U14630 ( .A(n18228), .ZN(n21272) );
  INV_X1 U14631 ( .A(n18229), .ZN(n21273) );
  INV_X1 U14632 ( .A(n18229), .ZN(n21274) );
  INV_X1 U14633 ( .A(n18230), .ZN(n21275) );
  INV_X1 U14634 ( .A(n18231), .ZN(n21276) );
  INV_X1 U14635 ( .A(n18231), .ZN(n21277) );
  INV_X1 U14636 ( .A(n18232), .ZN(n21278) );
  INV_X1 U14637 ( .A(n18233), .ZN(n21279) );
  INV_X1 U14638 ( .A(n18233), .ZN(n21280) );
  CLKBUF_X1 U14639 ( .A(n25609), .Z(n21281) );
  CLKBUF_X1 U14640 ( .A(n256101), .Z(n21282) );
  INV_X1 U14641 ( .A(n24775), .ZN(n21283) );
  INV_X1 U14642 ( .A(n25617), .ZN(n21284) );
  INV_X1 U14643 ( .A(n21284), .ZN(n21285) );
  INV_X1 U14644 ( .A(n18234), .ZN(n21286) );
  INV_X1 U14645 ( .A(n18234), .ZN(n21287) );
  INV_X1 U14646 ( .A(n25617), .ZN(n21288) );
  INV_X1 U14647 ( .A(n21288), .ZN(n21289) );
  INV_X1 U14648 ( .A(n18235), .ZN(n21290) );
  INV_X1 U14649 ( .A(n18235), .ZN(n21291) );
  INV_X1 U14650 ( .A(n18236), .ZN(n21292) );
  INV_X1 U14651 ( .A(n18237), .ZN(n21293) );
  INV_X1 U14652 ( .A(n18237), .ZN(n21294) );
  INV_X1 U14653 ( .A(n18238), .ZN(n21295) );
  INV_X1 U14654 ( .A(n18239), .ZN(n21296) );
  INV_X1 U14655 ( .A(n18239), .ZN(n21297) );
  INV_X1 U14656 ( .A(n18240), .ZN(n21298) );
  INV_X1 U14657 ( .A(n18241), .ZN(n21299) );
  INV_X1 U14658 ( .A(n18241), .ZN(n21300) );
  INV_X1 U14659 ( .A(n18242), .ZN(n21301) );
  INV_X1 U14660 ( .A(n18243), .ZN(n21302) );
  INV_X1 U14661 ( .A(n18243), .ZN(n21303) );
  INV_X1 U14662 ( .A(n18244), .ZN(n21304) );
  INV_X1 U14663 ( .A(n18245), .ZN(n21305) );
  INV_X1 U14664 ( .A(n18245), .ZN(n21306) );
  INV_X1 U14665 ( .A(n18246), .ZN(n21307) );
  INV_X1 U14666 ( .A(n18247), .ZN(n21308) );
  INV_X1 U14667 ( .A(n18247), .ZN(n21309) );
  INV_X1 U14668 ( .A(n18248), .ZN(n21310) );
  INV_X1 U14669 ( .A(n18249), .ZN(n21311) );
  INV_X1 U14670 ( .A(n18249), .ZN(n21312) );
  INV_X1 U14671 ( .A(n18250), .ZN(n21313) );
  INV_X1 U14672 ( .A(n18251), .ZN(n21314) );
  INV_X1 U14673 ( .A(n18251), .ZN(n21315) );
  INV_X1 U14674 ( .A(n18252), .ZN(n21316) );
  INV_X1 U14675 ( .A(n18253), .ZN(n21317) );
  INV_X1 U14676 ( .A(n18253), .ZN(n21318) );
  INV_X1 U14677 ( .A(n18254), .ZN(n21319) );
  INV_X1 U14678 ( .A(n18255), .ZN(n21320) );
  INV_X1 U14679 ( .A(n18255), .ZN(n21321) );
  INV_X1 U14680 ( .A(n18256), .ZN(n21322) );
  INV_X1 U14681 ( .A(n18257), .ZN(n21323) );
  INV_X1 U14682 ( .A(n18257), .ZN(n21324) );
  INV_X1 U14683 ( .A(n256301), .ZN(n21325) );
  INV_X1 U14684 ( .A(n21325), .ZN(n21326) );
  INV_X1 U14685 ( .A(n21325), .ZN(n21327) );
  INV_X1 U14686 ( .A(n18258), .ZN(n21328) );
  INV_X1 U14687 ( .A(n21328), .ZN(n21329) );
  INV_X1 U14688 ( .A(n21329), .ZN(n21330) );
  INV_X1 U14689 ( .A(n18258), .ZN(n21331) );
  INV_X1 U14690 ( .A(n18259), .ZN(n21332) );
  INV_X1 U14691 ( .A(n18260), .ZN(n21333) );
  INV_X1 U14692 ( .A(n18260), .ZN(n21334) );
  INV_X1 U14693 ( .A(n38060), .ZN(n21335) );
  INV_X1 U14694 ( .A(n25633), .ZN(n21336) );
  INV_X1 U14695 ( .A(n21336), .ZN(n21337) );
  INV_X1 U14696 ( .A(n21336), .ZN(n21338) );
  INV_X1 U14697 ( .A(n18261), .ZN(n21339) );
  INV_X1 U14698 ( .A(n18262), .ZN(n21340) );
  INV_X1 U14699 ( .A(n18262), .ZN(n21341) );
  INV_X1 U14700 ( .A(n18263), .ZN(n21342) );
  INV_X1 U14701 ( .A(n21342), .ZN(n21343) );
  INV_X1 U14702 ( .A(n18263), .ZN(n21344) );
  INV_X1 U14703 ( .A(n21343), .ZN(n21345) );
  INV_X1 U14704 ( .A(n18264), .ZN(n21346) );
  INV_X1 U14705 ( .A(n18265), .ZN(n21347) );
  INV_X1 U14706 ( .A(n18265), .ZN(n21348) );
  INV_X1 U14707 ( .A(n18266), .ZN(n21349) );
  INV_X1 U14708 ( .A(n18267), .ZN(n21350) );
  INV_X1 U14709 ( .A(n18267), .ZN(n21351) );
  INV_X1 U14710 ( .A(n25639), .ZN(n21352) );
  INV_X1 U14711 ( .A(n21352), .ZN(n21353) );
  INV_X1 U14712 ( .A(n25639), .ZN(n21354) );
  INV_X1 U14713 ( .A(n21353), .ZN(n21355) );
  INV_X1 U14714 ( .A(n18268), .ZN(n21356) );
  INV_X1 U14715 ( .A(n21356), .ZN(n21357) );
  INV_X1 U14716 ( .A(n18268), .ZN(n21358) );
  INV_X1 U14717 ( .A(n21357), .ZN(n21359) );
  INV_X1 U14718 ( .A(n18269), .ZN(n21360) );
  INV_X1 U14719 ( .A(n18270), .ZN(n21361) );
  INV_X1 U14720 ( .A(n18270), .ZN(n21362) );
  INV_X1 U14721 ( .A(n18271), .ZN(n21363) );
  INV_X1 U14722 ( .A(n21363), .ZN(n21364) );
  INV_X1 U14723 ( .A(n18271), .ZN(n21365) );
  INV_X1 U14724 ( .A(n21364), .ZN(n21366) );
  INV_X1 U14725 ( .A(n18950), .ZN(n21367) );
  INV_X1 U14726 ( .A(n21367), .ZN(n21368) );
  INV_X1 U14727 ( .A(n21367), .ZN(n21369) );
  INV_X1 U14728 ( .A(n18949), .ZN(n21370) );
  INV_X1 U14729 ( .A(n21370), .ZN(n21371) );
  INV_X1 U14730 ( .A(n21370), .ZN(n21372) );
  INV_X1 U14731 ( .A(n25644), .ZN(n21373) );
  INV_X1 U14732 ( .A(n21373), .ZN(n21374) );
  INV_X1 U14733 ( .A(n18272), .ZN(n21375) );
  INV_X1 U14734 ( .A(n21375), .ZN(n21376) );
  INV_X1 U14735 ( .A(n18272), .ZN(n21377) );
  INV_X1 U14736 ( .A(n21376), .ZN(n21378) );
  INV_X1 U14737 ( .A(n25651), .ZN(n21379) );
  INV_X1 U14738 ( .A(n21379), .ZN(n21380) );
  INV_X1 U14739 ( .A(n25651), .ZN(n21381) );
  INV_X1 U14740 ( .A(n21380), .ZN(n21382) );
  INV_X1 U14741 ( .A(n25653), .ZN(n21383) );
  INV_X1 U14742 ( .A(n21383), .ZN(n21384) );
  INV_X1 U14743 ( .A(n21384), .ZN(n21385) );
  INV_X1 U14744 ( .A(n25653), .ZN(n21386) );
  INV_X1 U14745 ( .A(n18273), .ZN(n21387) );
  INV_X1 U14746 ( .A(n18273), .ZN(n21388) );
  INV_X1 U14747 ( .A(n18274), .ZN(n21389) );
  INV_X1 U14748 ( .A(n18274), .ZN(n21390) );
  INV_X1 U14749 ( .A(n18275), .ZN(n21391) );
  INV_X1 U14750 ( .A(n18276), .ZN(n21392) );
  INV_X1 U14751 ( .A(n18276), .ZN(n21393) );
  INV_X1 U14752 ( .A(n17133), .ZN(n21394) );
  INV_X1 U14753 ( .A(n21394), .ZN(n21395) );
  INV_X1 U14754 ( .A(n25659), .ZN(n21396) );
  INV_X1 U14755 ( .A(n21396), .ZN(n21397) );
  INV_X1 U14756 ( .A(n21396), .ZN(n21398) );
  INV_X1 U14757 ( .A(n39800), .ZN(n21399) );
  INV_X1 U14758 ( .A(n39800), .ZN(n21400) );
  INV_X1 U14759 ( .A(n256601), .ZN(n21401) );
  INV_X1 U14760 ( .A(n21401), .ZN(n21402) );
  INV_X1 U14761 ( .A(n21401), .ZN(n21403) );
  INV_X1 U14762 ( .A(n18278), .ZN(n21404) );
  INV_X1 U14763 ( .A(n18279), .ZN(n21405) );
  INV_X1 U14764 ( .A(n18280), .ZN(n21406) );
  INV_X1 U14765 ( .A(n18280), .ZN(n21407) );
  INV_X1 U14766 ( .A(n19030), .ZN(n21408) );
  INV_X1 U14767 ( .A(n21408), .ZN(n21409) );
  INV_X1 U14768 ( .A(n21408), .ZN(n21410) );
  INV_X1 U14769 ( .A(n256601), .ZN(n21411) );
  INV_X1 U14770 ( .A(n21411), .ZN(n21412) );
  INV_X1 U14771 ( .A(n21411), .ZN(n21413) );
  INV_X1 U14772 ( .A(n18281), .ZN(n21414) );
  INV_X1 U14773 ( .A(n25832), .ZN(n21415) );
  INV_X1 U14774 ( .A(n21415), .ZN(n21416) );
  INV_X1 U14775 ( .A(n21415), .ZN(n21417) );
  INV_X1 U14776 ( .A(n25846), .ZN(n21418) );
  INV_X1 U14777 ( .A(n21418), .ZN(n21419) );
  INV_X1 U14778 ( .A(n21418), .ZN(n21420) );
  INV_X1 U14779 ( .A(n27221), .ZN(n21421) );
  INV_X1 U14780 ( .A(n21421), .ZN(n21422) );
  INV_X1 U14781 ( .A(n18282), .ZN(n21423) );
  INV_X1 U14782 ( .A(n18282), .ZN(n21424) );
  INV_X1 U14783 ( .A(n26728), .ZN(n21425) );
  INV_X1 U14784 ( .A(n21425), .ZN(n21426) );
  INV_X1 U14785 ( .A(n21425), .ZN(n21427) );
  INV_X1 U14786 ( .A(n24757), .ZN(n21428) );
  INV_X1 U14787 ( .A(n21428), .ZN(n21429) );
  INV_X1 U14788 ( .A(n18283), .ZN(n21430) );
  INV_X1 U14789 ( .A(n18283), .ZN(n21431) );
  INV_X1 U14790 ( .A(n25904), .ZN(n21432) );
  INV_X1 U14791 ( .A(n21432), .ZN(n21433) );
  INV_X1 U14792 ( .A(n21432), .ZN(n21434) );
  INV_X1 U14793 ( .A(n27739), .ZN(n21435) );
  INV_X1 U14794 ( .A(n21435), .ZN(n21436) );
  INV_X1 U14795 ( .A(n21435), .ZN(n21437) );
  INV_X1 U14796 ( .A(n23100), .ZN(n21438) );
  INV_X1 U14797 ( .A(n18284), .ZN(n21439) );
  INV_X1 U14798 ( .A(n18284), .ZN(n21440) );
  INV_X1 U14799 ( .A(n18285), .ZN(n21441) );
  INV_X1 U14800 ( .A(n18285), .ZN(n21442) );
  INV_X1 U14801 ( .A(n18286), .ZN(n21443) );
  INV_X1 U14802 ( .A(n18286), .ZN(n21444) );
  INV_X1 U14803 ( .A(n18287), .ZN(n21445) );
  INV_X1 U14804 ( .A(n18287), .ZN(n21446) );
  INV_X1 U14805 ( .A(n24520), .ZN(n21447) );
  INV_X1 U14806 ( .A(n21447), .ZN(n21448) );
  INV_X1 U14807 ( .A(n21447), .ZN(n21449) );
  INV_X1 U14808 ( .A(n18288), .ZN(n21450) );
  INV_X1 U14809 ( .A(n18288), .ZN(n21451) );
  INV_X1 U14810 ( .A(n18289), .ZN(n21452) );
  INV_X1 U14811 ( .A(n18289), .ZN(n21453) );
  INV_X1 U14812 ( .A(n18290), .ZN(n21454) );
  INV_X1 U14813 ( .A(n18290), .ZN(n21455) );
  INV_X1 U14814 ( .A(n18291), .ZN(n21456) );
  INV_X1 U14815 ( .A(n18291), .ZN(n21457) );
  INV_X1 U14816 ( .A(n18292), .ZN(n21458) );
  INV_X1 U14817 ( .A(n18292), .ZN(n21459) );
  INV_X1 U14818 ( .A(n18293), .ZN(n21460) );
  INV_X1 U14819 ( .A(n18293), .ZN(n21461) );
  INV_X1 U14820 ( .A(n18294), .ZN(n21462) );
  INV_X1 U14821 ( .A(n18294), .ZN(n21463) );
  INV_X1 U14822 ( .A(n22839), .ZN(n21464) );
  INV_X1 U14823 ( .A(n21464), .ZN(n21465) );
  INV_X1 U14824 ( .A(n21464), .ZN(n21466) );
  INV_X1 U14825 ( .A(n18295), .ZN(n21467) );
  INV_X1 U14826 ( .A(n18295), .ZN(n21468) );
  INV_X1 U14827 ( .A(n18296), .ZN(n21469) );
  INV_X1 U14828 ( .A(n18296), .ZN(n21470) );
  INV_X1 U14829 ( .A(n18297), .ZN(n21471) );
  INV_X1 U14830 ( .A(n18297), .ZN(n21472) );
  INV_X1 U14831 ( .A(n18298), .ZN(n21473) );
  INV_X1 U14832 ( .A(n18298), .ZN(n21474) );
  INV_X1 U14833 ( .A(n18299), .ZN(n21475) );
  INV_X1 U14834 ( .A(n18299), .ZN(n21476) );
  INV_X1 U14835 ( .A(n18300), .ZN(n21477) );
  INV_X1 U14836 ( .A(n18300), .ZN(n21478) );
  INV_X1 U14837 ( .A(n18301), .ZN(n21479) );
  INV_X1 U14838 ( .A(n18301), .ZN(n21480) );
  INV_X1 U14839 ( .A(n18302), .ZN(n21481) );
  INV_X1 U14840 ( .A(n18302), .ZN(n21482) );
  INV_X1 U14841 ( .A(n18303), .ZN(n21483) );
  INV_X1 U14842 ( .A(n18303), .ZN(n21484) );
  INV_X1 U14843 ( .A(n18304), .ZN(n21485) );
  INV_X1 U14844 ( .A(n18304), .ZN(n21486) );
  INV_X1 U14845 ( .A(n18305), .ZN(n21487) );
  INV_X1 U14846 ( .A(n18305), .ZN(n21488) );
  INV_X1 U14847 ( .A(n18306), .ZN(n21489) );
  INV_X1 U14848 ( .A(n18306), .ZN(n21490) );
  INV_X1 U14849 ( .A(n18307), .ZN(n21491) );
  INV_X1 U14850 ( .A(n18307), .ZN(n21492) );
  INV_X1 U14851 ( .A(n18308), .ZN(n21493) );
  INV_X1 U14852 ( .A(n18308), .ZN(n21494) );
  INV_X1 U14853 ( .A(n18309), .ZN(n21495) );
  INV_X1 U14854 ( .A(n18309), .ZN(n21496) );
  INV_X1 U14855 ( .A(n18310), .ZN(n21497) );
  INV_X1 U14856 ( .A(n18310), .ZN(n21498) );
  INV_X1 U14857 ( .A(n18311), .ZN(n21499) );
  INV_X1 U14858 ( .A(n18311), .ZN(n21500) );
  INV_X1 U14859 ( .A(n22828), .ZN(n21501) );
  INV_X1 U14860 ( .A(n21501), .ZN(n21502) );
  INV_X1 U14861 ( .A(n21501), .ZN(n21503) );
  INV_X1 U14862 ( .A(n18312), .ZN(n21504) );
  INV_X1 U14863 ( .A(n18312), .ZN(n21505) );
  INV_X1 U14864 ( .A(n18313), .ZN(n21506) );
  INV_X1 U14865 ( .A(n18313), .ZN(n21507) );
  INV_X1 U14866 ( .A(n18314), .ZN(n21508) );
  INV_X1 U14867 ( .A(n18314), .ZN(n21509) );
  INV_X1 U14868 ( .A(n18315), .ZN(n21510) );
  INV_X1 U14869 ( .A(n18315), .ZN(n21511) );
  INV_X1 U14870 ( .A(n18316), .ZN(n21512) );
  INV_X1 U14871 ( .A(n18316), .ZN(n21513) );
  INV_X1 U14872 ( .A(n26086), .ZN(n21514) );
  INV_X1 U14873 ( .A(n21514), .ZN(n21515) );
  INV_X1 U14874 ( .A(n21514), .ZN(n21516) );
  INV_X1 U14875 ( .A(n23221), .ZN(n21517) );
  INV_X1 U14876 ( .A(n18317), .ZN(n21518) );
  INV_X1 U14877 ( .A(n18317), .ZN(n21519) );
  INV_X1 U14878 ( .A(n18318), .ZN(n21520) );
  INV_X1 U14879 ( .A(n18318), .ZN(n21521) );
  INV_X1 U14880 ( .A(n18319), .ZN(n21522) );
  INV_X1 U14881 ( .A(n18319), .ZN(n21523) );
  INV_X1 U14882 ( .A(n26086), .ZN(n21524) );
  INV_X1 U14883 ( .A(n21524), .ZN(n21525) );
  INV_X1 U14884 ( .A(n21524), .ZN(n21526) );
  INV_X1 U14885 ( .A(n18320), .ZN(n21527) );
  INV_X1 U14886 ( .A(n18320), .ZN(n21528) );
  INV_X1 U14887 ( .A(n18321), .ZN(n21529) );
  INV_X1 U14888 ( .A(n18321), .ZN(n21530) );
  INV_X1 U14889 ( .A(n18322), .ZN(n21531) );
  INV_X1 U14890 ( .A(n18322), .ZN(n21532) );
  INV_X1 U14891 ( .A(n18323), .ZN(n21533) );
  INV_X1 U14892 ( .A(n18323), .ZN(n21534) );
  INV_X1 U14893 ( .A(n26097), .ZN(n21535) );
  INV_X1 U14894 ( .A(n21535), .ZN(n21536) );
  INV_X1 U14895 ( .A(n21535), .ZN(n21537) );
  INV_X1 U14896 ( .A(n18324), .ZN(n21538) );
  INV_X1 U14897 ( .A(n18324), .ZN(n21539) );
  INV_X1 U14898 ( .A(n18325), .ZN(n21540) );
  INV_X1 U14899 ( .A(n18325), .ZN(n21541) );
  INV_X1 U14900 ( .A(n26097), .ZN(n21542) );
  INV_X1 U14901 ( .A(n21542), .ZN(n21543) );
  INV_X1 U14902 ( .A(n21542), .ZN(n21544) );
  INV_X1 U14903 ( .A(n23234), .ZN(n21545) );
  INV_X1 U14904 ( .A(n23235), .ZN(n21546) );
  INV_X1 U14905 ( .A(n18326), .ZN(n21547) );
  INV_X1 U14906 ( .A(n18326), .ZN(n21548) );
  INV_X1 U14907 ( .A(n18327), .ZN(n21549) );
  INV_X1 U14908 ( .A(n18327), .ZN(n21550) );
  INV_X1 U14909 ( .A(n18328), .ZN(n21551) );
  INV_X1 U14910 ( .A(n18328), .ZN(n21552) );
  INV_X1 U14911 ( .A(n18329), .ZN(n21553) );
  INV_X1 U14912 ( .A(n18329), .ZN(n21554) );
  INV_X1 U14913 ( .A(n18330), .ZN(n21555) );
  INV_X1 U14914 ( .A(n18330), .ZN(n21556) );
  INV_X1 U14915 ( .A(n18331), .ZN(n21557) );
  INV_X1 U14916 ( .A(n18331), .ZN(n21558) );
  INV_X1 U14917 ( .A(n18332), .ZN(n21559) );
  INV_X1 U14918 ( .A(n18332), .ZN(n21560) );
  INV_X1 U14919 ( .A(n18333), .ZN(n21561) );
  INV_X1 U14920 ( .A(n18333), .ZN(n21562) );
  INV_X1 U14921 ( .A(n18334), .ZN(n21563) );
  INV_X1 U14922 ( .A(n18334), .ZN(n21564) );
  INV_X1 U14923 ( .A(n18335), .ZN(n21565) );
  INV_X1 U14924 ( .A(n18335), .ZN(n21566) );
  INV_X1 U14925 ( .A(n18336), .ZN(n21567) );
  INV_X1 U14926 ( .A(n18336), .ZN(n21568) );
  INV_X1 U14927 ( .A(n18337), .ZN(n21569) );
  INV_X1 U14928 ( .A(n18337), .ZN(n21570) );
  INV_X1 U14929 ( .A(n18338), .ZN(n21571) );
  INV_X1 U14930 ( .A(n18338), .ZN(n21572) );
  INV_X1 U14931 ( .A(n18339), .ZN(n21573) );
  INV_X1 U14932 ( .A(n18339), .ZN(n21574) );
  INV_X1 U14933 ( .A(n18340), .ZN(n21575) );
  INV_X1 U14934 ( .A(n18340), .ZN(n21576) );
  INV_X1 U14935 ( .A(n18341), .ZN(n21577) );
  INV_X1 U14936 ( .A(n18341), .ZN(n21578) );
  INV_X1 U14937 ( .A(n18342), .ZN(n21579) );
  INV_X1 U14938 ( .A(n18342), .ZN(n21580) );
  INV_X1 U14939 ( .A(n18343), .ZN(n21581) );
  INV_X1 U14940 ( .A(n18343), .ZN(n21582) );
  INV_X1 U14941 ( .A(n18344), .ZN(n21583) );
  INV_X1 U14942 ( .A(n18344), .ZN(n21584) );
  INV_X1 U14943 ( .A(n18345), .ZN(n21585) );
  INV_X1 U14944 ( .A(n18345), .ZN(n21586) );
  INV_X1 U14945 ( .A(n18346), .ZN(n21587) );
  INV_X1 U14946 ( .A(n18346), .ZN(n21588) );
  INV_X1 U14947 ( .A(n18347), .ZN(n21589) );
  INV_X1 U14948 ( .A(n18347), .ZN(n21590) );
  INV_X1 U14949 ( .A(n18348), .ZN(n21591) );
  INV_X1 U14950 ( .A(n18348), .ZN(n21592) );
  INV_X1 U14951 ( .A(n18349), .ZN(n21593) );
  INV_X1 U14952 ( .A(n18349), .ZN(n21594) );
  INV_X1 U14953 ( .A(n4715), .ZN(n21595) );
  INV_X1 U14954 ( .A(n21595), .ZN(n21596) );
  INV_X1 U14955 ( .A(n21595), .ZN(n21597) );
  INV_X1 U14956 ( .A(n26378), .ZN(n21598) );
  INV_X1 U14957 ( .A(n21598), .ZN(n21599) );
  INV_X1 U14958 ( .A(n21598), .ZN(n21600) );
  INV_X1 U14959 ( .A(n4716), .ZN(n21601) );
  INV_X1 U14960 ( .A(n21601), .ZN(n21602) );
  INV_X1 U14961 ( .A(n21601), .ZN(n21603) );
  INV_X1 U14962 ( .A(n26367), .ZN(n21604) );
  INV_X1 U14963 ( .A(n21604), .ZN(n21605) );
  INV_X1 U14964 ( .A(n21604), .ZN(n21606) );
  INV_X1 U14965 ( .A(n18350), .ZN(n21607) );
  INV_X1 U14966 ( .A(n18350), .ZN(n21608) );
  INV_X1 U14967 ( .A(n18351), .ZN(n21609) );
  INV_X1 U14968 ( .A(n18351), .ZN(n21610) );
  INV_X1 U14969 ( .A(n18352), .ZN(n21611) );
  INV_X1 U14970 ( .A(n18352), .ZN(n21612) );
  INV_X1 U14971 ( .A(n18353), .ZN(n21613) );
  INV_X1 U14972 ( .A(n18353), .ZN(n21614) );
  INV_X1 U14973 ( .A(n18354), .ZN(n21615) );
  INV_X1 U14974 ( .A(n18354), .ZN(n21616) );
  INV_X1 U14975 ( .A(n20564), .ZN(n21617) );
  INV_X1 U14976 ( .A(n21617), .ZN(n21618) );
  INV_X1 U14977 ( .A(n21617), .ZN(n21619) );
  INV_X1 U14978 ( .A(n18355), .ZN(n21620) );
  INV_X1 U14979 ( .A(n18355), .ZN(n21621) );
  INV_X1 U14980 ( .A(n20559), .ZN(n21622) );
  INV_X1 U14981 ( .A(n21622), .ZN(n21623) );
  INV_X1 U14982 ( .A(n21622), .ZN(n21624) );
  INV_X1 U14983 ( .A(n18356), .ZN(n21625) );
  INV_X1 U14984 ( .A(n18356), .ZN(n21626) );
  INV_X1 U14985 ( .A(n18357), .ZN(n21627) );
  INV_X1 U14986 ( .A(n18357), .ZN(n21628) );
  INV_X1 U14987 ( .A(n18358), .ZN(n21629) );
  INV_X1 U14988 ( .A(n18358), .ZN(n21630) );
  INV_X1 U14989 ( .A(n18359), .ZN(n21631) );
  INV_X1 U14990 ( .A(n18359), .ZN(n21632) );
  INV_X1 U14991 ( .A(n18360), .ZN(n21633) );
  INV_X1 U14992 ( .A(n18360), .ZN(n21634) );
  INV_X1 U14993 ( .A(n18361), .ZN(n21635) );
  INV_X1 U14994 ( .A(n18361), .ZN(n21636) );
  INV_X1 U14995 ( .A(n18362), .ZN(n21637) );
  INV_X1 U14996 ( .A(n18362), .ZN(n21638) );
  INV_X1 U14997 ( .A(n18363), .ZN(n21639) );
  INV_X1 U14998 ( .A(n18363), .ZN(n21640) );
  INV_X1 U14999 ( .A(n18364), .ZN(n21641) );
  INV_X1 U15000 ( .A(n18364), .ZN(n21642) );
  INV_X1 U15001 ( .A(n18365), .ZN(n21643) );
  INV_X1 U15002 ( .A(n18365), .ZN(n21644) );
  INV_X1 U15003 ( .A(n18366), .ZN(n21645) );
  INV_X1 U15004 ( .A(n18366), .ZN(n21646) );
  INV_X1 U15005 ( .A(n18367), .ZN(n21647) );
  INV_X1 U15006 ( .A(n18367), .ZN(n21648) );
  INV_X1 U15007 ( .A(n394), .ZN(n21649) );
  INV_X1 U15008 ( .A(n394), .ZN(n21650) );
  INV_X1 U15009 ( .A(n18368), .ZN(n21651) );
  INV_X1 U15010 ( .A(n18368), .ZN(n21652) );
  INV_X1 U15011 ( .A(n18369), .ZN(n21653) );
  INV_X1 U15012 ( .A(n18369), .ZN(n21654) );
  INV_X1 U15013 ( .A(n393), .ZN(n21655) );
  INV_X1 U15014 ( .A(n393), .ZN(n21656) );
  INV_X1 U15015 ( .A(n392), .ZN(n21657) );
  INV_X1 U15016 ( .A(n392), .ZN(n21658) );
  INV_X1 U15017 ( .A(n391), .ZN(n21659) );
  INV_X1 U15018 ( .A(n391), .ZN(n21660) );
  INV_X1 U15019 ( .A(n390), .ZN(n21661) );
  INV_X1 U15020 ( .A(n390), .ZN(n21662) );
  INV_X1 U15021 ( .A(n389), .ZN(n21663) );
  INV_X1 U15022 ( .A(n389), .ZN(n21664) );
  INV_X1 U15023 ( .A(n388), .ZN(n21665) );
  INV_X1 U15024 ( .A(n388), .ZN(n21666) );
  INV_X1 U15025 ( .A(n387), .ZN(n21667) );
  INV_X1 U15026 ( .A(n387), .ZN(n21668) );
  INV_X1 U15027 ( .A(n386), .ZN(n21669) );
  INV_X1 U15028 ( .A(n386), .ZN(n21670) );
  INV_X1 U15029 ( .A(n385), .ZN(n21671) );
  INV_X1 U15030 ( .A(n385), .ZN(n21672) );
  INV_X1 U15031 ( .A(n384), .ZN(n21673) );
  INV_X1 U15032 ( .A(n384), .ZN(n21674) );
  INV_X1 U15033 ( .A(n383), .ZN(n21675) );
  INV_X1 U15034 ( .A(n383), .ZN(n21676) );
  INV_X1 U15035 ( .A(n382), .ZN(n21677) );
  INV_X1 U15036 ( .A(n382), .ZN(n21678) );
  INV_X1 U15037 ( .A(n381), .ZN(n21679) );
  INV_X1 U15038 ( .A(n381), .ZN(n21680) );
  INV_X1 U15039 ( .A(n380), .ZN(n21681) );
  INV_X1 U15040 ( .A(n380), .ZN(n21682) );
  INV_X1 U15041 ( .A(n379), .ZN(n21683) );
  INV_X1 U15042 ( .A(n379), .ZN(n21684) );
  INV_X1 U15043 ( .A(n378), .ZN(n21685) );
  INV_X1 U15044 ( .A(n378), .ZN(n21686) );
  INV_X1 U15045 ( .A(n377), .ZN(n21687) );
  INV_X1 U15046 ( .A(n377), .ZN(n21688) );
  INV_X1 U15047 ( .A(n376), .ZN(n21689) );
  INV_X1 U15048 ( .A(n376), .ZN(n21690) );
  INV_X1 U15049 ( .A(n375), .ZN(n21691) );
  INV_X1 U15050 ( .A(n375), .ZN(n21692) );
  INV_X1 U15051 ( .A(n374), .ZN(n21693) );
  INV_X1 U15052 ( .A(n374), .ZN(n21694) );
  INV_X1 U15053 ( .A(n373), .ZN(n21695) );
  INV_X1 U15054 ( .A(n373), .ZN(n21696) );
  INV_X1 U15055 ( .A(n372), .ZN(n21697) );
  INV_X1 U15056 ( .A(n372), .ZN(n21698) );
  INV_X1 U15057 ( .A(n371), .ZN(n21699) );
  INV_X1 U15058 ( .A(n371), .ZN(n21700) );
  INV_X1 U15059 ( .A(n370), .ZN(n21701) );
  INV_X1 U15060 ( .A(n370), .ZN(n21702) );
  INV_X1 U15061 ( .A(n369), .ZN(n21703) );
  INV_X1 U15062 ( .A(n369), .ZN(n21704) );
  INV_X1 U15063 ( .A(n368), .ZN(n21705) );
  INV_X1 U15064 ( .A(n368), .ZN(n21706) );
  INV_X1 U15065 ( .A(n367), .ZN(n21707) );
  INV_X1 U15066 ( .A(n367), .ZN(n21708) );
  INV_X1 U15067 ( .A(n366), .ZN(n21709) );
  INV_X1 U15068 ( .A(n366), .ZN(n21710) );
  INV_X1 U15069 ( .A(n365), .ZN(n21711) );
  INV_X1 U15070 ( .A(n365), .ZN(n21712) );
  INV_X1 U15071 ( .A(n364), .ZN(n21713) );
  INV_X1 U15072 ( .A(n364), .ZN(n21714) );
  INV_X1 U15073 ( .A(n363), .ZN(n21715) );
  INV_X1 U15074 ( .A(n363), .ZN(n21716) );
  INV_X1 U15075 ( .A(n362), .ZN(n21717) );
  INV_X1 U15076 ( .A(n362), .ZN(n21718) );
  INV_X1 U15077 ( .A(n361), .ZN(n21719) );
  INV_X1 U15078 ( .A(n361), .ZN(n21720) );
  INV_X1 U15079 ( .A(n360), .ZN(n21721) );
  INV_X1 U15080 ( .A(n360), .ZN(n21722) );
  INV_X1 U15081 ( .A(n359), .ZN(n21723) );
  INV_X1 U15082 ( .A(n359), .ZN(n21724) );
  INV_X1 U15083 ( .A(n358), .ZN(n21725) );
  INV_X1 U15084 ( .A(n358), .ZN(n21726) );
  INV_X1 U15085 ( .A(n357), .ZN(n21727) );
  INV_X1 U15086 ( .A(n357), .ZN(n21728) );
  INV_X1 U15087 ( .A(n356), .ZN(n21729) );
  INV_X1 U15088 ( .A(n356), .ZN(n21730) );
  INV_X1 U15089 ( .A(n355), .ZN(n21731) );
  INV_X1 U15090 ( .A(n355), .ZN(n21732) );
  INV_X1 U15091 ( .A(n354), .ZN(n21733) );
  INV_X1 U15092 ( .A(n354), .ZN(n21734) );
  INV_X1 U15093 ( .A(n353), .ZN(n21735) );
  INV_X1 U15094 ( .A(n353), .ZN(n21736) );
  INV_X1 U15095 ( .A(n352), .ZN(n21737) );
  INV_X1 U15096 ( .A(n352), .ZN(n21738) );
  INV_X1 U15097 ( .A(n351), .ZN(n21739) );
  INV_X1 U15098 ( .A(n351), .ZN(n21740) );
  INV_X1 U15099 ( .A(n350), .ZN(n21741) );
  INV_X1 U15100 ( .A(n350), .ZN(n21742) );
  INV_X1 U15101 ( .A(n349), .ZN(n21743) );
  INV_X1 U15102 ( .A(n349), .ZN(n21744) );
  INV_X1 U15103 ( .A(n348), .ZN(n21745) );
  INV_X1 U15104 ( .A(n348), .ZN(n21746) );
  INV_X1 U15105 ( .A(n347), .ZN(n21747) );
  INV_X1 U15106 ( .A(n347), .ZN(n21748) );
  INV_X1 U15107 ( .A(n346), .ZN(n21749) );
  INV_X1 U15108 ( .A(n346), .ZN(n21750) );
  INV_X1 U15109 ( .A(n345), .ZN(n21751) );
  INV_X1 U15110 ( .A(n345), .ZN(n21752) );
  INV_X1 U15111 ( .A(n344), .ZN(n21753) );
  INV_X1 U15112 ( .A(n344), .ZN(n21754) );
  INV_X1 U15113 ( .A(n343), .ZN(n21755) );
  INV_X1 U15114 ( .A(n343), .ZN(n21756) );
  INV_X1 U15115 ( .A(n342), .ZN(n21757) );
  INV_X1 U15116 ( .A(n342), .ZN(n21758) );
  INV_X1 U15117 ( .A(n341), .ZN(n21759) );
  INV_X1 U15118 ( .A(n341), .ZN(n21760) );
  INV_X1 U15119 ( .A(n340), .ZN(n21761) );
  INV_X1 U15120 ( .A(n340), .ZN(n21762) );
  INV_X1 U15121 ( .A(n339), .ZN(n21763) );
  INV_X1 U15122 ( .A(n339), .ZN(n21764) );
  INV_X1 U15123 ( .A(n338), .ZN(n21765) );
  INV_X1 U15124 ( .A(n338), .ZN(n21766) );
  INV_X1 U15125 ( .A(n337), .ZN(n21767) );
  INV_X1 U15126 ( .A(n337), .ZN(n21768) );
  INV_X1 U15127 ( .A(n336), .ZN(n21769) );
  INV_X1 U15128 ( .A(n336), .ZN(n21770) );
  INV_X1 U15129 ( .A(n335), .ZN(n21771) );
  INV_X1 U15130 ( .A(n335), .ZN(n21772) );
  INV_X1 U15131 ( .A(n334), .ZN(n21773) );
  INV_X1 U15132 ( .A(n334), .ZN(n21774) );
  INV_X1 U15133 ( .A(n18370), .ZN(n21775) );
  INV_X1 U15134 ( .A(n18370), .ZN(n21776) );
  INV_X1 U15135 ( .A(n18371), .ZN(n21777) );
  INV_X1 U15136 ( .A(n18371), .ZN(n21778) );
  INV_X1 U15137 ( .A(n18372), .ZN(n21779) );
  INV_X1 U15138 ( .A(n18372), .ZN(n21780) );
  INV_X1 U15139 ( .A(n18373), .ZN(n21781) );
  INV_X1 U15140 ( .A(n18373), .ZN(n21782) );
  INV_X1 U15141 ( .A(n18374), .ZN(n21783) );
  INV_X1 U15142 ( .A(n18374), .ZN(n21784) );
  INV_X1 U15143 ( .A(n18375), .ZN(n21785) );
  INV_X1 U15144 ( .A(n18375), .ZN(n21786) );
  INV_X1 U15145 ( .A(n18376), .ZN(n21787) );
  INV_X1 U15146 ( .A(n18376), .ZN(n21788) );
  INV_X1 U15147 ( .A(n18377), .ZN(n21789) );
  INV_X1 U15148 ( .A(n18377), .ZN(n21790) );
  INV_X1 U15149 ( .A(n18378), .ZN(n21791) );
  INV_X1 U15150 ( .A(n18378), .ZN(n21792) );
  INV_X1 U15151 ( .A(n18379), .ZN(n21793) );
  INV_X1 U15152 ( .A(n18379), .ZN(n21794) );
  INV_X1 U15153 ( .A(n18380), .ZN(n21795) );
  INV_X1 U15154 ( .A(n18380), .ZN(n21796) );
  INV_X1 U15155 ( .A(n18381), .ZN(n21797) );
  INV_X1 U15156 ( .A(n18381), .ZN(n21798) );
  INV_X1 U15157 ( .A(n18382), .ZN(n21799) );
  INV_X1 U15158 ( .A(n18382), .ZN(n21800) );
  INV_X1 U15159 ( .A(n18383), .ZN(n21801) );
  INV_X1 U15160 ( .A(n18383), .ZN(n21802) );
  INV_X1 U15161 ( .A(n18384), .ZN(n21803) );
  INV_X1 U15162 ( .A(n18384), .ZN(n21804) );
  INV_X1 U15163 ( .A(n18385), .ZN(n21805) );
  INV_X1 U15164 ( .A(n18385), .ZN(n21806) );
  INV_X1 U15165 ( .A(n18386), .ZN(n21807) );
  INV_X1 U15166 ( .A(n18386), .ZN(n21808) );
  INV_X1 U15167 ( .A(n18387), .ZN(n21809) );
  INV_X1 U15168 ( .A(n18387), .ZN(n21810) );
  INV_X1 U15169 ( .A(n18388), .ZN(n21811) );
  INV_X1 U15170 ( .A(n18388), .ZN(n21812) );
  INV_X1 U15171 ( .A(n18389), .ZN(n21813) );
  INV_X1 U15172 ( .A(n18389), .ZN(n21814) );
  INV_X1 U15173 ( .A(n18390), .ZN(n21815) );
  INV_X1 U15174 ( .A(n18390), .ZN(n21816) );
  INV_X1 U15175 ( .A(n18391), .ZN(n21817) );
  INV_X1 U15176 ( .A(n18391), .ZN(n21818) );
  INV_X1 U15177 ( .A(n18392), .ZN(n21819) );
  INV_X1 U15178 ( .A(n18392), .ZN(n21820) );
  INV_X1 U15179 ( .A(n18393), .ZN(n21821) );
  INV_X1 U15180 ( .A(n18393), .ZN(n21822) );
  INV_X1 U15181 ( .A(n18394), .ZN(n21823) );
  INV_X1 U15182 ( .A(n18394), .ZN(n21824) );
  INV_X1 U15183 ( .A(n18395), .ZN(n21825) );
  INV_X1 U15184 ( .A(n18395), .ZN(n21826) );
  INV_X1 U15185 ( .A(n18396), .ZN(n21827) );
  INV_X1 U15186 ( .A(n18396), .ZN(n21828) );
  INV_X1 U15187 ( .A(n18397), .ZN(n21829) );
  INV_X1 U15188 ( .A(n18397), .ZN(n21830) );
  INV_X1 U15189 ( .A(n18398), .ZN(n21831) );
  INV_X1 U15190 ( .A(n18398), .ZN(n21832) );
  INV_X1 U15191 ( .A(n18399), .ZN(n21833) );
  INV_X1 U15192 ( .A(n18399), .ZN(n21834) );
  INV_X1 U15193 ( .A(n18400), .ZN(n21835) );
  INV_X1 U15194 ( .A(n18400), .ZN(n21836) );
  INV_X1 U15195 ( .A(n18401), .ZN(n21837) );
  INV_X1 U15196 ( .A(n18401), .ZN(n21838) );
  INV_X1 U15197 ( .A(n18402), .ZN(n21839) );
  INV_X1 U15198 ( .A(n18402), .ZN(n21840) );
  INV_X1 U15199 ( .A(n18403), .ZN(n21841) );
  INV_X1 U15200 ( .A(n18403), .ZN(n21842) );
  INV_X1 U15201 ( .A(n18404), .ZN(n21843) );
  INV_X1 U15202 ( .A(n18404), .ZN(n21844) );
  INV_X1 U15203 ( .A(n18405), .ZN(n21845) );
  INV_X1 U15204 ( .A(n18405), .ZN(n21846) );
  INV_X1 U15205 ( .A(n18406), .ZN(n21847) );
  INV_X1 U15206 ( .A(n18406), .ZN(n21848) );
  INV_X1 U15207 ( .A(n18407), .ZN(n21849) );
  INV_X1 U15208 ( .A(n18407), .ZN(n21850) );
  INV_X1 U15209 ( .A(n18408), .ZN(n21851) );
  INV_X1 U15210 ( .A(n18408), .ZN(n21852) );
  INV_X1 U15211 ( .A(n18409), .ZN(n21853) );
  INV_X1 U15212 ( .A(n18409), .ZN(n21854) );
  INV_X1 U15213 ( .A(n18410), .ZN(n21855) );
  INV_X1 U15214 ( .A(n18410), .ZN(n21856) );
  INV_X1 U15215 ( .A(n18411), .ZN(n21857) );
  INV_X1 U15216 ( .A(n18411), .ZN(n21858) );
  INV_X1 U15217 ( .A(n18412), .ZN(n21859) );
  INV_X1 U15218 ( .A(n18412), .ZN(n21860) );
  INV_X1 U15219 ( .A(n18413), .ZN(n21861) );
  INV_X1 U15220 ( .A(n18413), .ZN(n21862) );
  INV_X1 U15221 ( .A(n18414), .ZN(n21863) );
  INV_X1 U15222 ( .A(n18414), .ZN(n21864) );
  INV_X1 U15223 ( .A(n19752), .ZN(n21865) );
  INV_X1 U15224 ( .A(n21865), .ZN(n21866) );
  INV_X1 U15225 ( .A(n21865), .ZN(n21867) );
  INV_X1 U15226 ( .A(n18415), .ZN(n21868) );
  INV_X1 U15227 ( .A(n18415), .ZN(n21869) );
  INV_X1 U15228 ( .A(n18416), .ZN(n21870) );
  INV_X1 U15229 ( .A(n18416), .ZN(n21871) );
  INV_X1 U15230 ( .A(n18417), .ZN(n21872) );
  INV_X1 U15231 ( .A(n18417), .ZN(n21873) );
  INV_X1 U15232 ( .A(n26327), .ZN(n21874) );
  INV_X1 U15233 ( .A(n21874), .ZN(n21875) );
  INV_X1 U15234 ( .A(n21874), .ZN(n21876) );
  INV_X1 U15235 ( .A(n18418), .ZN(n21877) );
  INV_X1 U15236 ( .A(n18418), .ZN(n21878) );
  INV_X1 U15237 ( .A(n26331), .ZN(n21879) );
  INV_X1 U15238 ( .A(n21879), .ZN(n21880) );
  INV_X1 U15239 ( .A(n21879), .ZN(n21881) );
  INV_X1 U15240 ( .A(n18419), .ZN(n21882) );
  INV_X1 U15241 ( .A(n18419), .ZN(n21883) );
  INV_X1 U15242 ( .A(n26334), .ZN(n21884) );
  INV_X1 U15243 ( .A(n21884), .ZN(n21885) );
  INV_X1 U15244 ( .A(n21884), .ZN(n21886) );
  INV_X1 U15245 ( .A(n18420), .ZN(n21887) );
  INV_X1 U15246 ( .A(n18420), .ZN(n21888) );
  INV_X1 U15247 ( .A(n26336), .ZN(n21889) );
  INV_X1 U15248 ( .A(n21889), .ZN(n21890) );
  INV_X1 U15249 ( .A(n21889), .ZN(n21891) );
  INV_X1 U15250 ( .A(n18421), .ZN(n21892) );
  INV_X1 U15251 ( .A(n18421), .ZN(n21893) );
  INV_X1 U15252 ( .A(n26340), .ZN(n21894) );
  INV_X1 U15253 ( .A(n21894), .ZN(n21895) );
  INV_X1 U15254 ( .A(n21894), .ZN(n21896) );
  INV_X1 U15255 ( .A(n18422), .ZN(n21897) );
  INV_X1 U15256 ( .A(n18422), .ZN(n21898) );
  INV_X1 U15257 ( .A(n26342), .ZN(n21899) );
  INV_X1 U15258 ( .A(n21899), .ZN(n21900) );
  INV_X1 U15259 ( .A(n21899), .ZN(n21901) );
  INV_X1 U15260 ( .A(n18423), .ZN(n21902) );
  INV_X1 U15261 ( .A(n18423), .ZN(n21903) );
  INV_X1 U15262 ( .A(n26345), .ZN(n21904) );
  INV_X1 U15263 ( .A(n21904), .ZN(n21905) );
  INV_X1 U15264 ( .A(n21904), .ZN(n21906) );
  INV_X1 U15265 ( .A(n18424), .ZN(n21907) );
  INV_X1 U15266 ( .A(n18424), .ZN(n21908) );
  INV_X1 U15267 ( .A(n26348), .ZN(n21909) );
  INV_X1 U15268 ( .A(n21909), .ZN(n21910) );
  INV_X1 U15269 ( .A(n21909), .ZN(n21911) );
  INV_X1 U15270 ( .A(n18425), .ZN(n21912) );
  INV_X1 U15271 ( .A(n18425), .ZN(n21913) );
  INV_X1 U15272 ( .A(n26351), .ZN(n21914) );
  INV_X1 U15273 ( .A(n21914), .ZN(n21915) );
  INV_X1 U15274 ( .A(n21914), .ZN(n21916) );
  INV_X1 U15275 ( .A(n18426), .ZN(n21917) );
  INV_X1 U15276 ( .A(n18426), .ZN(n21918) );
  INV_X1 U15277 ( .A(n26354), .ZN(n21919) );
  INV_X1 U15278 ( .A(n21919), .ZN(n21920) );
  INV_X1 U15279 ( .A(n21919), .ZN(n21921) );
  INV_X1 U15280 ( .A(n18427), .ZN(n21922) );
  INV_X1 U15281 ( .A(n18427), .ZN(n21923) );
  INV_X1 U15282 ( .A(n26357), .ZN(n21924) );
  INV_X1 U15283 ( .A(n21924), .ZN(n21925) );
  INV_X1 U15284 ( .A(n21924), .ZN(n21926) );
  INV_X1 U15285 ( .A(n18428), .ZN(n21927) );
  INV_X1 U15286 ( .A(n18428), .ZN(n21928) );
  INV_X1 U15287 ( .A(n26360), .ZN(n21929) );
  INV_X1 U15288 ( .A(n21929), .ZN(n21930) );
  INV_X1 U15289 ( .A(n21929), .ZN(n21931) );
  INV_X1 U15290 ( .A(n18429), .ZN(n21932) );
  INV_X1 U15291 ( .A(n18429), .ZN(n21933) );
  INV_X1 U15292 ( .A(n26363), .ZN(n21934) );
  INV_X1 U15293 ( .A(n21934), .ZN(n21935) );
  INV_X1 U15294 ( .A(n21934), .ZN(n21936) );
  INV_X1 U15295 ( .A(n26367), .ZN(n21937) );
  INV_X1 U15296 ( .A(n21937), .ZN(n21938) );
  INV_X1 U15297 ( .A(n21937), .ZN(n21939) );
  INV_X1 U15298 ( .A(n18430), .ZN(n21940) );
  INV_X1 U15299 ( .A(n18430), .ZN(n21941) );
  INV_X1 U15300 ( .A(n263701), .ZN(n21942) );
  INV_X1 U15301 ( .A(n21942), .ZN(n21943) );
  INV_X1 U15302 ( .A(n21942), .ZN(n21944) );
  CLKBUF_X1 U15303 ( .A(n26374), .Z(n21945) );
  INV_X1 U15304 ( .A(n26378), .ZN(n21946) );
  INV_X1 U15305 ( .A(n21946), .ZN(n21947) );
  INV_X1 U15306 ( .A(n21946), .ZN(n21948) );
  INV_X1 U15307 ( .A(n20975), .ZN(n21949) );
  INV_X1 U15308 ( .A(n20981), .ZN(n21950) );
  INV_X1 U15309 ( .A(n18432), .ZN(n21951) );
  INV_X1 U15310 ( .A(n18432), .ZN(n21952) );
  INV_X1 U15311 ( .A(n18433), .ZN(n21953) );
  INV_X1 U15312 ( .A(n18433), .ZN(n21954) );
  INV_X1 U15313 ( .A(n20973), .ZN(n21955) );
  INV_X1 U15314 ( .A(n20983), .ZN(n21956) );
  INV_X1 U15315 ( .A(n18434), .ZN(n21957) );
  INV_X1 U15316 ( .A(n18434), .ZN(n21958) );
  INV_X1 U15317 ( .A(n18435), .ZN(n21959) );
  INV_X1 U15318 ( .A(n18435), .ZN(n21960) );
  INV_X1 U15319 ( .A(n20978), .ZN(n21961) );
  INV_X1 U15320 ( .A(n20985), .ZN(n21962) );
  INV_X1 U15321 ( .A(n18436), .ZN(n21963) );
  INV_X1 U15322 ( .A(n18436), .ZN(n21964) );
  INV_X1 U15323 ( .A(n21954), .ZN(n21965) );
  INV_X1 U15324 ( .A(n20989), .ZN(n21966) );
  INV_X1 U15325 ( .A(n18437), .ZN(n21967) );
  INV_X1 U15326 ( .A(n18437), .ZN(n21968) );
  INV_X1 U15327 ( .A(n26400), .ZN(n21969) );
  INV_X1 U15328 ( .A(n21969), .ZN(n21970) );
  INV_X1 U15329 ( .A(n21969), .ZN(n21971) );
  INV_X1 U15330 ( .A(n18438), .ZN(n21972) );
  INV_X1 U15331 ( .A(n18438), .ZN(n21973) );
  INV_X1 U15332 ( .A(n26403), .ZN(n21974) );
  INV_X1 U15333 ( .A(n21974), .ZN(n21975) );
  INV_X1 U15334 ( .A(n21974), .ZN(n21976) );
  INV_X1 U15335 ( .A(n333), .ZN(n21977) );
  INV_X1 U15336 ( .A(n333), .ZN(n21978) );
  INV_X1 U15337 ( .A(n332), .ZN(n21979) );
  INV_X1 U15338 ( .A(n332), .ZN(n21980) );
  INV_X1 U15339 ( .A(n331), .ZN(n21981) );
  INV_X1 U15340 ( .A(n331), .ZN(n21982) );
  INV_X1 U15341 ( .A(n330), .ZN(n21983) );
  INV_X1 U15342 ( .A(n330), .ZN(n21984) );
  INV_X1 U15343 ( .A(n329), .ZN(n21985) );
  INV_X1 U15344 ( .A(n329), .ZN(n21986) );
  INV_X1 U15345 ( .A(n328), .ZN(n21987) );
  INV_X1 U15346 ( .A(n328), .ZN(n21988) );
  INV_X1 U15347 ( .A(n327), .ZN(n21989) );
  INV_X1 U15348 ( .A(n327), .ZN(n21990) );
  INV_X1 U15349 ( .A(n326), .ZN(n21991) );
  INV_X1 U15350 ( .A(n326), .ZN(n21992) );
  INV_X1 U15351 ( .A(n325), .ZN(n21993) );
  INV_X1 U15352 ( .A(n325), .ZN(n21994) );
  INV_X1 U15353 ( .A(n324), .ZN(n21995) );
  INV_X1 U15354 ( .A(n324), .ZN(n21996) );
  INV_X1 U15355 ( .A(n323), .ZN(n21997) );
  INV_X1 U15356 ( .A(n323), .ZN(n21998) );
  INV_X1 U15357 ( .A(n322), .ZN(n21999) );
  INV_X1 U15358 ( .A(n322), .ZN(n22000) );
  INV_X1 U15359 ( .A(n321), .ZN(n22001) );
  INV_X1 U15360 ( .A(n321), .ZN(n22002) );
  INV_X1 U15361 ( .A(n320), .ZN(n22003) );
  INV_X1 U15362 ( .A(n320), .ZN(n22004) );
  INV_X1 U15363 ( .A(n319), .ZN(n22005) );
  INV_X1 U15364 ( .A(n319), .ZN(n22006) );
  INV_X1 U15365 ( .A(n318), .ZN(n22007) );
  INV_X1 U15366 ( .A(n318), .ZN(n22008) );
  INV_X1 U15367 ( .A(n317), .ZN(n22009) );
  INV_X1 U15368 ( .A(n317), .ZN(n22010) );
  INV_X1 U15369 ( .A(n316), .ZN(n22011) );
  INV_X1 U15370 ( .A(n316), .ZN(n22012) );
  INV_X1 U15371 ( .A(n315), .ZN(n22013) );
  INV_X1 U15372 ( .A(n315), .ZN(n22014) );
  INV_X1 U15373 ( .A(n314), .ZN(n22015) );
  INV_X1 U15374 ( .A(n314), .ZN(n22016) );
  INV_X1 U15375 ( .A(n313), .ZN(n22017) );
  INV_X1 U15376 ( .A(n313), .ZN(n22018) );
  INV_X1 U15377 ( .A(n312), .ZN(n22019) );
  INV_X1 U15378 ( .A(n312), .ZN(n22020) );
  INV_X1 U15379 ( .A(n311), .ZN(n22021) );
  INV_X1 U15380 ( .A(n311), .ZN(n22022) );
  INV_X1 U15381 ( .A(n310), .ZN(n22023) );
  INV_X1 U15382 ( .A(n310), .ZN(n22024) );
  INV_X1 U15383 ( .A(n309), .ZN(n22025) );
  INV_X1 U15384 ( .A(n309), .ZN(n22026) );
  INV_X1 U15385 ( .A(n308), .ZN(n22027) );
  INV_X1 U15386 ( .A(n308), .ZN(n22028) );
  INV_X1 U15387 ( .A(n307), .ZN(n22029) );
  INV_X1 U15388 ( .A(n307), .ZN(n22030) );
  INV_X1 U15389 ( .A(n306), .ZN(n22031) );
  INV_X1 U15390 ( .A(n306), .ZN(n22032) );
  INV_X1 U15391 ( .A(n305), .ZN(n22033) );
  INV_X1 U15392 ( .A(n305), .ZN(n22034) );
  INV_X1 U15393 ( .A(n304), .ZN(n22035) );
  INV_X1 U15394 ( .A(n304), .ZN(n22036) );
  INV_X1 U15395 ( .A(n303), .ZN(n22037) );
  INV_X1 U15396 ( .A(n303), .ZN(n22038) );
  INV_X1 U15397 ( .A(n302), .ZN(n22039) );
  INV_X1 U15398 ( .A(n302), .ZN(n22040) );
  INV_X1 U15399 ( .A(n301), .ZN(n22041) );
  INV_X1 U15400 ( .A(n301), .ZN(n22042) );
  INV_X1 U15401 ( .A(n300), .ZN(n22043) );
  INV_X1 U15402 ( .A(n300), .ZN(n22044) );
  INV_X1 U15403 ( .A(n299), .ZN(n22045) );
  INV_X1 U15404 ( .A(n299), .ZN(n22046) );
  INV_X1 U15405 ( .A(n298), .ZN(n22047) );
  INV_X1 U15406 ( .A(n298), .ZN(n22048) );
  INV_X1 U15407 ( .A(n297), .ZN(n22049) );
  INV_X1 U15408 ( .A(n297), .ZN(n22050) );
  INV_X1 U15409 ( .A(n296), .ZN(n22051) );
  INV_X1 U15410 ( .A(n296), .ZN(n22052) );
  INV_X1 U15411 ( .A(n295), .ZN(n22053) );
  INV_X1 U15412 ( .A(n295), .ZN(n22054) );
  INV_X1 U15413 ( .A(n294), .ZN(n22055) );
  INV_X1 U15414 ( .A(n294), .ZN(n22056) );
  INV_X1 U15415 ( .A(n293), .ZN(n22057) );
  INV_X1 U15416 ( .A(n293), .ZN(n22058) );
  INV_X1 U15417 ( .A(n292), .ZN(n22059) );
  INV_X1 U15418 ( .A(n292), .ZN(n22060) );
  INV_X1 U15419 ( .A(n291), .ZN(n22061) );
  INV_X1 U15420 ( .A(n291), .ZN(n22062) );
  INV_X1 U15421 ( .A(n290), .ZN(n22063) );
  INV_X1 U15422 ( .A(n290), .ZN(n22064) );
  INV_X1 U15423 ( .A(n289), .ZN(n22065) );
  INV_X1 U15424 ( .A(n289), .ZN(n22066) );
  INV_X1 U15425 ( .A(n288), .ZN(n22067) );
  INV_X1 U15426 ( .A(n288), .ZN(n22068) );
  INV_X1 U15427 ( .A(n287), .ZN(n22069) );
  INV_X1 U15428 ( .A(n287), .ZN(n22070) );
  INV_X1 U15429 ( .A(n286), .ZN(n22071) );
  INV_X1 U15430 ( .A(n286), .ZN(n22072) );
  INV_X1 U15431 ( .A(n285), .ZN(n22073) );
  INV_X1 U15432 ( .A(n285), .ZN(n22074) );
  INV_X1 U15433 ( .A(n284), .ZN(n22075) );
  INV_X1 U15434 ( .A(n284), .ZN(n22076) );
  INV_X1 U15435 ( .A(n283), .ZN(n22077) );
  INV_X1 U15436 ( .A(n283), .ZN(n22078) );
  INV_X1 U15437 ( .A(n282), .ZN(n22079) );
  INV_X1 U15438 ( .A(n282), .ZN(n22080) );
  INV_X1 U15439 ( .A(n281), .ZN(n22081) );
  INV_X1 U15440 ( .A(n281), .ZN(n22082) );
  INV_X1 U15441 ( .A(n280), .ZN(n22083) );
  INV_X1 U15442 ( .A(n280), .ZN(n22084) );
  INV_X1 U15443 ( .A(n279), .ZN(n22085) );
  INV_X1 U15444 ( .A(n279), .ZN(n22086) );
  INV_X1 U15445 ( .A(n278), .ZN(n22087) );
  INV_X1 U15446 ( .A(n278), .ZN(n22088) );
  INV_X1 U15447 ( .A(n277), .ZN(n22089) );
  INV_X1 U15448 ( .A(n277), .ZN(n22090) );
  INV_X1 U15449 ( .A(n276), .ZN(n22091) );
  INV_X1 U15450 ( .A(n276), .ZN(n22092) );
  INV_X1 U15451 ( .A(n275), .ZN(n22093) );
  INV_X1 U15452 ( .A(n275), .ZN(n22094) );
  INV_X1 U15453 ( .A(n274), .ZN(n22095) );
  INV_X1 U15454 ( .A(n274), .ZN(n22096) );
  INV_X1 U15455 ( .A(n273), .ZN(n22097) );
  INV_X1 U15456 ( .A(n273), .ZN(n22098) );
  INV_X1 U15457 ( .A(n272), .ZN(n22099) );
  INV_X1 U15458 ( .A(n272), .ZN(n22100) );
  INV_X1 U15459 ( .A(n271), .ZN(n22101) );
  INV_X1 U15460 ( .A(n271), .ZN(n22102) );
  INV_X1 U15461 ( .A(n270), .ZN(n22103) );
  INV_X1 U15462 ( .A(n270), .ZN(n22104) );
  INV_X1 U15463 ( .A(n269), .ZN(n22105) );
  INV_X1 U15464 ( .A(n269), .ZN(n22106) );
  INV_X1 U15465 ( .A(n268), .ZN(n22107) );
  INV_X1 U15466 ( .A(n268), .ZN(n22108) );
  INV_X1 U15467 ( .A(n267), .ZN(n22109) );
  INV_X1 U15468 ( .A(n267), .ZN(n22110) );
  INV_X1 U15469 ( .A(n266), .ZN(n22111) );
  INV_X1 U15470 ( .A(n266), .ZN(n22112) );
  INV_X1 U15471 ( .A(n265), .ZN(n22113) );
  INV_X1 U15472 ( .A(n265), .ZN(n22114) );
  INV_X1 U15473 ( .A(n264), .ZN(n22115) );
  INV_X1 U15474 ( .A(n264), .ZN(n22116) );
  INV_X1 U15475 ( .A(n263), .ZN(n22117) );
  INV_X1 U15476 ( .A(n263), .ZN(n22118) );
  INV_X1 U15477 ( .A(n262), .ZN(n22119) );
  INV_X1 U15478 ( .A(n262), .ZN(n22120) );
  INV_X1 U15479 ( .A(n261), .ZN(n22121) );
  INV_X1 U15480 ( .A(n261), .ZN(n22122) );
  INV_X1 U15481 ( .A(n260), .ZN(n22123) );
  INV_X1 U15482 ( .A(n260), .ZN(n22124) );
  INV_X1 U15483 ( .A(n259), .ZN(n22125) );
  INV_X1 U15484 ( .A(n259), .ZN(n22126) );
  INV_X1 U15485 ( .A(n258), .ZN(n22127) );
  INV_X1 U15486 ( .A(n258), .ZN(n22128) );
  INV_X1 U15487 ( .A(n257), .ZN(n22129) );
  INV_X1 U15488 ( .A(n257), .ZN(n22130) );
  INV_X1 U15489 ( .A(n26433), .ZN(n22131) );
  INV_X1 U15490 ( .A(n22131), .ZN(n22132) );
  INV_X1 U15491 ( .A(n22131), .ZN(n22133) );
  INV_X1 U15492 ( .A(n256), .ZN(n22134) );
  INV_X1 U15493 ( .A(n256), .ZN(n22135) );
  INV_X1 U15494 ( .A(n26434), .ZN(n22136) );
  INV_X1 U15495 ( .A(n22136), .ZN(n22137) );
  INV_X1 U15496 ( .A(n22136), .ZN(n22138) );
  INV_X1 U15497 ( .A(n255), .ZN(n22139) );
  INV_X1 U15498 ( .A(n255), .ZN(n22140) );
  INV_X1 U15499 ( .A(n26432), .ZN(n22141) );
  INV_X1 U15500 ( .A(n22141), .ZN(n22142) );
  INV_X1 U15501 ( .A(n22141), .ZN(n22143) );
  INV_X1 U15502 ( .A(n254), .ZN(n22144) );
  INV_X1 U15503 ( .A(n254), .ZN(n22145) );
  INV_X1 U15504 ( .A(n253), .ZN(n22146) );
  INV_X1 U15505 ( .A(n253), .ZN(n22147) );
  INV_X1 U15506 ( .A(n26432), .ZN(n22148) );
  INV_X1 U15507 ( .A(n22148), .ZN(n22149) );
  INV_X1 U15508 ( .A(n22148), .ZN(n22150) );
  INV_X1 U15509 ( .A(n26433), .ZN(n22151) );
  INV_X1 U15510 ( .A(n22151), .ZN(n22152) );
  INV_X1 U15511 ( .A(n22151), .ZN(n22153) );
  INV_X1 U15512 ( .A(n26434), .ZN(n22154) );
  INV_X1 U15513 ( .A(n22154), .ZN(n22155) );
  INV_X1 U15514 ( .A(n22154), .ZN(n22156) );
  INV_X1 U15515 ( .A(n252), .ZN(n22157) );
  INV_X1 U15516 ( .A(n252), .ZN(n22158) );
  INV_X1 U15517 ( .A(n26438), .ZN(n22159) );
  INV_X1 U15518 ( .A(n22159), .ZN(n22160) );
  INV_X1 U15519 ( .A(n22159), .ZN(n22161) );
  INV_X1 U15520 ( .A(n251), .ZN(n22162) );
  INV_X1 U15521 ( .A(n251), .ZN(n22163) );
  INV_X1 U15522 ( .A(n250), .ZN(n22164) );
  INV_X1 U15523 ( .A(n250), .ZN(n22165) );
  INV_X1 U15524 ( .A(n264401), .ZN(n22166) );
  INV_X1 U15525 ( .A(n22166), .ZN(n22167) );
  INV_X1 U15526 ( .A(n22166), .ZN(n22168) );
  INV_X1 U15527 ( .A(n249), .ZN(n22169) );
  INV_X1 U15528 ( .A(n249), .ZN(n22170) );
  INV_X1 U15529 ( .A(n248), .ZN(n22171) );
  INV_X1 U15530 ( .A(n248), .ZN(n22172) );
  INV_X1 U15531 ( .A(n247), .ZN(n22173) );
  INV_X1 U15532 ( .A(n247), .ZN(n22174) );
  INV_X1 U15533 ( .A(n26439), .ZN(n22175) );
  INV_X1 U15534 ( .A(n22175), .ZN(n22176) );
  INV_X1 U15535 ( .A(n22175), .ZN(n22177) );
  INV_X1 U15536 ( .A(n26438), .ZN(n22178) );
  INV_X1 U15537 ( .A(n22178), .ZN(n22179) );
  INV_X1 U15538 ( .A(n22178), .ZN(n22180) );
  INV_X1 U15539 ( .A(n26439), .ZN(n22181) );
  INV_X1 U15540 ( .A(n22181), .ZN(n22182) );
  INV_X1 U15541 ( .A(n22181), .ZN(n22183) );
  INV_X1 U15542 ( .A(n264401), .ZN(n22184) );
  INV_X1 U15543 ( .A(n22184), .ZN(n22185) );
  INV_X1 U15544 ( .A(n22184), .ZN(n22186) );
  INV_X1 U15545 ( .A(n26444), .ZN(n22187) );
  INV_X1 U15546 ( .A(n22187), .ZN(n22188) );
  INV_X1 U15547 ( .A(n22187), .ZN(n22189) );
  INV_X1 U15548 ( .A(n246), .ZN(n22190) );
  INV_X1 U15549 ( .A(n246), .ZN(n22191) );
  INV_X1 U15550 ( .A(n245), .ZN(n22192) );
  INV_X1 U15551 ( .A(n245), .ZN(n22193) );
  INV_X1 U15552 ( .A(n244), .ZN(n22194) );
  INV_X1 U15553 ( .A(n244), .ZN(n22195) );
  INV_X1 U15554 ( .A(n26442), .ZN(n22196) );
  INV_X1 U15555 ( .A(n22196), .ZN(n22197) );
  INV_X1 U15556 ( .A(n22196), .ZN(n22198) );
  INV_X1 U15557 ( .A(n26443), .ZN(n22199) );
  INV_X1 U15558 ( .A(n22199), .ZN(n22200) );
  INV_X1 U15559 ( .A(n22199), .ZN(n22201) );
  INV_X1 U15560 ( .A(n26442), .ZN(n22202) );
  INV_X1 U15561 ( .A(n22202), .ZN(n22203) );
  INV_X1 U15562 ( .A(n22202), .ZN(n22204) );
  INV_X1 U15563 ( .A(n26443), .ZN(n22205) );
  INV_X1 U15564 ( .A(n22205), .ZN(n22206) );
  INV_X1 U15565 ( .A(n22205), .ZN(n22207) );
  INV_X1 U15566 ( .A(n26444), .ZN(n22208) );
  INV_X1 U15567 ( .A(n22208), .ZN(n22209) );
  INV_X1 U15568 ( .A(n22208), .ZN(n22210) );
  INV_X1 U15569 ( .A(n243), .ZN(n22211) );
  INV_X1 U15570 ( .A(n243), .ZN(n22212) );
  INV_X1 U15571 ( .A(n242), .ZN(n22213) );
  INV_X1 U15572 ( .A(n242), .ZN(n22214) );
  INV_X1 U15573 ( .A(n241), .ZN(n22215) );
  INV_X1 U15574 ( .A(n241), .ZN(n22216) );
  INV_X1 U15575 ( .A(n240), .ZN(n22217) );
  INV_X1 U15576 ( .A(n240), .ZN(n22218) );
  INV_X1 U15577 ( .A(n239), .ZN(n22219) );
  INV_X1 U15578 ( .A(n239), .ZN(n22220) );
  INV_X1 U15579 ( .A(n238), .ZN(n22221) );
  INV_X1 U15580 ( .A(n238), .ZN(n22222) );
  INV_X1 U15581 ( .A(n237), .ZN(n22223) );
  INV_X1 U15582 ( .A(n237), .ZN(n22224) );
  INV_X1 U15583 ( .A(n236), .ZN(n22225) );
  INV_X1 U15584 ( .A(n236), .ZN(n22226) );
  INV_X1 U15585 ( .A(n235), .ZN(n22227) );
  INV_X1 U15586 ( .A(n235), .ZN(n22228) );
  INV_X1 U15587 ( .A(n234), .ZN(n22229) );
  INV_X1 U15588 ( .A(n234), .ZN(n22230) );
  INV_X1 U15589 ( .A(n233), .ZN(n22231) );
  INV_X1 U15590 ( .A(n233), .ZN(n22232) );
  INV_X1 U15591 ( .A(n232), .ZN(n22233) );
  INV_X1 U15592 ( .A(n232), .ZN(n22234) );
  INV_X1 U15593 ( .A(n231), .ZN(n22235) );
  INV_X1 U15594 ( .A(n231), .ZN(n22236) );
  INV_X1 U15595 ( .A(n230), .ZN(n22237) );
  INV_X1 U15596 ( .A(n230), .ZN(n22238) );
  INV_X1 U15597 ( .A(n229), .ZN(n22239) );
  INV_X1 U15598 ( .A(n229), .ZN(n22240) );
  INV_X1 U15599 ( .A(n228), .ZN(n22241) );
  INV_X1 U15600 ( .A(n228), .ZN(n22242) );
  INV_X1 U15601 ( .A(n227), .ZN(n22243) );
  INV_X1 U15602 ( .A(n227), .ZN(n22244) );
  INV_X1 U15603 ( .A(n226), .ZN(n22245) );
  INV_X1 U15604 ( .A(n226), .ZN(n22246) );
  INV_X1 U15605 ( .A(n225), .ZN(n22247) );
  INV_X1 U15606 ( .A(n225), .ZN(n22248) );
  INV_X1 U15607 ( .A(n224), .ZN(n22249) );
  INV_X1 U15608 ( .A(n224), .ZN(n22250) );
  INV_X1 U15609 ( .A(n223), .ZN(n22251) );
  INV_X1 U15610 ( .A(n223), .ZN(n22252) );
  INV_X1 U15611 ( .A(n222), .ZN(n22253) );
  INV_X1 U15612 ( .A(n222), .ZN(n22254) );
  INV_X1 U15613 ( .A(n221), .ZN(n22255) );
  INV_X1 U15614 ( .A(n220), .ZN(n22256) );
  INV_X1 U15615 ( .A(n220), .ZN(n22257) );
  INV_X1 U15616 ( .A(n219), .ZN(n22258) );
  INV_X1 U15617 ( .A(n219), .ZN(n22259) );
  INV_X1 U15618 ( .A(n218), .ZN(n22260) );
  INV_X1 U15619 ( .A(n218), .ZN(n22261) );
  INV_X1 U15620 ( .A(n217), .ZN(n22262) );
  INV_X1 U15621 ( .A(n217), .ZN(n22263) );
  INV_X1 U15622 ( .A(n27124), .ZN(n22264) );
  INV_X1 U15623 ( .A(n22264), .ZN(n22265) );
  INV_X1 U15624 ( .A(n22264), .ZN(n22266) );
  INV_X1 U15625 ( .A(n23587), .ZN(n22267) );
  INV_X1 U15626 ( .A(n23587), .ZN(n22268) );
  INV_X1 U15627 ( .A(n26829), .ZN(n22269) );
  INV_X1 U15628 ( .A(n22269), .ZN(n22270) );
  INV_X1 U15629 ( .A(n22269), .ZN(n22271) );
  INV_X1 U15630 ( .A(n22271), .ZN(n22272) );
  INV_X1 U15631 ( .A(n22272), .ZN(n22273) );
  INV_X1 U15632 ( .A(n22272), .ZN(n22274) );
  INV_X1 U15633 ( .A(n216), .ZN(n22275) );
  INV_X1 U15634 ( .A(n216), .ZN(n22276) );
  INV_X1 U15635 ( .A(n18861), .ZN(n22277) );
  INV_X1 U15636 ( .A(n22277), .ZN(n22278) );
  INV_X1 U15637 ( .A(n22277), .ZN(n22279) );
  INV_X1 U15638 ( .A(n26855), .ZN(n22280) );
  INV_X1 U15639 ( .A(n22280), .ZN(n22281) );
  INV_X1 U15640 ( .A(n22280), .ZN(n22282) );
  INV_X1 U15641 ( .A(n18439), .ZN(n22283) );
  INV_X1 U15642 ( .A(n18439), .ZN(n22284) );
  INV_X1 U15643 ( .A(n26456), .ZN(n22285) );
  INV_X1 U15644 ( .A(n22285), .ZN(n22286) );
  INV_X1 U15645 ( .A(n22285), .ZN(n22287) );
  INV_X1 U15646 ( .A(n18440), .ZN(n22288) );
  INV_X1 U15647 ( .A(n18440), .ZN(n22289) );
  INV_X1 U15648 ( .A(n26459), .ZN(n22290) );
  INV_X1 U15649 ( .A(n22290), .ZN(n22291) );
  INV_X1 U15650 ( .A(n22290), .ZN(n22292) );
  INV_X1 U15651 ( .A(n18441), .ZN(n22293) );
  INV_X1 U15652 ( .A(n18441), .ZN(n22294) );
  INV_X1 U15653 ( .A(n26462), .ZN(n22295) );
  INV_X1 U15654 ( .A(n22295), .ZN(n22296) );
  INV_X1 U15655 ( .A(n22295), .ZN(n22297) );
  INV_X1 U15656 ( .A(n18442), .ZN(n22298) );
  INV_X1 U15657 ( .A(n18442), .ZN(n22299) );
  INV_X1 U15658 ( .A(n26465), .ZN(n22300) );
  INV_X1 U15659 ( .A(n22300), .ZN(n22301) );
  INV_X1 U15660 ( .A(n22300), .ZN(n22302) );
  INV_X1 U15661 ( .A(n18443), .ZN(n22303) );
  INV_X1 U15662 ( .A(n18443), .ZN(n22304) );
  INV_X1 U15663 ( .A(n26468), .ZN(n22305) );
  INV_X1 U15664 ( .A(n22305), .ZN(n22306) );
  INV_X1 U15665 ( .A(n22305), .ZN(n22307) );
  INV_X1 U15666 ( .A(n18444), .ZN(n22308) );
  INV_X1 U15667 ( .A(n18444), .ZN(n22309) );
  INV_X1 U15668 ( .A(n26472), .ZN(n22310) );
  INV_X1 U15669 ( .A(n22310), .ZN(n22311) );
  INV_X1 U15670 ( .A(n22310), .ZN(n22312) );
  INV_X1 U15671 ( .A(n18445), .ZN(n22313) );
  INV_X1 U15672 ( .A(n18445), .ZN(n22314) );
  INV_X1 U15673 ( .A(n26474), .ZN(n22315) );
  INV_X1 U15674 ( .A(n22315), .ZN(n22316) );
  INV_X1 U15675 ( .A(n22315), .ZN(n22317) );
  INV_X1 U15676 ( .A(n18446), .ZN(n22318) );
  INV_X1 U15677 ( .A(n18446), .ZN(n22319) );
  INV_X1 U15678 ( .A(n26477), .ZN(n22320) );
  INV_X1 U15679 ( .A(n22320), .ZN(n22321) );
  INV_X1 U15680 ( .A(n22320), .ZN(n22322) );
  INV_X1 U15681 ( .A(n215), .ZN(n22323) );
  INV_X1 U15682 ( .A(n215), .ZN(n22324) );
  INV_X1 U15683 ( .A(n214), .ZN(n22325) );
  INV_X1 U15684 ( .A(n214), .ZN(n22326) );
  INV_X1 U15685 ( .A(n213), .ZN(n22327) );
  INV_X1 U15686 ( .A(n213), .ZN(n22328) );
  INV_X1 U15687 ( .A(n212), .ZN(n22329) );
  INV_X1 U15688 ( .A(n212), .ZN(n22330) );
  INV_X1 U15689 ( .A(n211), .ZN(n22331) );
  INV_X1 U15690 ( .A(n211), .ZN(n22332) );
  INV_X1 U15691 ( .A(n210), .ZN(n22333) );
  INV_X1 U15692 ( .A(n210), .ZN(n22334) );
  INV_X1 U15693 ( .A(n209), .ZN(n22335) );
  INV_X1 U15694 ( .A(n209), .ZN(n22336) );
  INV_X1 U15695 ( .A(n208), .ZN(n22337) );
  INV_X1 U15696 ( .A(n208), .ZN(n22338) );
  INV_X1 U15697 ( .A(n207), .ZN(n22339) );
  INV_X1 U15698 ( .A(n207), .ZN(n22340) );
  INV_X1 U15699 ( .A(n206), .ZN(n22341) );
  INV_X1 U15700 ( .A(n206), .ZN(n22342) );
  INV_X1 U15701 ( .A(n205), .ZN(n22343) );
  INV_X1 U15702 ( .A(n205), .ZN(n22344) );
  INV_X1 U15703 ( .A(n204), .ZN(n22345) );
  INV_X1 U15704 ( .A(n204), .ZN(n22346) );
  INV_X1 U15705 ( .A(n203), .ZN(n22347) );
  INV_X1 U15706 ( .A(n203), .ZN(n22348) );
  INV_X1 U15707 ( .A(n202), .ZN(n22349) );
  INV_X1 U15708 ( .A(n202), .ZN(n22350) );
  INV_X1 U15709 ( .A(n201), .ZN(n22351) );
  INV_X1 U15710 ( .A(n201), .ZN(n22352) );
  INV_X1 U15711 ( .A(n200), .ZN(n22353) );
  INV_X1 U15712 ( .A(n200), .ZN(n22354) );
  INV_X1 U15713 ( .A(n199), .ZN(n22355) );
  INV_X1 U15714 ( .A(n199), .ZN(n22356) );
  INV_X1 U15715 ( .A(n198), .ZN(n22357) );
  INV_X1 U15716 ( .A(n198), .ZN(n22358) );
  INV_X1 U15717 ( .A(n197), .ZN(n22359) );
  INV_X1 U15718 ( .A(n197), .ZN(n22360) );
  INV_X1 U15719 ( .A(n196), .ZN(n22361) );
  INV_X1 U15720 ( .A(n196), .ZN(n22362) );
  INV_X1 U15721 ( .A(n195), .ZN(n22363) );
  INV_X1 U15722 ( .A(n195), .ZN(n22364) );
  INV_X1 U15723 ( .A(n194), .ZN(n22365) );
  INV_X1 U15724 ( .A(n194), .ZN(n22366) );
  INV_X1 U15725 ( .A(n193), .ZN(n22367) );
  INV_X1 U15726 ( .A(n193), .ZN(n22368) );
  INV_X1 U15727 ( .A(n192), .ZN(n22369) );
  INV_X1 U15728 ( .A(n192), .ZN(n22370) );
  INV_X1 U15729 ( .A(n191), .ZN(n22371) );
  INV_X1 U15730 ( .A(n191), .ZN(n22372) );
  INV_X1 U15731 ( .A(n190), .ZN(n22373) );
  INV_X1 U15732 ( .A(n190), .ZN(n22374) );
  INV_X1 U15733 ( .A(n189), .ZN(n22375) );
  INV_X1 U15734 ( .A(n189), .ZN(n22376) );
  INV_X1 U15735 ( .A(n188), .ZN(n22377) );
  INV_X1 U15736 ( .A(n188), .ZN(n22378) );
  INV_X1 U15737 ( .A(n187), .ZN(n22379) );
  INV_X1 U15738 ( .A(n187), .ZN(n22380) );
  INV_X1 U15739 ( .A(n186), .ZN(n22381) );
  INV_X1 U15740 ( .A(n186), .ZN(n22382) );
  INV_X1 U15741 ( .A(n185), .ZN(n22383) );
  INV_X1 U15742 ( .A(n185), .ZN(n22384) );
  INV_X1 U15743 ( .A(n184), .ZN(n22385) );
  INV_X1 U15744 ( .A(n184), .ZN(n22386) );
  INV_X1 U15745 ( .A(n183), .ZN(n22387) );
  INV_X1 U15746 ( .A(n183), .ZN(n22388) );
  INV_X1 U15747 ( .A(n182), .ZN(n22389) );
  INV_X1 U15748 ( .A(n182), .ZN(n22390) );
  INV_X1 U15749 ( .A(n181), .ZN(n22391) );
  INV_X1 U15750 ( .A(n181), .ZN(n22392) );
  INV_X1 U15751 ( .A(n180), .ZN(n22393) );
  INV_X1 U15752 ( .A(n180), .ZN(n22394) );
  INV_X1 U15753 ( .A(n179), .ZN(n22395) );
  INV_X1 U15754 ( .A(n179), .ZN(n22396) );
  INV_X1 U15755 ( .A(n178), .ZN(n22397) );
  INV_X1 U15756 ( .A(n178), .ZN(n22398) );
  INV_X1 U15757 ( .A(n177), .ZN(n22399) );
  INV_X1 U15758 ( .A(n177), .ZN(n22400) );
  INV_X1 U15759 ( .A(n176), .ZN(n22401) );
  INV_X1 U15760 ( .A(n176), .ZN(n22402) );
  INV_X1 U15761 ( .A(n175), .ZN(n22403) );
  INV_X1 U15762 ( .A(n175), .ZN(n22404) );
  INV_X1 U15763 ( .A(n174), .ZN(n22405) );
  INV_X1 U15764 ( .A(n174), .ZN(n22406) );
  INV_X1 U15765 ( .A(n173), .ZN(n22407) );
  INV_X1 U15766 ( .A(n173), .ZN(n22408) );
  INV_X1 U15767 ( .A(n172), .ZN(n22409) );
  INV_X1 U15768 ( .A(n172), .ZN(n22410) );
  INV_X1 U15769 ( .A(n171), .ZN(n22411) );
  INV_X1 U15770 ( .A(n171), .ZN(n22412) );
  INV_X1 U15771 ( .A(n170), .ZN(n22413) );
  INV_X1 U15772 ( .A(n170), .ZN(n22414) );
  INV_X1 U15773 ( .A(n169), .ZN(n22415) );
  INV_X1 U15774 ( .A(n169), .ZN(n22416) );
  INV_X1 U15775 ( .A(n168), .ZN(n22417) );
  INV_X1 U15776 ( .A(n168), .ZN(n22418) );
  INV_X1 U15777 ( .A(n23642), .ZN(n22419) );
  INV_X1 U15778 ( .A(n23638), .ZN(n22420) );
  INV_X1 U15779 ( .A(n18447), .ZN(n22421) );
  INV_X1 U15780 ( .A(n18447), .ZN(n22422) );
  INV_X1 U15781 ( .A(n265001), .ZN(n22423) );
  INV_X1 U15782 ( .A(n22423), .ZN(n22424) );
  INV_X1 U15783 ( .A(n22423), .ZN(n22425) );
  INV_X1 U15784 ( .A(n24876), .ZN(n22426) );
  INV_X1 U15785 ( .A(n22426), .ZN(n22427) );
  INV_X1 U15786 ( .A(n22426), .ZN(n22428) );
  INV_X1 U15787 ( .A(n26503), .ZN(n22429) );
  INV_X1 U15788 ( .A(n22429), .ZN(n22430) );
  INV_X1 U15789 ( .A(n22429), .ZN(n22431) );
  INV_X1 U15790 ( .A(n18448), .ZN(n22432) );
  INV_X1 U15791 ( .A(n18448), .ZN(n22433) );
  INV_X1 U15792 ( .A(n17115), .ZN(n22434) );
  INV_X1 U15793 ( .A(n17115), .ZN(n22435) );
  INV_X1 U15794 ( .A(n18449), .ZN(n22436) );
  INV_X1 U15795 ( .A(n18449), .ZN(n22437) );
  INV_X1 U15796 ( .A(n26507), .ZN(n22438) );
  INV_X1 U15797 ( .A(n22438), .ZN(n22439) );
  INV_X1 U15798 ( .A(n22438), .ZN(n22440) );
  INV_X1 U15799 ( .A(n18450), .ZN(n22441) );
  INV_X1 U15800 ( .A(n18450), .ZN(n22442) );
  INV_X1 U15801 ( .A(n26511), .ZN(n22443) );
  INV_X1 U15802 ( .A(n22443), .ZN(n22444) );
  INV_X1 U15803 ( .A(n22443), .ZN(n22445) );
  INV_X1 U15804 ( .A(n21867), .ZN(n22446) );
  INV_X1 U15805 ( .A(n22446), .ZN(n22447) );
  INV_X1 U15806 ( .A(n22446), .ZN(n22448) );
  INV_X1 U15807 ( .A(n26516), .ZN(n22449) );
  INV_X1 U15808 ( .A(n22449), .ZN(n22450) );
  INV_X1 U15809 ( .A(n22449), .ZN(n22451) );
  INV_X1 U15810 ( .A(n26518), .ZN(n22452) );
  INV_X1 U15811 ( .A(n22452), .ZN(n22453) );
  INV_X1 U15812 ( .A(n22452), .ZN(n22454) );
  INV_X1 U15813 ( .A(n26521), .ZN(n22455) );
  INV_X1 U15814 ( .A(n22455), .ZN(n22456) );
  INV_X1 U15815 ( .A(n22455), .ZN(n22457) );
  INV_X1 U15816 ( .A(n26523), .ZN(n22458) );
  INV_X1 U15817 ( .A(n22458), .ZN(n22459) );
  INV_X1 U15818 ( .A(n22458), .ZN(n22460) );
  INV_X1 U15819 ( .A(n26993), .ZN(n22461) );
  INV_X1 U15820 ( .A(n22461), .ZN(n22462) );
  INV_X1 U15821 ( .A(n22461), .ZN(n22463) );
  INV_X1 U15822 ( .A(n26994), .ZN(n22464) );
  INV_X1 U15823 ( .A(n22464), .ZN(n22465) );
  INV_X1 U15824 ( .A(n22464), .ZN(n22466) );
  INV_X1 U15825 ( .A(n26529), .ZN(n22467) );
  INV_X1 U15826 ( .A(n22467), .ZN(n22468) );
  INV_X1 U15827 ( .A(n22467), .ZN(n22469) );
  INV_X1 U15828 ( .A(n26527), .ZN(n22470) );
  INV_X1 U15829 ( .A(n22470), .ZN(n22471) );
  INV_X1 U15830 ( .A(n22470), .ZN(n22472) );
  INV_X1 U15831 ( .A(n26532), .ZN(n22473) );
  INV_X1 U15832 ( .A(n22473), .ZN(n22474) );
  INV_X1 U15833 ( .A(n22473), .ZN(n22475) );
  INV_X1 U15834 ( .A(n26534), .ZN(n22476) );
  INV_X1 U15835 ( .A(n22476), .ZN(n22477) );
  INV_X1 U15836 ( .A(n22476), .ZN(n22478) );
  INV_X1 U15837 ( .A(n26536), .ZN(n22479) );
  INV_X1 U15838 ( .A(n22479), .ZN(n22480) );
  INV_X1 U15839 ( .A(n22479), .ZN(n22481) );
  INV_X1 U15840 ( .A(n26102), .ZN(n22482) );
  INV_X1 U15841 ( .A(n22482), .ZN(n22483) );
  INV_X1 U15842 ( .A(n22482), .ZN(n22484) );
  INV_X1 U15843 ( .A(n26538), .ZN(n22485) );
  INV_X1 U15844 ( .A(n22485), .ZN(n22486) );
  INV_X1 U15845 ( .A(n22485), .ZN(n22487) );
  INV_X1 U15846 ( .A(n26091), .ZN(n22488) );
  INV_X1 U15847 ( .A(n22488), .ZN(n22489) );
  INV_X1 U15848 ( .A(n22488), .ZN(n22490) );
  INV_X1 U15849 ( .A(n27203), .ZN(n22491) );
  INV_X1 U15850 ( .A(n22491), .ZN(n22492) );
  INV_X1 U15851 ( .A(n22491), .ZN(n22493) );
  INV_X1 U15852 ( .A(n26542), .ZN(n22494) );
  INV_X1 U15853 ( .A(n22494), .ZN(n22495) );
  INV_X1 U15854 ( .A(n22494), .ZN(n22496) );
  INV_X1 U15855 ( .A(n26543), .ZN(n22497) );
  INV_X1 U15856 ( .A(n22497), .ZN(n22498) );
  INV_X1 U15857 ( .A(n22497), .ZN(n22499) );
  INV_X1 U15858 ( .A(n18451), .ZN(n22500) );
  INV_X1 U15859 ( .A(n18451), .ZN(n22501) );
  INV_X1 U15860 ( .A(n26551), .ZN(n22502) );
  INV_X1 U15861 ( .A(n22502), .ZN(n22503) );
  INV_X1 U15862 ( .A(n22502), .ZN(n22504) );
  INV_X1 U15863 ( .A(n26555), .ZN(n22505) );
  INV_X1 U15864 ( .A(n22505), .ZN(n22506) );
  INV_X1 U15865 ( .A(n22505), .ZN(n22507) );
  INV_X1 U15866 ( .A(n26554), .ZN(n22508) );
  INV_X1 U15867 ( .A(n22508), .ZN(n22509) );
  INV_X1 U15868 ( .A(n22508), .ZN(n22510) );
  INV_X1 U15869 ( .A(n26557), .ZN(n22511) );
  INV_X1 U15870 ( .A(n22511), .ZN(n22512) );
  INV_X1 U15871 ( .A(n22511), .ZN(n22513) );
  INV_X1 U15872 ( .A(n26563), .ZN(n22514) );
  INV_X1 U15873 ( .A(n22514), .ZN(n22515) );
  INV_X1 U15874 ( .A(n22514), .ZN(n22516) );
  INV_X1 U15875 ( .A(n26567), .ZN(n22517) );
  INV_X1 U15876 ( .A(n22517), .ZN(n22518) );
  INV_X1 U15877 ( .A(n22517), .ZN(n22519) );
  INV_X1 U15878 ( .A(n26571), .ZN(n22520) );
  INV_X1 U15879 ( .A(n22520), .ZN(n22521) );
  INV_X1 U15880 ( .A(n22520), .ZN(n22522) );
  INV_X1 U15881 ( .A(n26576), .ZN(n22523) );
  INV_X1 U15882 ( .A(n22523), .ZN(n22524) );
  INV_X1 U15883 ( .A(n22523), .ZN(n22525) );
  INV_X1 U15884 ( .A(n26580), .ZN(n22526) );
  INV_X1 U15885 ( .A(n22526), .ZN(n22527) );
  INV_X1 U15886 ( .A(n22526), .ZN(n22528) );
  INV_X1 U15887 ( .A(n269401), .ZN(n22529) );
  INV_X1 U15888 ( .A(n22529), .ZN(n22530) );
  INV_X1 U15889 ( .A(n22529), .ZN(n22531) );
  INV_X1 U15890 ( .A(n26587), .ZN(n22532) );
  INV_X1 U15891 ( .A(n22532), .ZN(n22533) );
  INV_X1 U15892 ( .A(n22532), .ZN(n22534) );
  INV_X1 U15893 ( .A(n18452), .ZN(n22535) );
  INV_X1 U15894 ( .A(n18452), .ZN(n22536) );
  INV_X1 U15895 ( .A(n26592), .ZN(n22537) );
  INV_X1 U15896 ( .A(n22537), .ZN(n22538) );
  INV_X1 U15897 ( .A(n22537), .ZN(n22539) );
  INV_X1 U15898 ( .A(r899_B_2_), .ZN(n22540) );
  INV_X1 U15899 ( .A(n22540), .ZN(n22541) );
  INV_X1 U15900 ( .A(n22540), .ZN(n22542) );
  INV_X1 U15901 ( .A(n18721), .ZN(n22543) );
  INV_X1 U15902 ( .A(n22543), .ZN(n22544) );
  INV_X1 U15903 ( .A(n22543), .ZN(n22545) );
  INV_X1 U15904 ( .A(n167), .ZN(n22546) );
  INV_X1 U15905 ( .A(n167), .ZN(n22547) );
  INV_X1 U15906 ( .A(n166), .ZN(n22548) );
  INV_X1 U15907 ( .A(n166), .ZN(n22549) );
  INV_X1 U15908 ( .A(n165), .ZN(n22550) );
  INV_X1 U15909 ( .A(n165), .ZN(n22551) );
  INV_X1 U15910 ( .A(n164), .ZN(n22552) );
  INV_X1 U15911 ( .A(n164), .ZN(n22553) );
  INV_X1 U15912 ( .A(n163), .ZN(n22554) );
  INV_X1 U15913 ( .A(n163), .ZN(n22555) );
  INV_X1 U15914 ( .A(n162), .ZN(n22556) );
  INV_X1 U15915 ( .A(n162), .ZN(n22557) );
  INV_X1 U15916 ( .A(n161), .ZN(n22558) );
  INV_X1 U15917 ( .A(n161), .ZN(n22559) );
  INV_X1 U15918 ( .A(n160), .ZN(n22560) );
  INV_X1 U15919 ( .A(n160), .ZN(n22561) );
  INV_X1 U15920 ( .A(n159), .ZN(n22562) );
  INV_X1 U15921 ( .A(n159), .ZN(n22563) );
  INV_X1 U15922 ( .A(n158), .ZN(n22564) );
  INV_X1 U15923 ( .A(n158), .ZN(n22565) );
  INV_X1 U15924 ( .A(n157), .ZN(n22566) );
  INV_X1 U15925 ( .A(n157), .ZN(n22567) );
  INV_X1 U15926 ( .A(n156), .ZN(n22568) );
  INV_X1 U15927 ( .A(n156), .ZN(n22569) );
  INV_X1 U15928 ( .A(n155), .ZN(n22570) );
  INV_X1 U15929 ( .A(n155), .ZN(n22571) );
  INV_X1 U15930 ( .A(n154), .ZN(n22572) );
  INV_X1 U15931 ( .A(n154), .ZN(n22573) );
  INV_X1 U15932 ( .A(n153), .ZN(n22574) );
  INV_X1 U15933 ( .A(n153), .ZN(n22575) );
  INV_X1 U15934 ( .A(n152), .ZN(n22576) );
  INV_X1 U15935 ( .A(n152), .ZN(n22577) );
  INV_X1 U15936 ( .A(n151), .ZN(n22578) );
  INV_X1 U15937 ( .A(n151), .ZN(n22579) );
  INV_X1 U15938 ( .A(n150), .ZN(n22580) );
  INV_X1 U15939 ( .A(n150), .ZN(n22581) );
  INV_X1 U15940 ( .A(n149), .ZN(n22582) );
  INV_X1 U15941 ( .A(n149), .ZN(n22583) );
  INV_X1 U15942 ( .A(n148), .ZN(n22584) );
  INV_X1 U15943 ( .A(n148), .ZN(n22585) );
  INV_X1 U15944 ( .A(n147), .ZN(n22586) );
  INV_X1 U15945 ( .A(n147), .ZN(n22587) );
  INV_X1 U15946 ( .A(n146), .ZN(n22588) );
  INV_X1 U15947 ( .A(n146), .ZN(n22589) );
  INV_X1 U15948 ( .A(n145), .ZN(n22590) );
  INV_X1 U15949 ( .A(n145), .ZN(n22591) );
  INV_X1 U15950 ( .A(n144), .ZN(n22592) );
  INV_X1 U15951 ( .A(n144), .ZN(n22593) );
  INV_X1 U15952 ( .A(n143), .ZN(n22594) );
  INV_X1 U15953 ( .A(n143), .ZN(n22595) );
  INV_X1 U15954 ( .A(n142), .ZN(n22596) );
  INV_X1 U15955 ( .A(n142), .ZN(n22597) );
  INV_X1 U15956 ( .A(n141), .ZN(n22598) );
  INV_X1 U15957 ( .A(n141), .ZN(n22599) );
  INV_X1 U15958 ( .A(n140), .ZN(n22600) );
  INV_X1 U15959 ( .A(n140), .ZN(n22601) );
  INV_X1 U15960 ( .A(n139), .ZN(n22602) );
  INV_X1 U15961 ( .A(n139), .ZN(n22603) );
  INV_X1 U15962 ( .A(n138), .ZN(n22604) );
  INV_X1 U15963 ( .A(n138), .ZN(n22605) );
  INV_X1 U15964 ( .A(n137), .ZN(n22606) );
  INV_X1 U15965 ( .A(n137), .ZN(n22607) );
  INV_X1 U15966 ( .A(n136), .ZN(n22608) );
  INV_X1 U15967 ( .A(n136), .ZN(n22609) );
  INV_X1 U15968 ( .A(n135), .ZN(n22610) );
  INV_X1 U15969 ( .A(n135), .ZN(n22611) );
  INV_X1 U15970 ( .A(n134), .ZN(n22612) );
  INV_X1 U15971 ( .A(n134), .ZN(n22613) );
  INV_X1 U15972 ( .A(n133), .ZN(n22614) );
  INV_X1 U15973 ( .A(n133), .ZN(n22615) );
  INV_X1 U15974 ( .A(n132), .ZN(n22616) );
  INV_X1 U15975 ( .A(n132), .ZN(n22617) );
  INV_X1 U15976 ( .A(n131), .ZN(n22618) );
  INV_X1 U15977 ( .A(n131), .ZN(n22619) );
  INV_X1 U15978 ( .A(n130), .ZN(n22620) );
  INV_X1 U15979 ( .A(n130), .ZN(n22621) );
  INV_X1 U15980 ( .A(n129), .ZN(n22622) );
  INV_X1 U15981 ( .A(n129), .ZN(n22623) );
  INV_X1 U15982 ( .A(n128), .ZN(n22624) );
  INV_X1 U15983 ( .A(n128), .ZN(n22625) );
  INV_X1 U15984 ( .A(n127), .ZN(n22626) );
  INV_X1 U15985 ( .A(n127), .ZN(n22627) );
  INV_X1 U15986 ( .A(n126), .ZN(n22628) );
  INV_X1 U15987 ( .A(n126), .ZN(n22629) );
  INV_X1 U15988 ( .A(n125), .ZN(n22630) );
  INV_X1 U15989 ( .A(n125), .ZN(n22631) );
  INV_X1 U15990 ( .A(n124), .ZN(n22632) );
  INV_X1 U15991 ( .A(n124), .ZN(n22633) );
  INV_X1 U15992 ( .A(n123), .ZN(n22634) );
  INV_X1 U15993 ( .A(n123), .ZN(n22635) );
  INV_X1 U15994 ( .A(n122), .ZN(n22636) );
  INV_X1 U15995 ( .A(n122), .ZN(n22637) );
  INV_X1 U15996 ( .A(n121), .ZN(n22638) );
  INV_X1 U15997 ( .A(n121), .ZN(n22639) );
  INV_X1 U15998 ( .A(n120), .ZN(n22640) );
  INV_X1 U15999 ( .A(n120), .ZN(n22641) );
  INV_X1 U16000 ( .A(n119), .ZN(n22642) );
  INV_X1 U16001 ( .A(n119), .ZN(n22643) );
  INV_X1 U16002 ( .A(n118), .ZN(n22644) );
  INV_X1 U16003 ( .A(n118), .ZN(n22645) );
  INV_X1 U16004 ( .A(n117), .ZN(n22646) );
  INV_X1 U16005 ( .A(n117), .ZN(n22647) );
  INV_X1 U16006 ( .A(n116), .ZN(n22648) );
  INV_X1 U16007 ( .A(n116), .ZN(n22649) );
  INV_X1 U16008 ( .A(n115), .ZN(n22650) );
  INV_X1 U16009 ( .A(n115), .ZN(n22651) );
  INV_X1 U16010 ( .A(n114), .ZN(n22652) );
  INV_X1 U16011 ( .A(n114), .ZN(n22653) );
  INV_X1 U16012 ( .A(n113), .ZN(n22654) );
  INV_X1 U16013 ( .A(n113), .ZN(n22655) );
  INV_X1 U16014 ( .A(n112), .ZN(n22656) );
  INV_X1 U16015 ( .A(n112), .ZN(n22657) );
  INV_X1 U16016 ( .A(n111), .ZN(n22658) );
  INV_X1 U16017 ( .A(n111), .ZN(n22659) );
  INV_X1 U16018 ( .A(n110), .ZN(n22660) );
  INV_X1 U16019 ( .A(n110), .ZN(n22661) );
  INV_X1 U16020 ( .A(n109), .ZN(n22662) );
  INV_X1 U16021 ( .A(n109), .ZN(n22663) );
  INV_X1 U16022 ( .A(n108), .ZN(n22664) );
  INV_X1 U16023 ( .A(n108), .ZN(n22665) );
  INV_X1 U16024 ( .A(n107), .ZN(n22666) );
  INV_X1 U16025 ( .A(n107), .ZN(n22667) );
  INV_X1 U16026 ( .A(n106), .ZN(n22668) );
  INV_X1 U16027 ( .A(n106), .ZN(n22669) );
  INV_X1 U16028 ( .A(n105), .ZN(n22670) );
  INV_X1 U16029 ( .A(n105), .ZN(n22671) );
  INV_X1 U16030 ( .A(n104), .ZN(n22672) );
  INV_X1 U16031 ( .A(n104), .ZN(n22673) );
  OAI21_X1 U16032 ( .B1(n17999), .B2(n27299), .A(n24680), .ZN(r899_B_6_) );
  INV_X1 U16033 ( .A(n103), .ZN(n22674) );
  INV_X1 U16034 ( .A(n103), .ZN(n22675) );
  INV_X1 U16035 ( .A(n18453), .ZN(n22676) );
  INV_X1 U16036 ( .A(n18453), .ZN(n22677) );
  INV_X1 U16037 ( .A(n18454), .ZN(n22678) );
  INV_X1 U16038 ( .A(n18454), .ZN(n22679) );
  INV_X1 U16039 ( .A(n18455), .ZN(n22680) );
  INV_X1 U16040 ( .A(n18456), .ZN(n22681) );
  INV_X1 U16041 ( .A(n18457), .ZN(n22682) );
  INV_X1 U16042 ( .A(n18457), .ZN(n22683) );
  INV_X1 U16043 ( .A(n27260), .ZN(n22684) );
  INV_X1 U16044 ( .A(n22684), .ZN(n22685) );
  INV_X1 U16045 ( .A(n22684), .ZN(n22686) );
  INV_X1 U16046 ( .A(n18458), .ZN(n22687) );
  INV_X1 U16047 ( .A(n18459), .ZN(n22688) );
  INV_X1 U16048 ( .A(n18460), .ZN(n22689) );
  INV_X1 U16049 ( .A(n3988), .ZN(n22690) );
  INV_X1 U16050 ( .A(n22690), .ZN(n22691) );
  INV_X1 U16051 ( .A(n22690), .ZN(n22692) );
  INV_X1 U16052 ( .A(n18461), .ZN(n22693) );
  INV_X1 U16053 ( .A(n26637), .ZN(n22694) );
  INV_X1 U16054 ( .A(n26638), .ZN(n22695) );
  INV_X1 U16055 ( .A(n22695), .ZN(n22696) );
  INV_X1 U16056 ( .A(n18462), .ZN(n22697) );
  INV_X1 U16057 ( .A(n18462), .ZN(n22698) );
  INV_X1 U16058 ( .A(n26640), .ZN(n22699) );
  INV_X1 U16059 ( .A(n22699), .ZN(n22700) );
  INV_X1 U16060 ( .A(n18463), .ZN(n22701) );
  INV_X1 U16061 ( .A(n18463), .ZN(n22702) );
  INV_X1 U16062 ( .A(n18464), .ZN(n22703) );
  INV_X1 U16063 ( .A(n18465), .ZN(n22704) );
  INV_X1 U16064 ( .A(n18465), .ZN(n22705) );
  INV_X1 U16065 ( .A(n18466), .ZN(n22706) );
  INV_X1 U16066 ( .A(n18467), .ZN(n22707) );
  INV_X1 U16067 ( .A(n18467), .ZN(n22708) );
  INV_X1 U16068 ( .A(n26644), .ZN(n22709) );
  INV_X1 U16069 ( .A(n22709), .ZN(n22710) );
  INV_X1 U16070 ( .A(n18468), .ZN(n22711) );
  INV_X1 U16071 ( .A(n18468), .ZN(n22712) );
  INV_X1 U16072 ( .A(n18469), .ZN(n22713) );
  INV_X1 U16073 ( .A(n18470), .ZN(n22714) );
  INV_X1 U16074 ( .A(n18470), .ZN(n22715) );
  INV_X1 U16075 ( .A(n18471), .ZN(n22716) );
  INV_X1 U16076 ( .A(n18472), .ZN(n22717) );
  INV_X1 U16077 ( .A(n18472), .ZN(n22718) );
  INV_X1 U16078 ( .A(n18473), .ZN(n22719) );
  INV_X1 U16079 ( .A(n18474), .ZN(n22720) );
  INV_X1 U16080 ( .A(n18474), .ZN(n22721) );
  INV_X1 U16081 ( .A(n18475), .ZN(n22722) );
  INV_X1 U16082 ( .A(n18476), .ZN(n22723) );
  INV_X1 U16083 ( .A(n18476), .ZN(n22724) );
  INV_X1 U16084 ( .A(n18477), .ZN(n22725) );
  INV_X1 U16085 ( .A(n26652), .ZN(n22726) );
  INV_X1 U16086 ( .A(n22726), .ZN(n22727) );
  INV_X1 U16087 ( .A(n22726), .ZN(n22728) );
  INV_X1 U16088 ( .A(n18478), .ZN(n22729) );
  INV_X1 U16089 ( .A(n18479), .ZN(n22730) );
  INV_X1 U16090 ( .A(n18479), .ZN(n22731) );
  INV_X1 U16091 ( .A(n18480), .ZN(n22732) );
  INV_X1 U16092 ( .A(n19290), .ZN(n22733) );
  INV_X1 U16093 ( .A(n22733), .ZN(n22734) );
  INV_X1 U16094 ( .A(n22733), .ZN(n22735) );
  INV_X1 U16095 ( .A(n26666), .ZN(n22736) );
  INV_X1 U16096 ( .A(n22736), .ZN(n22737) );
  INV_X1 U16097 ( .A(n26667), .ZN(n22738) );
  INV_X1 U16098 ( .A(n22738), .ZN(n22739) );
  INV_X1 U16099 ( .A(n22738), .ZN(n22740) );
  INV_X1 U16100 ( .A(n26669), .ZN(n22741) );
  INV_X1 U16101 ( .A(n22741), .ZN(n22742) );
  INV_X1 U16102 ( .A(n19292), .ZN(n22743) );
  INV_X1 U16103 ( .A(n22743), .ZN(n22744) );
  INV_X1 U16104 ( .A(n22743), .ZN(n22745) );
  INV_X1 U16105 ( .A(n20498), .ZN(n22746) );
  INV_X1 U16106 ( .A(n22746), .ZN(n22747) );
  INV_X1 U16107 ( .A(n18481), .ZN(n22748) );
  INV_X1 U16108 ( .A(n18481), .ZN(n22749) );
  INV_X1 U16109 ( .A(n20496), .ZN(n22750) );
  INV_X1 U16110 ( .A(n22750), .ZN(n22751) );
  INV_X1 U16111 ( .A(n18482), .ZN(n22752) );
  INV_X1 U16112 ( .A(n18482), .ZN(n22753) );
  INV_X1 U16113 ( .A(n18483), .ZN(n22754) );
  INV_X1 U16114 ( .A(n19295), .ZN(n22755) );
  INV_X1 U16115 ( .A(n22755), .ZN(n22756) );
  INV_X1 U16116 ( .A(n22755), .ZN(n22757) );
  INV_X1 U16117 ( .A(n26679), .ZN(n22758) );
  INV_X1 U16118 ( .A(n22758), .ZN(n22759) );
  INV_X1 U16119 ( .A(n22758), .ZN(n22760) );
  INV_X1 U16120 ( .A(n26683), .ZN(n22761) );
  INV_X1 U16121 ( .A(n22761), .ZN(n22762) );
  INV_X1 U16122 ( .A(n22761), .ZN(n22763) );
  INV_X1 U16123 ( .A(n18484), .ZN(n22764) );
  INV_X1 U16124 ( .A(n26687), .ZN(n22765) );
  INV_X1 U16125 ( .A(n22765), .ZN(n22766) );
  INV_X1 U16126 ( .A(n22765), .ZN(n22767) );
  INV_X1 U16127 ( .A(n26693), .ZN(n22768) );
  INV_X1 U16128 ( .A(n22768), .ZN(n22769) );
  INV_X1 U16129 ( .A(n22768), .ZN(n22770) );
  INV_X1 U16130 ( .A(n18485), .ZN(n22771) );
  INV_X1 U16131 ( .A(n26696), .ZN(n22772) );
  INV_X1 U16132 ( .A(n22772), .ZN(n22773) );
  INV_X1 U16133 ( .A(n22772), .ZN(n22774) );
  INV_X1 U16134 ( .A(n26699), .ZN(n22775) );
  INV_X1 U16135 ( .A(n22775), .ZN(n22776) );
  INV_X1 U16136 ( .A(n22775), .ZN(n22777) );
  INV_X1 U16137 ( .A(n26702), .ZN(n22778) );
  INV_X1 U16138 ( .A(n22778), .ZN(n22779) );
  INV_X1 U16139 ( .A(n26705), .ZN(n22780) );
  INV_X1 U16140 ( .A(n22780), .ZN(n22781) );
  INV_X1 U16141 ( .A(n26708), .ZN(n22782) );
  INV_X1 U16142 ( .A(n22782), .ZN(n22783) );
  INV_X1 U16143 ( .A(n50780), .ZN(n22784) );
  INV_X1 U16144 ( .A(n22784), .ZN(n22785) );
  INV_X1 U16145 ( .A(n18486), .ZN(n22786) );
  INV_X1 U16146 ( .A(n18486), .ZN(n22787) );
  INV_X1 U16147 ( .A(n26712), .ZN(n22788) );
  INV_X1 U16148 ( .A(n22788), .ZN(n22789) );
  INV_X1 U16149 ( .A(n18487), .ZN(n22790) );
  INV_X1 U16150 ( .A(n18487), .ZN(n22791) );
  INV_X1 U16151 ( .A(n18488), .ZN(n22792) );
  INV_X1 U16152 ( .A(n18488), .ZN(n22793) );
  INV_X1 U16153 ( .A(n18489), .ZN(n22794) );
  INV_X1 U16154 ( .A(n18489), .ZN(n22795) );
  INV_X1 U16155 ( .A(n18490), .ZN(n22796) );
  INV_X1 U16156 ( .A(n18490), .ZN(n22797) );
  INV_X1 U16157 ( .A(n18491), .ZN(n22798) );
  INV_X1 U16158 ( .A(n18492), .ZN(n22799) );
  INV_X1 U16159 ( .A(n18492), .ZN(n22800) );
  INV_X1 U16160 ( .A(n18493), .ZN(n22801) );
  INV_X1 U16161 ( .A(n18494), .ZN(n22802) );
  INV_X1 U16162 ( .A(n18494), .ZN(n22803) );
  INV_X1 U16163 ( .A(n25288), .ZN(n22804) );
  INV_X1 U16164 ( .A(n22804), .ZN(n22805) );
  INV_X1 U16165 ( .A(n22804), .ZN(n22806) );
  INV_X1 U16166 ( .A(n3236), .ZN(n22807) );
  INV_X1 U16167 ( .A(n22807), .ZN(n22808) );
  INV_X1 U16168 ( .A(n3443), .ZN(n22809) );
  INV_X1 U16169 ( .A(n22809), .ZN(n22810) );
  INV_X1 U16170 ( .A(n26738), .ZN(n22811) );
  INV_X1 U16171 ( .A(n22811), .ZN(n22812) );
  INV_X1 U16172 ( .A(n22811), .ZN(n22813) );
  INV_X1 U16173 ( .A(n26744), .ZN(n22814) );
  INV_X1 U16174 ( .A(n22814), .ZN(n22815) );
  INV_X1 U16175 ( .A(n22814), .ZN(n22816) );
  INV_X1 U16176 ( .A(n18495), .ZN(n22817) );
  INV_X1 U16177 ( .A(n18495), .ZN(n22818) );
  INV_X1 U16178 ( .A(n256301), .ZN(n22819) );
  INV_X1 U16179 ( .A(n22819), .ZN(n22820) );
  INV_X1 U16180 ( .A(n22819), .ZN(n22821) );
  INV_X1 U16181 ( .A(n25633), .ZN(n22822) );
  INV_X1 U16182 ( .A(n22822), .ZN(n22823) );
  INV_X1 U16183 ( .A(n22822), .ZN(n22824) );
  INV_X1 U16184 ( .A(n26754), .ZN(n22825) );
  INV_X1 U16185 ( .A(n22825), .ZN(n22826) );
  INV_X1 U16186 ( .A(n22825), .ZN(n22827) );
  INV_X1 U16187 ( .A(n26998), .ZN(n22828) );
  INV_X1 U16188 ( .A(n26757), .ZN(n22829) );
  INV_X1 U16189 ( .A(n22829), .ZN(n22830) );
  INV_X1 U16190 ( .A(n22829), .ZN(n22831) );
  INV_X1 U16191 ( .A(n18497), .ZN(n22832) );
  INV_X1 U16192 ( .A(n18497), .ZN(n22833) );
  INV_X1 U16193 ( .A(n26064), .ZN(n22834) );
  INV_X1 U16194 ( .A(n22834), .ZN(n22835) );
  INV_X1 U16195 ( .A(n22834), .ZN(n22836) );
  INV_X1 U16196 ( .A(n26552), .ZN(n22837) );
  INV_X1 U16197 ( .A(n22837), .ZN(n22838) );
  INV_X1 U16198 ( .A(n22837), .ZN(n22839) );
  INV_X1 U16199 ( .A(n18498), .ZN(n22840) );
  INV_X1 U16200 ( .A(n18498), .ZN(n22841) );
  INV_X1 U16201 ( .A(n18499), .ZN(n22842) );
  INV_X1 U16202 ( .A(n18499), .ZN(n22843) );
  INV_X1 U16203 ( .A(n18500), .ZN(n22844) );
  INV_X1 U16204 ( .A(n18500), .ZN(n22845) );
  INV_X1 U16205 ( .A(n26034), .ZN(n22846) );
  INV_X1 U16206 ( .A(n22846), .ZN(n22847) );
  INV_X1 U16207 ( .A(n22846), .ZN(n22848) );
  INV_X1 U16208 ( .A(n20715), .ZN(n22849) );
  INV_X1 U16209 ( .A(n18115), .ZN(n22850) );
  INV_X1 U16210 ( .A(n18501), .ZN(n22851) );
  INV_X1 U16211 ( .A(n18501), .ZN(n22852) );
  INV_X1 U16212 ( .A(n26021), .ZN(n22853) );
  INV_X1 U16213 ( .A(n22853), .ZN(n22854) );
  INV_X1 U16214 ( .A(n22853), .ZN(n22855) );
  INV_X1 U16215 ( .A(n18502), .ZN(n22856) );
  INV_X1 U16216 ( .A(n18502), .ZN(n22857) );
  INV_X1 U16217 ( .A(n26017), .ZN(n22858) );
  INV_X1 U16218 ( .A(n22858), .ZN(n22859) );
  INV_X1 U16219 ( .A(n22858), .ZN(n22860) );
  INV_X1 U16220 ( .A(n18503), .ZN(n22861) );
  INV_X1 U16221 ( .A(n18503), .ZN(n22862) );
  INV_X1 U16222 ( .A(n26012), .ZN(n22863) );
  INV_X1 U16223 ( .A(n22863), .ZN(n22864) );
  INV_X1 U16224 ( .A(n22863), .ZN(n22865) );
  INV_X1 U16225 ( .A(n18504), .ZN(n22866) );
  INV_X1 U16226 ( .A(n18504), .ZN(n22867) );
  INV_X1 U16227 ( .A(n26008), .ZN(n22868) );
  INV_X1 U16228 ( .A(n22868), .ZN(n22869) );
  INV_X1 U16229 ( .A(n22868), .ZN(n22870) );
  INV_X1 U16230 ( .A(n24430), .ZN(n22871) );
  INV_X1 U16231 ( .A(n18505), .ZN(n22872) );
  INV_X1 U16232 ( .A(n18505), .ZN(n22873) );
  INV_X1 U16233 ( .A(n25998), .ZN(n22874) );
  INV_X1 U16234 ( .A(n22874), .ZN(n22875) );
  INV_X1 U16235 ( .A(n22874), .ZN(n22876) );
  INV_X1 U16236 ( .A(n18506), .ZN(n22877) );
  INV_X1 U16237 ( .A(n18506), .ZN(n22878) );
  INV_X1 U16238 ( .A(n18507), .ZN(n22879) );
  INV_X1 U16239 ( .A(n18507), .ZN(n22880) );
  INV_X1 U16240 ( .A(n18508), .ZN(n22881) );
  INV_X1 U16241 ( .A(n18508), .ZN(n22882) );
  INV_X1 U16242 ( .A(n18509), .ZN(n22883) );
  INV_X1 U16243 ( .A(n18509), .ZN(n22884) );
  INV_X1 U16244 ( .A(n18510), .ZN(n22885) );
  INV_X1 U16245 ( .A(n18510), .ZN(n22886) );
  INV_X1 U16246 ( .A(n18511), .ZN(n22887) );
  INV_X1 U16247 ( .A(n18511), .ZN(n22888) );
  INV_X1 U16248 ( .A(n18903), .ZN(n22889) );
  INV_X1 U16249 ( .A(n22889), .ZN(n22890) );
  INV_X1 U16250 ( .A(n22889), .ZN(n22891) );
  INV_X1 U16251 ( .A(n18512), .ZN(n22892) );
  INV_X1 U16252 ( .A(n18512), .ZN(n22893) );
  INV_X1 U16253 ( .A(n5305), .ZN(n22894) );
  INV_X1 U16254 ( .A(n22894), .ZN(n22895) );
  INV_X1 U16255 ( .A(n22894), .ZN(n22896) );
  CLKBUF_X1 U16256 ( .A(n27177), .Z(n22897) );
  INV_X1 U16257 ( .A(n19316), .ZN(n22898) );
  INV_X1 U16258 ( .A(n22898), .ZN(n22899) );
  INV_X1 U16259 ( .A(n22898), .ZN(n22900) );
  CLKBUF_X1 U16260 ( .A(n27232), .Z(n22901) );
  INV_X1 U16261 ( .A(n19317), .ZN(n22902) );
  INV_X1 U16262 ( .A(n22902), .ZN(n22903) );
  INV_X1 U16263 ( .A(n22902), .ZN(n22904) );
  INV_X1 U16264 ( .A(n27186), .ZN(n22905) );
  INV_X1 U16265 ( .A(n22905), .ZN(n22906) );
  INV_X1 U16266 ( .A(n22905), .ZN(n22907) );
  INV_X1 U16267 ( .A(n27184), .ZN(n22908) );
  INV_X1 U16268 ( .A(n22908), .ZN(n22909) );
  INV_X1 U16269 ( .A(n22908), .ZN(n22910) );
  INV_X1 U16270 ( .A(n27182), .ZN(n22911) );
  INV_X1 U16271 ( .A(n22911), .ZN(n22912) );
  INV_X1 U16272 ( .A(n22911), .ZN(n22913) );
  INV_X1 U16273 ( .A(n27180), .ZN(n22914) );
  INV_X1 U16274 ( .A(n22914), .ZN(n22915) );
  INV_X1 U16275 ( .A(n22914), .ZN(n22916) );
  INV_X1 U16276 ( .A(n27241), .ZN(n22917) );
  INV_X1 U16277 ( .A(n22917), .ZN(n22918) );
  INV_X1 U16278 ( .A(n22917), .ZN(n22919) );
  INV_X1 U16279 ( .A(n27239), .ZN(n22920) );
  INV_X1 U16280 ( .A(n22920), .ZN(n22921) );
  INV_X1 U16281 ( .A(n22920), .ZN(n22922) );
  INV_X1 U16282 ( .A(n27237), .ZN(n22923) );
  INV_X1 U16283 ( .A(n22923), .ZN(n22924) );
  INV_X1 U16284 ( .A(n22923), .ZN(n22925) );
  INV_X1 U16285 ( .A(n27235), .ZN(n22926) );
  INV_X1 U16286 ( .A(n22926), .ZN(n22927) );
  INV_X1 U16287 ( .A(n22926), .ZN(n22928) );
  INV_X1 U16288 ( .A(n27164), .ZN(n22929) );
  INV_X1 U16289 ( .A(n22929), .ZN(n22930) );
  INV_X1 U16290 ( .A(n22929), .ZN(n22931) );
  INV_X1 U16291 ( .A(n27162), .ZN(n22932) );
  INV_X1 U16292 ( .A(n22932), .ZN(n22933) );
  INV_X1 U16293 ( .A(n22932), .ZN(n22934) );
  INV_X1 U16294 ( .A(n27252), .ZN(n22935) );
  INV_X1 U16295 ( .A(n22935), .ZN(n22936) );
  INV_X1 U16296 ( .A(n22935), .ZN(n22937) );
  INV_X1 U16297 ( .A(n27250), .ZN(n22938) );
  INV_X1 U16298 ( .A(n22938), .ZN(n22939) );
  INV_X1 U16299 ( .A(n22938), .ZN(n22940) );
  INV_X1 U16300 ( .A(n27073), .ZN(n22941) );
  INV_X1 U16301 ( .A(n22941), .ZN(n22942) );
  INV_X1 U16302 ( .A(n22941), .ZN(n22943) );
  INV_X1 U16303 ( .A(n21397), .ZN(n22944) );
  INV_X1 U16304 ( .A(n22944), .ZN(n22945) );
  INV_X1 U16305 ( .A(n22944), .ZN(n22946) );
  INV_X1 U16306 ( .A(n26993), .ZN(n22947) );
  INV_X1 U16307 ( .A(n22947), .ZN(n22948) );
  INV_X1 U16308 ( .A(n22947), .ZN(n22949) );
  INV_X1 U16309 ( .A(n18513), .ZN(n22950) );
  INV_X1 U16310 ( .A(n18513), .ZN(n22951) );
  INV_X1 U16311 ( .A(n18515), .ZN(n22952) );
  INV_X1 U16312 ( .A(n18515), .ZN(n22953) );
  INV_X1 U16313 ( .A(n18516), .ZN(n22954) );
  INV_X1 U16314 ( .A(n18516), .ZN(n22955) );
  INV_X1 U16315 ( .A(n19318), .ZN(n22956) );
  INV_X1 U16316 ( .A(n22956), .ZN(n22957) );
  INV_X1 U16317 ( .A(n22956), .ZN(n22958) );
  INV_X1 U16318 ( .A(n27072), .ZN(n22959) );
  INV_X1 U16319 ( .A(n22959), .ZN(n22960) );
  INV_X1 U16320 ( .A(n22959), .ZN(n22961) );
  INV_X1 U16321 ( .A(n22943), .ZN(n22962) );
  INV_X1 U16322 ( .A(n22943), .ZN(n22963) );
  INV_X1 U16323 ( .A(n27109), .ZN(n22964) );
  INV_X1 U16324 ( .A(n22964), .ZN(n22965) );
  INV_X1 U16325 ( .A(n22964), .ZN(n22966) );
  INV_X1 U16326 ( .A(n27129), .ZN(n22967) );
  INV_X1 U16327 ( .A(n22967), .ZN(n22968) );
  INV_X1 U16328 ( .A(n25088), .ZN(n22969) );
  INV_X1 U16329 ( .A(n27277), .ZN(n22970) );
  INV_X1 U16330 ( .A(n22970), .ZN(n22971) );
  INV_X1 U16331 ( .A(n25085), .ZN(n22972) );
  INV_X1 U16332 ( .A(n277901), .ZN(n22973) );
  INV_X1 U16333 ( .A(n277901), .ZN(n22974) );
  INV_X1 U16334 ( .A(n18517), .ZN(n22975) );
  INV_X1 U16335 ( .A(n18517), .ZN(n22976) );
  INV_X1 U16336 ( .A(n18518), .ZN(n22977) );
  INV_X1 U16337 ( .A(n18518), .ZN(n22978) );
  INV_X1 U16338 ( .A(n18519), .ZN(n22979) );
  INV_X1 U16339 ( .A(n18519), .ZN(n22980) );
  INV_X1 U16340 ( .A(n25682), .ZN(n22981) );
  INV_X1 U16341 ( .A(n22981), .ZN(n22982) );
  INV_X1 U16342 ( .A(n22981), .ZN(n22983) );
  INV_X1 U16343 ( .A(n18520), .ZN(n22984) );
  INV_X1 U16344 ( .A(n18520), .ZN(n22985) );
  INV_X1 U16345 ( .A(n18521), .ZN(n22986) );
  INV_X1 U16346 ( .A(n18521), .ZN(n22987) );
  INV_X1 U16347 ( .A(n25695), .ZN(n22988) );
  INV_X1 U16348 ( .A(n22988), .ZN(n22989) );
  INV_X1 U16349 ( .A(n22988), .ZN(n22990) );
  INV_X1 U16350 ( .A(n25682), .ZN(n22991) );
  INV_X1 U16351 ( .A(n22991), .ZN(n22992) );
  INV_X1 U16352 ( .A(n22991), .ZN(n22993) );
  INV_X1 U16353 ( .A(n18522), .ZN(n22994) );
  INV_X1 U16354 ( .A(n18522), .ZN(n22995) );
  INV_X1 U16355 ( .A(n25946), .ZN(n22996) );
  INV_X1 U16356 ( .A(n25946), .ZN(n22997) );
  INV_X1 U16357 ( .A(n25695), .ZN(n22998) );
  INV_X1 U16358 ( .A(n22998), .ZN(n22999) );
  INV_X1 U16359 ( .A(n22998), .ZN(n23000) );
  INV_X1 U16360 ( .A(n27146), .ZN(n23001) );
  INV_X1 U16361 ( .A(n27146), .ZN(n23002) );
  INV_X1 U16362 ( .A(n18523), .ZN(n23003) );
  INV_X1 U16363 ( .A(n18523), .ZN(n23004) );
  INV_X1 U16364 ( .A(n25954), .ZN(n23005) );
  INV_X1 U16365 ( .A(n25954), .ZN(n23006) );
  INV_X1 U16366 ( .A(n27145), .ZN(n23007) );
  INV_X1 U16367 ( .A(n27145), .ZN(n23008) );
  INV_X1 U16368 ( .A(n18524), .ZN(n23009) );
  INV_X1 U16369 ( .A(n18524), .ZN(n23010) );
  INV_X1 U16370 ( .A(n19030), .ZN(n23011) );
  INV_X1 U16371 ( .A(n23011), .ZN(n23012) );
  INV_X1 U16372 ( .A(n23011), .ZN(n23013) );
  INV_X1 U16373 ( .A(n21400), .ZN(n23014) );
  INV_X1 U16374 ( .A(n23014), .ZN(n23015) );
  INV_X1 U16375 ( .A(n18525), .ZN(n23016) );
  INV_X1 U16376 ( .A(n18525), .ZN(n23017) );
  INV_X1 U16377 ( .A(n18526), .ZN(n23018) );
  INV_X1 U16378 ( .A(n18526), .ZN(n23019) );
  INV_X1 U16379 ( .A(n20492), .ZN(n23020) );
  INV_X1 U16380 ( .A(n20492), .ZN(n23021) );
  INV_X1 U16381 ( .A(n18527), .ZN(n23022) );
  INV_X1 U16382 ( .A(n18527), .ZN(n23023) );
  INV_X1 U16383 ( .A(n18528), .ZN(n23024) );
  INV_X1 U16384 ( .A(n18528), .ZN(n23025) );
  INV_X1 U16385 ( .A(n18529), .ZN(n23026) );
  INV_X1 U16386 ( .A(n18529), .ZN(n23027) );
  INV_X1 U16387 ( .A(n18530), .ZN(n23028) );
  INV_X1 U16388 ( .A(n18530), .ZN(n23029) );
  INV_X1 U16389 ( .A(n18531), .ZN(n23030) );
  INV_X1 U16390 ( .A(n18531), .ZN(n23031) );
  INV_X1 U16391 ( .A(n18532), .ZN(n23032) );
  INV_X1 U16392 ( .A(n18532), .ZN(n23033) );
  INV_X1 U16393 ( .A(n18533), .ZN(n23034) );
  INV_X1 U16394 ( .A(n18533), .ZN(n23035) );
  INV_X1 U16395 ( .A(n18534), .ZN(n23036) );
  INV_X1 U16396 ( .A(n18534), .ZN(n23037) );
  INV_X1 U16397 ( .A(n18535), .ZN(n23038) );
  INV_X1 U16398 ( .A(n18535), .ZN(n23039) );
  INV_X1 U16399 ( .A(n18536), .ZN(n23040) );
  INV_X1 U16400 ( .A(n18536), .ZN(n23041) );
  INV_X1 U16401 ( .A(n18537), .ZN(n23042) );
  INV_X1 U16402 ( .A(n18537), .ZN(n23043) );
  INV_X1 U16403 ( .A(n18538), .ZN(n23044) );
  INV_X1 U16404 ( .A(n18538), .ZN(n23045) );
  INV_X1 U16405 ( .A(n18539), .ZN(n23046) );
  INV_X1 U16406 ( .A(n18539), .ZN(n23047) );
  INV_X1 U16407 ( .A(n18540), .ZN(n23048) );
  INV_X1 U16408 ( .A(n18540), .ZN(n23049) );
  INV_X1 U16409 ( .A(n18541), .ZN(n23050) );
  INV_X1 U16410 ( .A(n18541), .ZN(n23051) );
  INV_X1 U16411 ( .A(n18542), .ZN(n23052) );
  INV_X1 U16412 ( .A(n18542), .ZN(n23053) );
  INV_X1 U16413 ( .A(n18543), .ZN(n23054) );
  INV_X1 U16414 ( .A(n18543), .ZN(n23055) );
  INV_X1 U16415 ( .A(n18544), .ZN(n23056) );
  INV_X1 U16416 ( .A(n18544), .ZN(n23057) );
  INV_X1 U16417 ( .A(n18545), .ZN(n23058) );
  INV_X1 U16418 ( .A(n18545), .ZN(n23059) );
  INV_X1 U16419 ( .A(n18546), .ZN(n23060) );
  INV_X1 U16420 ( .A(n18546), .ZN(n23061) );
  INV_X1 U16421 ( .A(n32600), .ZN(n23062) );
  INV_X1 U16422 ( .A(n32600), .ZN(n23063) );
  INV_X1 U16423 ( .A(n18547), .ZN(n23064) );
  INV_X1 U16424 ( .A(n18547), .ZN(n23065) );
  INV_X1 U16425 ( .A(n18548), .ZN(n23066) );
  INV_X1 U16426 ( .A(n18548), .ZN(n23067) );
  INV_X1 U16427 ( .A(n25883), .ZN(n23068) );
  INV_X1 U16428 ( .A(n23068), .ZN(n23069) );
  INV_X1 U16429 ( .A(n23068), .ZN(n23070) );
  INV_X1 U16430 ( .A(n18549), .ZN(n23071) );
  INV_X1 U16431 ( .A(n18549), .ZN(n23072) );
  INV_X1 U16432 ( .A(n18550), .ZN(n23073) );
  INV_X1 U16433 ( .A(n18550), .ZN(n23074) );
  INV_X1 U16434 ( .A(n18551), .ZN(n23075) );
  INV_X1 U16435 ( .A(n18551), .ZN(n23076) );
  INV_X1 U16436 ( .A(n18552), .ZN(n23077) );
  INV_X1 U16437 ( .A(n18552), .ZN(n23078) );
  INV_X1 U16438 ( .A(n18553), .ZN(n23079) );
  INV_X1 U16439 ( .A(n18553), .ZN(n23080) );
  INV_X1 U16440 ( .A(n18554), .ZN(n23081) );
  INV_X1 U16441 ( .A(n18554), .ZN(n23082) );
  INV_X1 U16442 ( .A(n18555), .ZN(n23083) );
  INV_X1 U16443 ( .A(n18555), .ZN(n23084) );
  INV_X1 U16444 ( .A(n18556), .ZN(n23085) );
  INV_X1 U16445 ( .A(n18556), .ZN(n23086) );
  INV_X1 U16446 ( .A(n18557), .ZN(n23087) );
  INV_X1 U16447 ( .A(n18557), .ZN(n23088) );
  INV_X1 U16448 ( .A(n3160), .ZN(n23089) );
  INV_X1 U16449 ( .A(n3987), .ZN(n23090) );
  INV_X1 U16450 ( .A(n17128), .ZN(n23091) );
  INV_X1 U16451 ( .A(n17126), .ZN(n23092) );
  INV_X1 U16452 ( .A(n17128), .ZN(n23093) );
  INV_X1 U16453 ( .A(n4163), .ZN(n23094) );
  INV_X1 U16454 ( .A(n4163), .ZN(n23095) );
  INV_X1 U16455 ( .A(n18558), .ZN(n23096) );
  INV_X1 U16456 ( .A(n18558), .ZN(n23097) );
  INV_X1 U16457 ( .A(n31280), .ZN(n23098) );
  INV_X1 U16458 ( .A(n31280), .ZN(n23099) );
  INV_X1 U16459 ( .A(n18559), .ZN(n23100) );
  INV_X1 U16460 ( .A(n18560), .ZN(n23101) );
  INV_X1 U16461 ( .A(n18560), .ZN(n23102) );
  INV_X1 U16462 ( .A(n18561), .ZN(n23103) );
  INV_X1 U16463 ( .A(n18561), .ZN(n23104) );
  INV_X1 U16464 ( .A(n18562), .ZN(n23105) );
  INV_X1 U16465 ( .A(n18562), .ZN(n23106) );
  INV_X1 U16466 ( .A(n18563), .ZN(n23107) );
  INV_X1 U16467 ( .A(n18563), .ZN(n23108) );
  INV_X1 U16468 ( .A(n18564), .ZN(n23109) );
  INV_X1 U16469 ( .A(n18564), .ZN(n23110) );
  INV_X1 U16470 ( .A(n18565), .ZN(n23111) );
  INV_X1 U16471 ( .A(n18565), .ZN(n23112) );
  INV_X1 U16472 ( .A(n18566), .ZN(n23113) );
  INV_X1 U16473 ( .A(n27804), .ZN(n23114) );
  INV_X1 U16474 ( .A(n23114), .ZN(n23115) );
  INV_X1 U16475 ( .A(n23114), .ZN(n23116) );
  INV_X1 U16476 ( .A(n18567), .ZN(n23117) );
  INV_X1 U16477 ( .A(n18567), .ZN(n23118) );
  INV_X1 U16478 ( .A(n18568), .ZN(n23119) );
  INV_X1 U16479 ( .A(n18568), .ZN(n23120) );
  INV_X1 U16480 ( .A(n18569), .ZN(n23121) );
  INV_X1 U16481 ( .A(n18569), .ZN(n23122) );
  INV_X1 U16482 ( .A(n18570), .ZN(n23123) );
  INV_X1 U16483 ( .A(n18570), .ZN(n23124) );
  INV_X1 U16484 ( .A(n18571), .ZN(n23125) );
  INV_X1 U16485 ( .A(n18571), .ZN(n23126) );
  INV_X1 U16486 ( .A(n18572), .ZN(n23127) );
  INV_X1 U16487 ( .A(n18572), .ZN(n23128) );
  INV_X1 U16488 ( .A(n18573), .ZN(n23129) );
  INV_X1 U16489 ( .A(n18573), .ZN(n23130) );
  INV_X1 U16490 ( .A(n259901), .ZN(n23131) );
  INV_X1 U16491 ( .A(n23131), .ZN(n23132) );
  INV_X1 U16492 ( .A(n23131), .ZN(n23133) );
  INV_X1 U16493 ( .A(n18574), .ZN(n23134) );
  INV_X1 U16494 ( .A(n18574), .ZN(n23135) );
  INV_X1 U16495 ( .A(n18575), .ZN(n23136) );
  INV_X1 U16496 ( .A(n18575), .ZN(n23137) );
  INV_X1 U16497 ( .A(n18576), .ZN(n23138) );
  INV_X1 U16498 ( .A(n18576), .ZN(n23139) );
  INV_X1 U16499 ( .A(n25994), .ZN(n23140) );
  INV_X1 U16500 ( .A(n23140), .ZN(n23141) );
  INV_X1 U16501 ( .A(n23140), .ZN(n23142) );
  INV_X1 U16502 ( .A(n18577), .ZN(n23143) );
  INV_X1 U16503 ( .A(n18577), .ZN(n23144) );
  INV_X1 U16504 ( .A(n25999), .ZN(n23145) );
  INV_X1 U16505 ( .A(n23145), .ZN(n23146) );
  INV_X1 U16506 ( .A(n23145), .ZN(n23147) );
  INV_X1 U16507 ( .A(n18578), .ZN(n23148) );
  INV_X1 U16508 ( .A(n18578), .ZN(n23149) );
  INV_X1 U16509 ( .A(n18579), .ZN(n23150) );
  INV_X1 U16510 ( .A(n18579), .ZN(n23151) );
  INV_X1 U16511 ( .A(n27196), .ZN(n23152) );
  INV_X1 U16512 ( .A(n23152), .ZN(n23153) );
  INV_X1 U16513 ( .A(n23152), .ZN(n23154) );
  INV_X1 U16514 ( .A(n18580), .ZN(n23155) );
  INV_X1 U16515 ( .A(n18580), .ZN(n23156) );
  INV_X1 U16516 ( .A(n26013), .ZN(n23157) );
  INV_X1 U16517 ( .A(n23157), .ZN(n23158) );
  INV_X1 U16518 ( .A(n23157), .ZN(n23159) );
  INV_X1 U16519 ( .A(n18581), .ZN(n23160) );
  INV_X1 U16520 ( .A(n18581), .ZN(n23161) );
  INV_X1 U16521 ( .A(n27218), .ZN(n23162) );
  INV_X1 U16522 ( .A(n23162), .ZN(n23163) );
  INV_X1 U16523 ( .A(n23162), .ZN(n23164) );
  INV_X1 U16524 ( .A(n18582), .ZN(n23165) );
  INV_X1 U16525 ( .A(n18582), .ZN(n23166) );
  INV_X1 U16526 ( .A(n25999), .ZN(n23167) );
  INV_X1 U16527 ( .A(n23167), .ZN(n23168) );
  INV_X1 U16528 ( .A(n23167), .ZN(n23169) );
  INV_X1 U16529 ( .A(n27799), .ZN(n23170) );
  INV_X1 U16530 ( .A(n23170), .ZN(n23171) );
  INV_X1 U16531 ( .A(n23170), .ZN(n23172) );
  INV_X1 U16532 ( .A(n27174), .ZN(n23173) );
  INV_X1 U16533 ( .A(n23173), .ZN(n23174) );
  INV_X1 U16534 ( .A(n23173), .ZN(n23175) );
  INV_X1 U16535 ( .A(n18583), .ZN(n23176) );
  INV_X1 U16536 ( .A(n18583), .ZN(n23177) );
  INV_X1 U16537 ( .A(n18584), .ZN(n23178) );
  INV_X1 U16538 ( .A(n18584), .ZN(n23179) );
  INV_X1 U16539 ( .A(n27218), .ZN(n23180) );
  INV_X1 U16540 ( .A(n23180), .ZN(n23181) );
  INV_X1 U16541 ( .A(n23180), .ZN(n23182) );
  INV_X1 U16542 ( .A(n27196), .ZN(n23183) );
  INV_X1 U16543 ( .A(n23183), .ZN(n23184) );
  INV_X1 U16544 ( .A(n23183), .ZN(n23185) );
  INV_X1 U16545 ( .A(n18585), .ZN(n23186) );
  INV_X1 U16546 ( .A(n18585), .ZN(n23187) );
  INV_X1 U16547 ( .A(n18586), .ZN(n23188) );
  INV_X1 U16548 ( .A(n18586), .ZN(n23189) );
  INV_X1 U16549 ( .A(n27801), .ZN(n23190) );
  INV_X1 U16550 ( .A(n23190), .ZN(n23191) );
  INV_X1 U16551 ( .A(n23190), .ZN(n23192) );
  INV_X1 U16552 ( .A(n27228), .ZN(n23193) );
  INV_X1 U16553 ( .A(n23193), .ZN(n23194) );
  INV_X1 U16554 ( .A(n23193), .ZN(n23195) );
  INV_X1 U16555 ( .A(n18587), .ZN(n23196) );
  INV_X1 U16556 ( .A(n18587), .ZN(n23197) );
  INV_X1 U16557 ( .A(n18588), .ZN(n23198) );
  INV_X1 U16558 ( .A(n18588), .ZN(n23199) );
  INV_X1 U16559 ( .A(n18589), .ZN(n23200) );
  INV_X1 U16560 ( .A(n18589), .ZN(n23201) );
  INV_X1 U16561 ( .A(n26065), .ZN(n23202) );
  INV_X1 U16562 ( .A(n23202), .ZN(n23203) );
  INV_X1 U16563 ( .A(n23202), .ZN(n23204) );
  INV_X1 U16564 ( .A(n18590), .ZN(n23205) );
  INV_X1 U16565 ( .A(n18590), .ZN(n23206) );
  INV_X1 U16566 ( .A(n18591), .ZN(n23207) );
  INV_X1 U16567 ( .A(n18591), .ZN(n23208) );
  INV_X1 U16568 ( .A(n18592), .ZN(n23209) );
  INV_X1 U16569 ( .A(n18592), .ZN(n23210) );
  INV_X1 U16570 ( .A(n18593), .ZN(n23211) );
  INV_X1 U16571 ( .A(n26077), .ZN(n23212) );
  INV_X1 U16572 ( .A(n23212), .ZN(n23213) );
  INV_X1 U16573 ( .A(n23212), .ZN(n23214) );
  INV_X1 U16574 ( .A(n18594), .ZN(n23215) );
  INV_X1 U16575 ( .A(n18594), .ZN(n23216) );
  INV_X1 U16576 ( .A(n26669), .ZN(n23217) );
  INV_X1 U16577 ( .A(n24696), .ZN(n23218) );
  INV_X1 U16578 ( .A(n27273), .ZN(n23219) );
  INV_X1 U16579 ( .A(n26526), .ZN(n23220) );
  INV_X1 U16580 ( .A(n23220), .ZN(n23221) );
  INV_X1 U16581 ( .A(n23220), .ZN(n23222) );
  INV_X1 U16582 ( .A(n26091), .ZN(n23223) );
  INV_X1 U16583 ( .A(n23223), .ZN(n23224) );
  INV_X1 U16584 ( .A(n23223), .ZN(n23225) );
  INV_X1 U16585 ( .A(n18595), .ZN(n23226) );
  INV_X1 U16586 ( .A(n18596), .ZN(n23227) );
  INV_X1 U16587 ( .A(n18596), .ZN(n23228) );
  INV_X1 U16588 ( .A(n24694), .ZN(n23229) );
  INV_X1 U16589 ( .A(n27125), .ZN(n23230) );
  INV_X1 U16590 ( .A(n18597), .ZN(n23231) );
  INV_X1 U16591 ( .A(n18597), .ZN(n23232) );
  INV_X1 U16592 ( .A(n26102), .ZN(n23233) );
  INV_X1 U16593 ( .A(n23233), .ZN(n23234) );
  INV_X1 U16594 ( .A(n23233), .ZN(n23235) );
  INV_X1 U16595 ( .A(n18598), .ZN(n23236) );
  INV_X1 U16596 ( .A(n18598), .ZN(n23237) );
  INV_X1 U16597 ( .A(n18599), .ZN(n23238) );
  INV_X1 U16598 ( .A(n18599), .ZN(n23239) );
  INV_X1 U16599 ( .A(n26732), .ZN(n23240) );
  INV_X1 U16600 ( .A(n23240), .ZN(n23241) );
  INV_X1 U16601 ( .A(n23240), .ZN(n23242) );
  INV_X1 U16602 ( .A(n18600), .ZN(n23243) );
  INV_X1 U16603 ( .A(n18600), .ZN(n23244) );
  INV_X1 U16604 ( .A(n18601), .ZN(n23245) );
  INV_X1 U16605 ( .A(n18601), .ZN(n23246) );
  INV_X1 U16606 ( .A(n18602), .ZN(n23247) );
  INV_X1 U16607 ( .A(n18602), .ZN(n23248) );
  INV_X1 U16608 ( .A(n18603), .ZN(n23249) );
  INV_X1 U16609 ( .A(n18603), .ZN(n23250) );
  INV_X1 U16610 ( .A(n18604), .ZN(n23251) );
  INV_X1 U16611 ( .A(n18604), .ZN(n23252) );
  INV_X1 U16612 ( .A(n18605), .ZN(n23253) );
  INV_X1 U16613 ( .A(n18605), .ZN(n23254) );
  INV_X1 U16614 ( .A(n26739), .ZN(n23255) );
  INV_X1 U16615 ( .A(n23255), .ZN(n23256) );
  INV_X1 U16616 ( .A(n23255), .ZN(n23257) );
  INV_X1 U16617 ( .A(n18606), .ZN(n23258) );
  INV_X1 U16618 ( .A(n18606), .ZN(n23259) );
  INV_X1 U16619 ( .A(n18607), .ZN(n23260) );
  INV_X1 U16620 ( .A(n18607), .ZN(n23261) );
  INV_X1 U16621 ( .A(n18608), .ZN(n23262) );
  INV_X1 U16622 ( .A(n18608), .ZN(n23263) );
  INV_X1 U16623 ( .A(n26137), .ZN(n23264) );
  INV_X1 U16624 ( .A(n23264), .ZN(n23265) );
  INV_X1 U16625 ( .A(n23264), .ZN(n23266) );
  INV_X1 U16626 ( .A(n26138), .ZN(n23267) );
  INV_X1 U16627 ( .A(n23267), .ZN(n23268) );
  INV_X1 U16628 ( .A(n23267), .ZN(n23269) );
  INV_X1 U16629 ( .A(n18609), .ZN(n23270) );
  INV_X1 U16630 ( .A(n18609), .ZN(n23271) );
  INV_X1 U16631 ( .A(n26141), .ZN(n23272) );
  INV_X1 U16632 ( .A(n23272), .ZN(n23273) );
  INV_X1 U16633 ( .A(n23272), .ZN(n23274) );
  INV_X1 U16634 ( .A(n26142), .ZN(n23275) );
  INV_X1 U16635 ( .A(n23275), .ZN(n23276) );
  INV_X1 U16636 ( .A(n23275), .ZN(n23277) );
  INV_X1 U16637 ( .A(n18610), .ZN(n23278) );
  INV_X1 U16638 ( .A(n18611), .ZN(n23279) );
  INV_X1 U16639 ( .A(n18612), .ZN(n23280) );
  INV_X1 U16640 ( .A(n18612), .ZN(n23281) );
  INV_X1 U16641 ( .A(n18613), .ZN(n23282) );
  INV_X1 U16642 ( .A(n18613), .ZN(n23283) );
  INV_X1 U16643 ( .A(n25197), .ZN(n23284) );
  INV_X1 U16644 ( .A(n25197), .ZN(n23285) );
  INV_X1 U16645 ( .A(n18614), .ZN(n23286) );
  INV_X1 U16646 ( .A(n18614), .ZN(n23287) );
  INV_X1 U16647 ( .A(n18615), .ZN(n23288) );
  INV_X1 U16648 ( .A(n18615), .ZN(n23289) );
  INV_X1 U16649 ( .A(n18616), .ZN(n23290) );
  INV_X1 U16650 ( .A(n18616), .ZN(n23291) );
  INV_X1 U16651 ( .A(n18617), .ZN(n23292) );
  INV_X1 U16652 ( .A(n18617), .ZN(n23293) );
  INV_X1 U16653 ( .A(n18618), .ZN(n23294) );
  INV_X1 U16654 ( .A(n18618), .ZN(n23295) );
  INV_X1 U16655 ( .A(n25194), .ZN(n23296) );
  INV_X1 U16656 ( .A(n25194), .ZN(n23297) );
  INV_X1 U16657 ( .A(n18619), .ZN(n23298) );
  INV_X1 U16658 ( .A(n18619), .ZN(n23299) );
  INV_X1 U16659 ( .A(n102), .ZN(n23300) );
  INV_X1 U16660 ( .A(n102), .ZN(n23301) );
  INV_X1 U16661 ( .A(n18620), .ZN(n23302) );
  INV_X1 U16662 ( .A(n18620), .ZN(n23303) );
  INV_X1 U16663 ( .A(n101), .ZN(n23304) );
  INV_X1 U16664 ( .A(n101), .ZN(n23305) );
  INV_X1 U16665 ( .A(n100), .ZN(n23306) );
  INV_X1 U16666 ( .A(n100), .ZN(n23307) );
  INV_X1 U16667 ( .A(n26884), .ZN(n23308) );
  INV_X1 U16668 ( .A(n26884), .ZN(n23309) );
  INV_X1 U16669 ( .A(n99), .ZN(n23310) );
  INV_X1 U16670 ( .A(n99), .ZN(n23311) );
  INV_X1 U16671 ( .A(n26876), .ZN(n23312) );
  INV_X1 U16672 ( .A(n26876), .ZN(n23313) );
  INV_X1 U16673 ( .A(n268801), .ZN(n23314) );
  INV_X1 U16674 ( .A(n268801), .ZN(n23315) );
  INV_X1 U16675 ( .A(n1), .ZN(n23316) );
  INV_X1 U16676 ( .A(n1), .ZN(n23317) );
  INV_X1 U16677 ( .A(n26872), .ZN(n23318) );
  INV_X1 U16678 ( .A(n26872), .ZN(n23319) );
  INV_X1 U16679 ( .A(n26836), .ZN(n23320) );
  INV_X1 U16680 ( .A(n26827), .ZN(n23321) );
  INV_X1 U16681 ( .A(n2), .ZN(n23322) );
  INV_X1 U16682 ( .A(n2), .ZN(n23323) );
  INV_X1 U16683 ( .A(n98), .ZN(n23324) );
  INV_X1 U16684 ( .A(n98), .ZN(n23325) );
  INV_X1 U16685 ( .A(n67), .ZN(n23326) );
  INV_X1 U16686 ( .A(n67), .ZN(n23327) );
  INV_X1 U16687 ( .A(n97), .ZN(n23328) );
  INV_X1 U16688 ( .A(n97), .ZN(n23329) );
  INV_X1 U16689 ( .A(n96), .ZN(n23330) );
  INV_X1 U16690 ( .A(n96), .ZN(n23331) );
  INV_X1 U16691 ( .A(n27206), .ZN(n23332) );
  INV_X1 U16692 ( .A(n23332), .ZN(n23333) );
  INV_X1 U16693 ( .A(n23332), .ZN(n23334) );
  INV_X1 U16694 ( .A(n27205), .ZN(n23335) );
  INV_X1 U16695 ( .A(n23335), .ZN(n23336) );
  INV_X1 U16696 ( .A(n23335), .ZN(n23337) );
  INV_X1 U16697 ( .A(n27206), .ZN(n23338) );
  INV_X1 U16698 ( .A(n23338), .ZN(n23339) );
  INV_X1 U16699 ( .A(n23338), .ZN(n23340) );
  INV_X1 U16700 ( .A(n27205), .ZN(n23341) );
  INV_X1 U16701 ( .A(n23341), .ZN(n23342) );
  INV_X1 U16702 ( .A(n23341), .ZN(n23343) );
  INV_X1 U16703 ( .A(n95), .ZN(n23344) );
  INV_X1 U16704 ( .A(n95), .ZN(n23345) );
  INV_X1 U16705 ( .A(n94), .ZN(n23346) );
  INV_X1 U16706 ( .A(n94), .ZN(n23347) );
  INV_X1 U16707 ( .A(n93), .ZN(n23348) );
  INV_X1 U16708 ( .A(n93), .ZN(n23349) );
  INV_X1 U16709 ( .A(n92), .ZN(n23350) );
  INV_X1 U16710 ( .A(n92), .ZN(n23351) );
  INV_X1 U16711 ( .A(n91), .ZN(n23352) );
  INV_X1 U16712 ( .A(n91), .ZN(n23353) );
  INV_X1 U16713 ( .A(n90), .ZN(n23354) );
  INV_X1 U16714 ( .A(n90), .ZN(n23355) );
  INV_X1 U16715 ( .A(n89), .ZN(n23356) );
  INV_X1 U16716 ( .A(n89), .ZN(n23357) );
  INV_X1 U16717 ( .A(n88), .ZN(n23358) );
  INV_X1 U16718 ( .A(n88), .ZN(n23359) );
  INV_X1 U16719 ( .A(n87), .ZN(n23360) );
  INV_X1 U16720 ( .A(n87), .ZN(n23361) );
  INV_X1 U16721 ( .A(n86), .ZN(n23362) );
  INV_X1 U16722 ( .A(n86), .ZN(n23363) );
  INV_X1 U16723 ( .A(n85), .ZN(n23364) );
  INV_X1 U16724 ( .A(n85), .ZN(n23365) );
  INV_X1 U16725 ( .A(n84), .ZN(n23366) );
  INV_X1 U16726 ( .A(n84), .ZN(n23367) );
  INV_X1 U16727 ( .A(n83), .ZN(n23368) );
  INV_X1 U16728 ( .A(n83), .ZN(n23369) );
  INV_X1 U16729 ( .A(n82), .ZN(n23370) );
  INV_X1 U16730 ( .A(n82), .ZN(n23371) );
  INV_X1 U16731 ( .A(n81), .ZN(n23372) );
  INV_X1 U16732 ( .A(n81), .ZN(n23373) );
  INV_X1 U16733 ( .A(n80), .ZN(n23374) );
  INV_X1 U16734 ( .A(n80), .ZN(n23375) );
  INV_X1 U16735 ( .A(n277401), .ZN(n23376) );
  INV_X1 U16736 ( .A(n23376), .ZN(n23377) );
  INV_X1 U16737 ( .A(n23376), .ZN(n23378) );
  INV_X1 U16738 ( .A(n26246), .ZN(n23379) );
  INV_X1 U16739 ( .A(n23379), .ZN(n23380) );
  INV_X1 U16740 ( .A(n23379), .ZN(n23381) );
  INV_X1 U16741 ( .A(n24874), .ZN(n23382) );
  INV_X1 U16742 ( .A(n23382), .ZN(n23383) );
  INV_X1 U16743 ( .A(n23382), .ZN(n23384) );
  INV_X1 U16744 ( .A(n18621), .ZN(n23385) );
  INV_X1 U16745 ( .A(n18621), .ZN(n23386) );
  INV_X1 U16746 ( .A(n27171), .ZN(n23387) );
  INV_X1 U16747 ( .A(n23387), .ZN(n23388) );
  INV_X1 U16748 ( .A(n23387), .ZN(n23389) );
  INV_X1 U16749 ( .A(n18622), .ZN(n23390) );
  INV_X1 U16750 ( .A(n18622), .ZN(n23391) );
  INV_X1 U16751 ( .A(n18623), .ZN(n23392) );
  INV_X1 U16752 ( .A(n18623), .ZN(n23393) );
  INV_X1 U16753 ( .A(n26263), .ZN(n23394) );
  INV_X1 U16754 ( .A(n23394), .ZN(n23395) );
  INV_X1 U16755 ( .A(n23394), .ZN(n23396) );
  INV_X1 U16756 ( .A(n24879), .ZN(n23397) );
  INV_X1 U16757 ( .A(n23397), .ZN(n23398) );
  INV_X1 U16758 ( .A(n23397), .ZN(n23399) );
  INV_X1 U16759 ( .A(n18624), .ZN(n23400) );
  INV_X1 U16760 ( .A(n18624), .ZN(n23401) );
  INV_X1 U16761 ( .A(n23673), .ZN(n23402) );
  INV_X1 U16762 ( .A(n23402), .ZN(n23403) );
  INV_X1 U16763 ( .A(n23402), .ZN(n23404) );
  INV_X1 U16764 ( .A(n18625), .ZN(n23405) );
  INV_X1 U16765 ( .A(n18625), .ZN(n23406) );
  INV_X1 U16766 ( .A(n18626), .ZN(n23407) );
  INV_X1 U16767 ( .A(n18626), .ZN(n23408) );
  INV_X1 U16768 ( .A(n27259), .ZN(n23409) );
  INV_X1 U16769 ( .A(n23409), .ZN(n23410) );
  INV_X1 U16770 ( .A(n23409), .ZN(n23411) );
  INV_X1 U16771 ( .A(n18627), .ZN(n23412) );
  INV_X1 U16772 ( .A(n18627), .ZN(n23413) );
  INV_X1 U16773 ( .A(n18628), .ZN(n23414) );
  INV_X1 U16774 ( .A(n18628), .ZN(n23415) );
  INV_X1 U16775 ( .A(n26288), .ZN(n23416) );
  INV_X1 U16776 ( .A(n23416), .ZN(n23417) );
  INV_X1 U16777 ( .A(n23416), .ZN(n23418) );
  INV_X1 U16778 ( .A(n18629), .ZN(n23419) );
  INV_X1 U16779 ( .A(n18629), .ZN(n23420) );
  INV_X1 U16780 ( .A(n18630), .ZN(n23421) );
  INV_X1 U16781 ( .A(n18630), .ZN(n23422) );
  INV_X1 U16782 ( .A(n26297), .ZN(n23423) );
  INV_X1 U16783 ( .A(n23423), .ZN(n23424) );
  INV_X1 U16784 ( .A(n18631), .ZN(n23425) );
  INV_X1 U16785 ( .A(n18631), .ZN(n23426) );
  INV_X1 U16786 ( .A(n18632), .ZN(n23427) );
  INV_X1 U16787 ( .A(n18632), .ZN(n23428) );
  INV_X1 U16788 ( .A(n18633), .ZN(n23429) );
  INV_X1 U16789 ( .A(n18633), .ZN(n23430) );
  INV_X1 U16790 ( .A(n18634), .ZN(n23431) );
  INV_X1 U16791 ( .A(n18634), .ZN(n23432) );
  INV_X1 U16792 ( .A(n18635), .ZN(n23433) );
  INV_X1 U16793 ( .A(n18635), .ZN(n23434) );
  INV_X1 U16794 ( .A(n18636), .ZN(n23435) );
  INV_X1 U16795 ( .A(n18636), .ZN(n23436) );
  INV_X1 U16796 ( .A(n18637), .ZN(n23437) );
  INV_X1 U16797 ( .A(n18637), .ZN(n23438) );
  INV_X1 U16798 ( .A(n18638), .ZN(n23439) );
  INV_X1 U16799 ( .A(n18638), .ZN(n23440) );
  INV_X1 U16800 ( .A(n18639), .ZN(n23441) );
  INV_X1 U16801 ( .A(n18639), .ZN(n23442) );
  INV_X1 U16802 ( .A(n36250), .ZN(n23443) );
  INV_X1 U16803 ( .A(n32110), .ZN(n23444) );
  INV_X1 U16804 ( .A(n18986), .ZN(n23445) );
  INV_X1 U16805 ( .A(n17135), .ZN(n23446) );
  INV_X1 U16806 ( .A(n17134), .ZN(n23447) );
  INV_X1 U16807 ( .A(n26644), .ZN(n23448) );
  INV_X1 U16808 ( .A(n26329), .ZN(n23449) );
  INV_X1 U16809 ( .A(n23449), .ZN(n23450) );
  INV_X1 U16810 ( .A(n23449), .ZN(n23451) );
  INV_X1 U16811 ( .A(n27045), .ZN(n23452) );
  INV_X1 U16812 ( .A(n27045), .ZN(n23453) );
  INV_X1 U16813 ( .A(n27046), .ZN(n23454) );
  INV_X1 U16814 ( .A(n27046), .ZN(n23455) );
  INV_X1 U16815 ( .A(n18640), .ZN(n23456) );
  INV_X1 U16816 ( .A(n18640), .ZN(n23457) );
  INV_X1 U16817 ( .A(n27044), .ZN(n23458) );
  INV_X1 U16818 ( .A(n27044), .ZN(n23459) );
  INV_X1 U16819 ( .A(n18641), .ZN(n23460) );
  INV_X1 U16820 ( .A(n18641), .ZN(n23461) );
  INV_X1 U16821 ( .A(n18642), .ZN(n23462) );
  INV_X1 U16822 ( .A(n18642), .ZN(n23463) );
  INV_X1 U16823 ( .A(n18643), .ZN(n23464) );
  INV_X1 U16824 ( .A(n18643), .ZN(n23465) );
  INV_X1 U16825 ( .A(n18644), .ZN(n23466) );
  INV_X1 U16826 ( .A(n18644), .ZN(n23467) );
  INV_X1 U16827 ( .A(n18645), .ZN(n23468) );
  INV_X1 U16828 ( .A(n18645), .ZN(n23469) );
  INV_X1 U16829 ( .A(n18646), .ZN(n23470) );
  INV_X1 U16830 ( .A(n18646), .ZN(n23471) );
  INV_X1 U16831 ( .A(n18647), .ZN(n23472) );
  INV_X1 U16832 ( .A(n18647), .ZN(n23473) );
  INV_X1 U16833 ( .A(n18648), .ZN(n23474) );
  INV_X1 U16834 ( .A(n18648), .ZN(n23475) );
  INV_X1 U16835 ( .A(n26996), .ZN(n23476) );
  INV_X1 U16836 ( .A(n26996), .ZN(n23477) );
  INV_X1 U16837 ( .A(n18649), .ZN(n23478) );
  INV_X1 U16838 ( .A(n18649), .ZN(n23479) );
  INV_X1 U16839 ( .A(n18650), .ZN(n23480) );
  INV_X1 U16840 ( .A(n18650), .ZN(n23481) );
  INV_X1 U16841 ( .A(n26995), .ZN(n23482) );
  INV_X1 U16842 ( .A(n26995), .ZN(n23483) );
  INV_X1 U16843 ( .A(n25207), .ZN(n23484) );
  INV_X1 U16844 ( .A(n23484), .ZN(n23485) );
  INV_X1 U16845 ( .A(n23484), .ZN(n23486) );
  INV_X1 U16846 ( .A(n18651), .ZN(n23487) );
  INV_X1 U16847 ( .A(n18651), .ZN(n23488) );
  INV_X1 U16848 ( .A(n25219), .ZN(n23489) );
  INV_X1 U16849 ( .A(n23489), .ZN(n23490) );
  INV_X1 U16850 ( .A(n23489), .ZN(n23491) );
  INV_X1 U16851 ( .A(n18652), .ZN(n23492) );
  INV_X1 U16852 ( .A(n18652), .ZN(n23493) );
  INV_X1 U16853 ( .A(n18653), .ZN(n23494) );
  INV_X1 U16854 ( .A(n18653), .ZN(n23495) );
  INV_X1 U16855 ( .A(n18654), .ZN(n23496) );
  INV_X1 U16856 ( .A(n18654), .ZN(n23497) );
  INV_X1 U16857 ( .A(n18655), .ZN(n23498) );
  INV_X1 U16858 ( .A(n18655), .ZN(n23499) );
  INV_X1 U16859 ( .A(n17109), .ZN(n23500) );
  INV_X1 U16860 ( .A(n17109), .ZN(n23501) );
  INV_X1 U16861 ( .A(n17108), .ZN(n23502) );
  INV_X1 U16862 ( .A(n17108), .ZN(n23503) );
  INV_X1 U16863 ( .A(n17107), .ZN(n23504) );
  INV_X1 U16864 ( .A(n17107), .ZN(n23505) );
  INV_X1 U16865 ( .A(n17106), .ZN(n23506) );
  INV_X1 U16866 ( .A(n17106), .ZN(n23507) );
  INV_X1 U16867 ( .A(n18656), .ZN(n23508) );
  INV_X1 U16868 ( .A(n18656), .ZN(n23509) );
  INV_X1 U16869 ( .A(n18657), .ZN(n23510) );
  INV_X1 U16870 ( .A(n18657), .ZN(n23511) );
  INV_X1 U16871 ( .A(n18658), .ZN(n23512) );
  INV_X1 U16872 ( .A(n18658), .ZN(n23513) );
  INV_X1 U16873 ( .A(n18659), .ZN(n23514) );
  INV_X1 U16874 ( .A(n18659), .ZN(n23515) );
  INV_X1 U16875 ( .A(n18660), .ZN(n23516) );
  INV_X1 U16876 ( .A(n18660), .ZN(n23517) );
  INV_X1 U16877 ( .A(n18661), .ZN(n23518) );
  INV_X1 U16878 ( .A(n18661), .ZN(n23519) );
  INV_X1 U16879 ( .A(n18662), .ZN(n23520) );
  INV_X1 U16880 ( .A(n18662), .ZN(n23521) );
  INV_X1 U16881 ( .A(n18663), .ZN(n23522) );
  INV_X1 U16882 ( .A(n18663), .ZN(n23523) );
  INV_X1 U16883 ( .A(n26882), .ZN(n23524) );
  INV_X1 U16884 ( .A(n26882), .ZN(n23525) );
  INV_X1 U16885 ( .A(n26883), .ZN(n23526) );
  INV_X1 U16886 ( .A(n26883), .ZN(n23527) );
  INV_X1 U16887 ( .A(n26879), .ZN(n23528) );
  INV_X1 U16888 ( .A(n26879), .ZN(n23529) );
  INV_X1 U16889 ( .A(n26881), .ZN(n23530) );
  INV_X1 U16890 ( .A(n26881), .ZN(n23531) );
  INV_X1 U16891 ( .A(n26877), .ZN(n23532) );
  INV_X1 U16892 ( .A(n26877), .ZN(n23533) );
  INV_X1 U16893 ( .A(n26878), .ZN(n23534) );
  INV_X1 U16894 ( .A(n26878), .ZN(n23535) );
  INV_X1 U16895 ( .A(n26874), .ZN(n23536) );
  INV_X1 U16896 ( .A(n26874), .ZN(n23537) );
  INV_X1 U16897 ( .A(n26875), .ZN(n23538) );
  INV_X1 U16898 ( .A(n26875), .ZN(n23539) );
  INV_X1 U16899 ( .A(n26871), .ZN(n23540) );
  INV_X1 U16900 ( .A(n26871), .ZN(n23541) );
  INV_X1 U16901 ( .A(n26873), .ZN(n23542) );
  INV_X1 U16902 ( .A(n26873), .ZN(n23543) );
  INV_X1 U16903 ( .A(n26869), .ZN(n23544) );
  INV_X1 U16904 ( .A(n26869), .ZN(n23545) );
  INV_X1 U16905 ( .A(n268701), .ZN(n23546) );
  INV_X1 U16906 ( .A(n268701), .ZN(n23547) );
  INV_X1 U16907 ( .A(n26835), .ZN(n23548) );
  INV_X1 U16908 ( .A(n268401), .ZN(n23549) );
  INV_X1 U16909 ( .A(n18664), .ZN(n23550) );
  INV_X1 U16910 ( .A(n26868), .ZN(n23551) );
  INV_X1 U16911 ( .A(n26868), .ZN(n23552) );
  INV_X1 U16912 ( .A(n18863), .ZN(n23553) );
  INV_X1 U16913 ( .A(n26833), .ZN(n23554) );
  INV_X1 U16914 ( .A(n26825), .ZN(n23555) );
  INV_X1 U16915 ( .A(n18665), .ZN(n23556) );
  INV_X1 U16916 ( .A(n18665), .ZN(n23557) );
  INV_X1 U16917 ( .A(n18666), .ZN(n23558) );
  INV_X1 U16918 ( .A(n26834), .ZN(n23559) );
  INV_X1 U16919 ( .A(n26838), .ZN(n23560) );
  INV_X1 U16920 ( .A(n18667), .ZN(n23561) );
  INV_X1 U16921 ( .A(n26837), .ZN(n23562) );
  INV_X1 U16922 ( .A(n268301), .ZN(n23563) );
  INV_X1 U16923 ( .A(n18668), .ZN(n23564) );
  INV_X1 U16924 ( .A(n18668), .ZN(n23565) );
  INV_X1 U16925 ( .A(n18669), .ZN(n23566) );
  INV_X1 U16926 ( .A(n18669), .ZN(n23567) );
  INV_X1 U16927 ( .A(n18670), .ZN(n23568) );
  INV_X1 U16928 ( .A(n18670), .ZN(n23569) );
  INV_X1 U16929 ( .A(n18671), .ZN(n23570) );
  INV_X1 U16930 ( .A(n18671), .ZN(n23571) );
  INV_X1 U16931 ( .A(n18672), .ZN(n23572) );
  INV_X1 U16932 ( .A(n18672), .ZN(n23573) );
  INV_X1 U16933 ( .A(n18673), .ZN(n23574) );
  INV_X1 U16934 ( .A(n18673), .ZN(n23575) );
  INV_X1 U16935 ( .A(n18674), .ZN(n23576) );
  INV_X1 U16936 ( .A(n18674), .ZN(n23577) );
  INV_X1 U16937 ( .A(n18675), .ZN(n23578) );
  INV_X1 U16938 ( .A(n18675), .ZN(n23579) );
  INV_X1 U16939 ( .A(n18676), .ZN(n23580) );
  INV_X1 U16940 ( .A(n18676), .ZN(n23581) );
  INV_X1 U16941 ( .A(n18677), .ZN(n23582) );
  INV_X1 U16942 ( .A(n18677), .ZN(n23583) );
  INV_X1 U16943 ( .A(n27121), .ZN(n23584) );
  INV_X1 U16944 ( .A(n23584), .ZN(n23585) );
  INV_X1 U16945 ( .A(n23584), .ZN(n23586) );
  INV_X1 U16946 ( .A(n18678), .ZN(n23587) );
  INV_X1 U16947 ( .A(n26856), .ZN(n23588) );
  INV_X1 U16948 ( .A(n18679), .ZN(n23589) );
  INV_X1 U16949 ( .A(n18679), .ZN(n23590) );
  INV_X1 U16950 ( .A(n18680), .ZN(n23591) );
  INV_X1 U16951 ( .A(n18680), .ZN(n23592) );
  INV_X1 U16952 ( .A(n18681), .ZN(n23593) );
  INV_X1 U16953 ( .A(n18681), .ZN(n23594) );
  INV_X1 U16954 ( .A(n18682), .ZN(n23595) );
  INV_X1 U16955 ( .A(n18682), .ZN(n23596) );
  INV_X1 U16956 ( .A(n18683), .ZN(n23597) );
  INV_X1 U16957 ( .A(n18683), .ZN(n23598) );
  INV_X1 U16958 ( .A(n18684), .ZN(n23599) );
  INV_X1 U16959 ( .A(n18684), .ZN(n23600) );
  INV_X1 U16960 ( .A(n18685), .ZN(n23601) );
  INV_X1 U16961 ( .A(n18685), .ZN(n23602) );
  INV_X1 U16962 ( .A(n18686), .ZN(n23603) );
  INV_X1 U16963 ( .A(n18686), .ZN(n23604) );
  INV_X1 U16964 ( .A(n18687), .ZN(n23605) );
  INV_X1 U16965 ( .A(n18687), .ZN(n23606) );
  INV_X1 U16966 ( .A(n18688), .ZN(n23607) );
  INV_X1 U16967 ( .A(n18688), .ZN(n23608) );
  INV_X1 U16968 ( .A(n18689), .ZN(n23609) );
  INV_X1 U16969 ( .A(n18689), .ZN(n23610) );
  INV_X1 U16970 ( .A(n18690), .ZN(n23611) );
  INV_X1 U16971 ( .A(n18690), .ZN(n23612) );
  INV_X1 U16972 ( .A(n18691), .ZN(n23613) );
  INV_X1 U16973 ( .A(n18691), .ZN(n23614) );
  INV_X1 U16974 ( .A(n18692), .ZN(n23615) );
  INV_X1 U16975 ( .A(n18692), .ZN(n23616) );
  INV_X1 U16976 ( .A(n18693), .ZN(n23617) );
  INV_X1 U16977 ( .A(n18693), .ZN(n23618) );
  INV_X1 U16978 ( .A(n18694), .ZN(n23619) );
  INV_X1 U16979 ( .A(n18694), .ZN(n23620) );
  INV_X1 U16980 ( .A(n18695), .ZN(n23621) );
  INV_X1 U16981 ( .A(n18695), .ZN(n23622) );
  INV_X1 U16982 ( .A(n18696), .ZN(n23623) );
  INV_X1 U16983 ( .A(n18696), .ZN(n23624) );
  INV_X1 U16984 ( .A(n18697), .ZN(n23625) );
  INV_X1 U16985 ( .A(n18697), .ZN(n23626) );
  INV_X1 U16986 ( .A(n18698), .ZN(n23627) );
  INV_X1 U16987 ( .A(n18698), .ZN(n23628) );
  INV_X1 U16988 ( .A(n18699), .ZN(n23629) );
  INV_X1 U16989 ( .A(n18699), .ZN(n23630) );
  INV_X1 U16990 ( .A(n18700), .ZN(n23631) );
  INV_X1 U16991 ( .A(n18700), .ZN(n23632) );
  INV_X1 U16992 ( .A(n18701), .ZN(n23633) );
  INV_X1 U16993 ( .A(n18701), .ZN(n23634) );
  INV_X1 U16994 ( .A(n18702), .ZN(n23635) );
  INV_X1 U16995 ( .A(n18702), .ZN(n23636) );
  INV_X1 U16996 ( .A(n18703), .ZN(n23637) );
  INV_X1 U16997 ( .A(n18703), .ZN(n23638) );
  INV_X1 U16998 ( .A(n4979), .ZN(n23639) );
  INV_X1 U16999 ( .A(n4979), .ZN(n23640) );
  INV_X1 U17000 ( .A(n23377), .ZN(n23641) );
  INV_X1 U17001 ( .A(n22428), .ZN(n23642) );
  INV_X1 U17002 ( .A(n26513), .ZN(n23643) );
  INV_X1 U17003 ( .A(n23643), .ZN(n23644) );
  INV_X1 U17004 ( .A(n23643), .ZN(n23645) );
  INV_X1 U17005 ( .A(r899_B_1_), .ZN(n23646) );
  INV_X1 U17006 ( .A(r899_B_1_), .ZN(n23647) );
  INV_X1 U17007 ( .A(n17134), .ZN(n23648) );
  INV_X1 U17008 ( .A(n17135), .ZN(n23649) );
  INV_X1 U17009 ( .A(n26321), .ZN(n23650) );
  INV_X1 U17010 ( .A(n23650), .ZN(n23651) );
  INV_X1 U17011 ( .A(n18704), .ZN(n23652) );
  INV_X1 U17012 ( .A(n18704), .ZN(n23653) );
  INV_X1 U17013 ( .A(n265201), .ZN(n23654) );
  INV_X1 U17014 ( .A(n23654), .ZN(n23655) );
  INV_X1 U17015 ( .A(n23654), .ZN(n23656) );
  INV_X1 U17016 ( .A(n25644), .ZN(n23657) );
  INV_X1 U17017 ( .A(n23657), .ZN(n23658) );
  INV_X1 U17018 ( .A(n26526), .ZN(n23659) );
  INV_X1 U17019 ( .A(n23659), .ZN(n23660) );
  INV_X1 U17020 ( .A(n23659), .ZN(n23661) );
  INV_X1 U17021 ( .A(n26531), .ZN(n23662) );
  INV_X1 U17022 ( .A(n23662), .ZN(n23663) );
  INV_X1 U17023 ( .A(n23662), .ZN(n23664) );
  INV_X1 U17024 ( .A(n18705), .ZN(n23665) );
  INV_X1 U17025 ( .A(n18706), .ZN(n23666) );
  INV_X1 U17026 ( .A(n18707), .ZN(n23667) );
  INV_X1 U17027 ( .A(n18707), .ZN(n23668) );
  INV_X1 U17028 ( .A(n18708), .ZN(n23669) );
  INV_X1 U17029 ( .A(n18708), .ZN(n23670) );
  INV_X1 U17030 ( .A(n24698), .ZN(n23671) );
  INV_X1 U17031 ( .A(n23671), .ZN(n23672) );
  INV_X1 U17032 ( .A(n23671), .ZN(n23673) );
  INV_X1 U17033 ( .A(n18709), .ZN(n23674) );
  INV_X1 U17034 ( .A(n18709), .ZN(n23675) );
  INV_X1 U17035 ( .A(n26549), .ZN(n23676) );
  INV_X1 U17036 ( .A(n23676), .ZN(n23677) );
  INV_X1 U17037 ( .A(n23676), .ZN(n23678) );
  INV_X1 U17038 ( .A(n23678), .ZN(n23679) );
  INV_X1 U17039 ( .A(n23678), .ZN(n23680) );
  INV_X1 U17040 ( .A(n26552), .ZN(n23681) );
  INV_X1 U17041 ( .A(n23681), .ZN(n23682) );
  INV_X1 U17042 ( .A(n23681), .ZN(n23683) );
  INV_X1 U17043 ( .A(n26553), .ZN(n23684) );
  INV_X1 U17044 ( .A(n23684), .ZN(n23685) );
  INV_X1 U17045 ( .A(n23684), .ZN(n23686) );
  INV_X1 U17046 ( .A(n18710), .ZN(n23687) );
  INV_X1 U17047 ( .A(n18710), .ZN(n23688) );
  INV_X1 U17048 ( .A(n26558), .ZN(n23689) );
  INV_X1 U17049 ( .A(n23689), .ZN(n23690) );
  INV_X1 U17050 ( .A(n23689), .ZN(n23691) );
  INV_X1 U17051 ( .A(n18711), .ZN(n23692) );
  INV_X1 U17052 ( .A(n18711), .ZN(n23693) );
  INV_X1 U17053 ( .A(n26564), .ZN(n23694) );
  INV_X1 U17054 ( .A(n23694), .ZN(n23695) );
  INV_X1 U17055 ( .A(n23694), .ZN(n23696) );
  INV_X1 U17056 ( .A(n18712), .ZN(n23697) );
  INV_X1 U17057 ( .A(n18712), .ZN(n23698) );
  INV_X1 U17058 ( .A(n26568), .ZN(n23699) );
  INV_X1 U17059 ( .A(n23699), .ZN(n23700) );
  INV_X1 U17060 ( .A(n23699), .ZN(n23701) );
  INV_X1 U17061 ( .A(n18713), .ZN(n23702) );
  INV_X1 U17062 ( .A(n18713), .ZN(n23703) );
  INV_X1 U17063 ( .A(n26572), .ZN(n23704) );
  INV_X1 U17064 ( .A(n23704), .ZN(n23705) );
  INV_X1 U17065 ( .A(n23704), .ZN(n23706) );
  INV_X1 U17066 ( .A(n18714), .ZN(n23707) );
  INV_X1 U17067 ( .A(n18714), .ZN(n23708) );
  INV_X1 U17068 ( .A(n26577), .ZN(n23709) );
  INV_X1 U17069 ( .A(n23709), .ZN(n23710) );
  INV_X1 U17070 ( .A(n23709), .ZN(n23711) );
  INV_X1 U17071 ( .A(n18715), .ZN(n23712) );
  INV_X1 U17072 ( .A(n18715), .ZN(n23713) );
  INV_X1 U17073 ( .A(n26581), .ZN(n23714) );
  INV_X1 U17074 ( .A(n23714), .ZN(n23715) );
  INV_X1 U17075 ( .A(n23714), .ZN(n23716) );
  INV_X1 U17076 ( .A(n18716), .ZN(n23717) );
  INV_X1 U17077 ( .A(n18716), .ZN(n23718) );
  INV_X1 U17078 ( .A(n26583), .ZN(n23719) );
  INV_X1 U17079 ( .A(n23719), .ZN(n23720) );
  INV_X1 U17080 ( .A(n23719), .ZN(n23721) );
  INV_X1 U17081 ( .A(n18717), .ZN(n23722) );
  INV_X1 U17082 ( .A(n18717), .ZN(n23723) );
  INV_X1 U17083 ( .A(n26586), .ZN(n23724) );
  INV_X1 U17084 ( .A(n23724), .ZN(n23725) );
  INV_X1 U17085 ( .A(n23724), .ZN(n23726) );
  INV_X1 U17086 ( .A(n25515), .ZN(n23727) );
  INV_X1 U17087 ( .A(n23727), .ZN(n23728) );
  INV_X1 U17088 ( .A(n23727), .ZN(n23729) );
  INV_X1 U17089 ( .A(n18718), .ZN(n23730) );
  INV_X1 U17090 ( .A(n18718), .ZN(n23731) );
  INV_X1 U17091 ( .A(n18719), .ZN(n23732) );
  INV_X1 U17092 ( .A(n18719), .ZN(n23733) );
  INV_X1 U17093 ( .A(n26595), .ZN(n23734) );
  INV_X1 U17094 ( .A(n23734), .ZN(n23735) );
  INV_X1 U17095 ( .A(n23734), .ZN(n23736) );
  INV_X1 U17096 ( .A(n26593), .ZN(n23737) );
  INV_X1 U17097 ( .A(n23737), .ZN(n23738) );
  INV_X1 U17098 ( .A(n23737), .ZN(n23739) );
  INV_X1 U17099 ( .A(n19271), .ZN(n23740) );
  INV_X1 U17100 ( .A(n23740), .ZN(n23741) );
  INV_X1 U17101 ( .A(n23740), .ZN(n23742) );
  INV_X1 U17102 ( .A(n18722), .ZN(n23743) );
  INV_X1 U17103 ( .A(n18722), .ZN(n23744) );
  INV_X1 U17104 ( .A(n18723), .ZN(n23745) );
  INV_X1 U17105 ( .A(n18723), .ZN(n23746) );
  INV_X1 U17106 ( .A(n18724), .ZN(n23747) );
  INV_X1 U17107 ( .A(n18724), .ZN(n23748) );
  INV_X1 U17108 ( .A(n18725), .ZN(n23749) );
  INV_X1 U17109 ( .A(n18725), .ZN(n23750) );
  INV_X1 U17110 ( .A(n18726), .ZN(n23751) );
  INV_X1 U17111 ( .A(n18726), .ZN(n23752) );
  INV_X1 U17112 ( .A(n18727), .ZN(n23753) );
  INV_X1 U17113 ( .A(n18727), .ZN(n23754) );
  INV_X1 U17114 ( .A(n18728), .ZN(n23755) );
  INV_X1 U17115 ( .A(n18728), .ZN(n23756) );
  INV_X1 U17116 ( .A(n18729), .ZN(n23757) );
  INV_X1 U17117 ( .A(n18729), .ZN(n23758) );
  INV_X1 U17118 ( .A(n18730), .ZN(n23759) );
  INV_X1 U17119 ( .A(n18730), .ZN(n23760) );
  INV_X1 U17120 ( .A(n18731), .ZN(n23761) );
  INV_X1 U17121 ( .A(n18731), .ZN(n23762) );
  INV_X1 U17122 ( .A(n18732), .ZN(n23763) );
  INV_X1 U17123 ( .A(n18732), .ZN(n23764) );
  INV_X1 U17124 ( .A(n18733), .ZN(n23765) );
  INV_X1 U17125 ( .A(n18733), .ZN(n23766) );
  INV_X1 U17126 ( .A(n18734), .ZN(n23767) );
  INV_X1 U17127 ( .A(n18734), .ZN(n23768) );
  INV_X1 U17128 ( .A(n18735), .ZN(n23769) );
  INV_X1 U17129 ( .A(n18735), .ZN(n23770) );
  INV_X1 U17130 ( .A(n18736), .ZN(n23771) );
  INV_X1 U17131 ( .A(n18736), .ZN(n23772) );
  INV_X1 U17132 ( .A(n18737), .ZN(n23773) );
  INV_X1 U17133 ( .A(n18737), .ZN(n23774) );
  INV_X1 U17134 ( .A(n18738), .ZN(n23775) );
  INV_X1 U17135 ( .A(n18738), .ZN(n23776) );
  INV_X1 U17136 ( .A(n18739), .ZN(n23777) );
  INV_X1 U17137 ( .A(n18739), .ZN(n23778) );
  INV_X1 U17138 ( .A(n18740), .ZN(n23779) );
  INV_X1 U17139 ( .A(n18740), .ZN(n23780) );
  INV_X1 U17140 ( .A(n18741), .ZN(n23781) );
  INV_X1 U17141 ( .A(n18741), .ZN(n23782) );
  INV_X1 U17142 ( .A(n18742), .ZN(n23783) );
  INV_X1 U17143 ( .A(n18742), .ZN(n23784) );
  INV_X1 U17144 ( .A(n18743), .ZN(n23785) );
  INV_X1 U17145 ( .A(n18743), .ZN(n23786) );
  INV_X1 U17146 ( .A(n18744), .ZN(n23787) );
  INV_X1 U17147 ( .A(n18744), .ZN(n23788) );
  INV_X1 U17148 ( .A(n18745), .ZN(n23789) );
  INV_X1 U17149 ( .A(n18745), .ZN(n23790) );
  INV_X1 U17150 ( .A(n18746), .ZN(n23791) );
  INV_X1 U17151 ( .A(n18746), .ZN(n23792) );
  INV_X1 U17152 ( .A(n18747), .ZN(n23793) );
  INV_X1 U17153 ( .A(n18747), .ZN(n23794) );
  INV_X1 U17154 ( .A(n18748), .ZN(n23795) );
  INV_X1 U17155 ( .A(n18748), .ZN(n23796) );
  INV_X1 U17156 ( .A(n18749), .ZN(n23797) );
  INV_X1 U17157 ( .A(n18749), .ZN(n23798) );
  INV_X1 U17158 ( .A(n18750), .ZN(n23799) );
  INV_X1 U17159 ( .A(n18750), .ZN(n23800) );
  INV_X1 U17160 ( .A(n18751), .ZN(n23801) );
  INV_X1 U17161 ( .A(n18751), .ZN(n23802) );
  INV_X1 U17162 ( .A(n18752), .ZN(n23803) );
  INV_X1 U17163 ( .A(n18752), .ZN(n23804) );
  INV_X1 U17164 ( .A(n18753), .ZN(n23805) );
  INV_X1 U17165 ( .A(n18753), .ZN(n23806) );
  INV_X1 U17166 ( .A(n18754), .ZN(n23807) );
  INV_X1 U17167 ( .A(n18754), .ZN(n23808) );
  INV_X1 U17168 ( .A(n18755), .ZN(n23809) );
  INV_X1 U17169 ( .A(n18755), .ZN(n23810) );
  INV_X1 U17170 ( .A(n18756), .ZN(n23811) );
  INV_X1 U17171 ( .A(n18756), .ZN(n23812) );
  INV_X1 U17172 ( .A(n18757), .ZN(n23813) );
  INV_X1 U17173 ( .A(n18757), .ZN(n23814) );
  INV_X1 U17174 ( .A(n18758), .ZN(n23815) );
  INV_X1 U17175 ( .A(n18758), .ZN(n23816) );
  INV_X1 U17176 ( .A(n18759), .ZN(n23817) );
  INV_X1 U17177 ( .A(n18759), .ZN(n23818) );
  INV_X1 U17178 ( .A(n18760), .ZN(n23819) );
  INV_X1 U17179 ( .A(n18760), .ZN(n23820) );
  INV_X1 U17180 ( .A(n18761), .ZN(n23821) );
  INV_X1 U17181 ( .A(n18761), .ZN(n23822) );
  INV_X1 U17182 ( .A(n18762), .ZN(n23823) );
  INV_X1 U17183 ( .A(n18762), .ZN(n23824) );
  INV_X1 U17184 ( .A(n18763), .ZN(n23825) );
  INV_X1 U17185 ( .A(n18763), .ZN(n23826) );
  INV_X1 U17186 ( .A(n18764), .ZN(n23827) );
  INV_X1 U17187 ( .A(n18764), .ZN(n23828) );
  INV_X1 U17188 ( .A(n18765), .ZN(n23829) );
  INV_X1 U17189 ( .A(n18765), .ZN(n23830) );
  INV_X1 U17190 ( .A(n18766), .ZN(n23831) );
  INV_X1 U17191 ( .A(n18766), .ZN(n23832) );
  INV_X1 U17192 ( .A(n18767), .ZN(n23833) );
  INV_X1 U17193 ( .A(n18767), .ZN(n23834) );
  INV_X1 U17194 ( .A(n18768), .ZN(n23835) );
  INV_X1 U17195 ( .A(n18768), .ZN(n23836) );
  INV_X1 U17196 ( .A(n18769), .ZN(n23837) );
  INV_X1 U17197 ( .A(n18769), .ZN(n23838) );
  INV_X1 U17198 ( .A(n18770), .ZN(n23839) );
  INV_X1 U17199 ( .A(n18770), .ZN(n23840) );
  INV_X1 U17200 ( .A(n18771), .ZN(n23841) );
  INV_X1 U17201 ( .A(n18771), .ZN(n23842) );
  INV_X1 U17202 ( .A(n18772), .ZN(n23843) );
  INV_X1 U17203 ( .A(n18772), .ZN(n23844) );
  INV_X1 U17204 ( .A(n18773), .ZN(n23845) );
  INV_X1 U17205 ( .A(n18773), .ZN(n23846) );
  INV_X1 U17206 ( .A(n18774), .ZN(n23847) );
  INV_X1 U17207 ( .A(n18774), .ZN(n23848) );
  INV_X1 U17208 ( .A(n18775), .ZN(n23849) );
  INV_X1 U17209 ( .A(n18775), .ZN(n23850) );
  INV_X1 U17210 ( .A(n18776), .ZN(n23851) );
  INV_X1 U17211 ( .A(n18776), .ZN(n23852) );
  INV_X1 U17212 ( .A(n18777), .ZN(n23853) );
  INV_X1 U17213 ( .A(n18777), .ZN(n23854) );
  INV_X1 U17214 ( .A(n18778), .ZN(n23855) );
  INV_X1 U17215 ( .A(n18778), .ZN(n23856) );
  INV_X1 U17216 ( .A(n18779), .ZN(n23857) );
  INV_X1 U17217 ( .A(n18779), .ZN(n23858) );
  INV_X1 U17218 ( .A(n18780), .ZN(n23859) );
  INV_X1 U17219 ( .A(n18780), .ZN(n23860) );
  INV_X1 U17220 ( .A(n18781), .ZN(n23861) );
  INV_X1 U17221 ( .A(n18781), .ZN(n23862) );
  INV_X1 U17222 ( .A(n18782), .ZN(n23863) );
  INV_X1 U17223 ( .A(n18782), .ZN(n23864) );
  INV_X1 U17224 ( .A(n18783), .ZN(n23865) );
  INV_X1 U17225 ( .A(n18783), .ZN(n23866) );
  INV_X1 U17226 ( .A(n18784), .ZN(n23867) );
  INV_X1 U17227 ( .A(n18784), .ZN(n23868) );
  INV_X1 U17228 ( .A(n18785), .ZN(n23869) );
  INV_X1 U17229 ( .A(n18785), .ZN(n23870) );
  INV_X1 U17230 ( .A(n18786), .ZN(n23871) );
  INV_X1 U17231 ( .A(n18786), .ZN(n23872) );
  INV_X1 U17232 ( .A(n18787), .ZN(n23873) );
  INV_X1 U17233 ( .A(n18787), .ZN(n23874) );
  INV_X1 U17234 ( .A(n18788), .ZN(n23875) );
  INV_X1 U17235 ( .A(n18788), .ZN(n23876) );
  INV_X1 U17236 ( .A(n18789), .ZN(n23877) );
  INV_X1 U17237 ( .A(n18789), .ZN(n23878) );
  INV_X1 U17238 ( .A(n18790), .ZN(n23879) );
  INV_X1 U17239 ( .A(n18790), .ZN(n23880) );
  INV_X1 U17240 ( .A(n18791), .ZN(n23881) );
  INV_X1 U17241 ( .A(n18791), .ZN(n23882) );
  INV_X1 U17242 ( .A(n18792), .ZN(n23883) );
  INV_X1 U17243 ( .A(n18792), .ZN(n23884) );
  INV_X1 U17244 ( .A(n18793), .ZN(n23885) );
  INV_X1 U17245 ( .A(n18793), .ZN(n23886) );
  INV_X1 U17246 ( .A(n18794), .ZN(n23887) );
  INV_X1 U17247 ( .A(n18794), .ZN(n23888) );
  INV_X1 U17248 ( .A(n18795), .ZN(n23889) );
  INV_X1 U17249 ( .A(n18795), .ZN(n23890) );
  INV_X1 U17250 ( .A(n18796), .ZN(n23891) );
  INV_X1 U17251 ( .A(n18796), .ZN(n23892) );
  INV_X1 U17252 ( .A(n18797), .ZN(n23893) );
  INV_X1 U17253 ( .A(n18797), .ZN(n23894) );
  INV_X1 U17254 ( .A(n18798), .ZN(n23895) );
  INV_X1 U17255 ( .A(n18798), .ZN(n23896) );
  INV_X1 U17256 ( .A(n18799), .ZN(n23897) );
  INV_X1 U17257 ( .A(n18799), .ZN(n23898) );
  INV_X1 U17258 ( .A(n18800), .ZN(n23899) );
  INV_X1 U17259 ( .A(n18800), .ZN(n23900) );
  INV_X1 U17260 ( .A(n18801), .ZN(n23901) );
  INV_X1 U17261 ( .A(n18801), .ZN(n23902) );
  INV_X1 U17262 ( .A(n18802), .ZN(n23903) );
  INV_X1 U17263 ( .A(n18802), .ZN(n23904) );
  INV_X1 U17264 ( .A(n18803), .ZN(n23905) );
  INV_X1 U17265 ( .A(n18803), .ZN(n23906) );
  INV_X1 U17266 ( .A(n18804), .ZN(n23907) );
  INV_X1 U17267 ( .A(n18804), .ZN(n23908) );
  INV_X1 U17268 ( .A(n18805), .ZN(n23909) );
  INV_X1 U17269 ( .A(n18805), .ZN(n23910) );
  INV_X1 U17270 ( .A(n18806), .ZN(n23911) );
  INV_X1 U17271 ( .A(n18806), .ZN(n23912) );
  INV_X1 U17272 ( .A(n18807), .ZN(n23913) );
  INV_X1 U17273 ( .A(n18807), .ZN(n23914) );
  INV_X1 U17274 ( .A(n18808), .ZN(n23915) );
  INV_X1 U17275 ( .A(n18808), .ZN(n23916) );
  INV_X1 U17276 ( .A(n18809), .ZN(n23917) );
  INV_X1 U17277 ( .A(n18809), .ZN(n23918) );
  INV_X1 U17278 ( .A(n18810), .ZN(n23919) );
  INV_X1 U17279 ( .A(n18810), .ZN(n23920) );
  INV_X1 U17280 ( .A(n18811), .ZN(n23921) );
  INV_X1 U17281 ( .A(n18811), .ZN(n23922) );
  INV_X1 U17282 ( .A(n18812), .ZN(n23923) );
  INV_X1 U17283 ( .A(n18812), .ZN(n23924) );
  INV_X1 U17284 ( .A(n18813), .ZN(n23925) );
  INV_X1 U17285 ( .A(n18813), .ZN(n23926) );
  INV_X1 U17286 ( .A(n18814), .ZN(n23927) );
  INV_X1 U17287 ( .A(n18814), .ZN(n23928) );
  INV_X1 U17288 ( .A(n18815), .ZN(n23929) );
  INV_X1 U17289 ( .A(n18815), .ZN(n23930) );
  INV_X1 U17290 ( .A(n18816), .ZN(n23931) );
  INV_X1 U17291 ( .A(n18816), .ZN(n23932) );
  INV_X1 U17292 ( .A(n18817), .ZN(n23933) );
  INV_X1 U17293 ( .A(n18817), .ZN(n23934) );
  INV_X1 U17294 ( .A(n17072), .ZN(n23935) );
  INV_X1 U17295 ( .A(n23935), .ZN(n23936) );
  INV_X1 U17296 ( .A(n23935), .ZN(n23937) );
  INV_X1 U17297 ( .A(r899_B_7_), .ZN(n23938) );
  INV_X1 U17298 ( .A(n17069), .ZN(n23939) );
  INV_X1 U17299 ( .A(n23939), .ZN(n23940) );
  INV_X1 U17300 ( .A(n23939), .ZN(n23941) );
  INV_X1 U17301 ( .A(r899_B_6_), .ZN(n23942) );
  INV_X1 U17302 ( .A(n23942), .ZN(n23943) );
  INV_X1 U17303 ( .A(n23945), .ZN(n23944) );
  INV_X1 U17304 ( .A(n26605), .ZN(n23945) );
  INV_X1 U17305 ( .A(n23945), .ZN(n23946) );
  INV_X1 U17306 ( .A(r899_B_3_), .ZN(n23947) );
  INV_X1 U17307 ( .A(r899_B_3_), .ZN(n23948) );
  INV_X1 U17308 ( .A(n26606), .ZN(n23949) );
  INV_X1 U17309 ( .A(n23949), .ZN(n23950) );
  INV_X1 U17310 ( .A(n26607), .ZN(n23951) );
  INV_X1 U17311 ( .A(n23951), .ZN(n23952) );
  INV_X1 U17312 ( .A(n23951), .ZN(n23953) );
  INV_X1 U17313 ( .A(n26611), .ZN(n23954) );
  INV_X1 U17314 ( .A(n23954), .ZN(n23955) );
  INV_X1 U17315 ( .A(n23954), .ZN(n23956) );
  INV_X1 U17316 ( .A(n26612), .ZN(n23957) );
  INV_X1 U17317 ( .A(n23957), .ZN(n23958) );
  INV_X1 U17318 ( .A(n23957), .ZN(n23959) );
  INV_X1 U17319 ( .A(n26962), .ZN(n23960) );
  INV_X1 U17320 ( .A(n18820), .ZN(n23961) );
  INV_X1 U17321 ( .A(n18820), .ZN(n23962) );
  INV_X1 U17322 ( .A(n18821), .ZN(n23963) );
  INV_X1 U17323 ( .A(n18821), .ZN(n23964) );
  INV_X1 U17324 ( .A(n18822), .ZN(n23965) );
  INV_X1 U17325 ( .A(n18822), .ZN(n23966) );
  CLKBUF_X1 U17326 ( .A(n23968), .Z(n23967) );
  CLKBUF_X1 U17327 ( .A(n21063), .Z(n23968) );
  INV_X1 U17328 ( .A(n26621), .ZN(n23969) );
  INV_X1 U17329 ( .A(n23969), .ZN(n23970) );
  INV_X1 U17330 ( .A(n23969), .ZN(n23971) );
  INV_X1 U17331 ( .A(n19273), .ZN(n23972) );
  INV_X1 U17332 ( .A(n23972), .ZN(n23973) );
  INV_X1 U17333 ( .A(n23972), .ZN(n23974) );
  CLKBUF_X1 U17334 ( .A(n23976), .Z(n23975) );
  CLKBUF_X1 U17335 ( .A(n21001), .Z(n23976) );
  INV_X1 U17336 ( .A(n26623), .ZN(n23977) );
  INV_X1 U17337 ( .A(n23977), .ZN(n23978) );
  INV_X1 U17338 ( .A(n23977), .ZN(n23979) );
  INV_X1 U17339 ( .A(n19274), .ZN(n23980) );
  INV_X1 U17340 ( .A(n23980), .ZN(n23981) );
  INV_X1 U17341 ( .A(n23980), .ZN(n23982) );
  CLKBUF_X1 U17342 ( .A(n23984), .Z(n23983) );
  CLKBUF_X1 U17343 ( .A(n22686), .Z(n23984) );
  INV_X1 U17344 ( .A(n26629), .ZN(n23985) );
  INV_X1 U17345 ( .A(n23985), .ZN(n23986) );
  INV_X1 U17346 ( .A(n23985), .ZN(n23987) );
  INV_X1 U17347 ( .A(n23984), .ZN(n23988) );
  INV_X1 U17348 ( .A(n23988), .ZN(n23989) );
  INV_X1 U17349 ( .A(n23988), .ZN(n23990) );
  CLKBUF_X1 U17350 ( .A(n23992), .Z(n23991) );
  CLKBUF_X1 U17351 ( .A(n21066), .Z(n23992) );
  INV_X1 U17352 ( .A(n26631), .ZN(n23993) );
  INV_X1 U17353 ( .A(n23993), .ZN(n23994) );
  INV_X1 U17354 ( .A(n23993), .ZN(n23995) );
  INV_X1 U17355 ( .A(n23992), .ZN(n23996) );
  INV_X1 U17356 ( .A(n23996), .ZN(n23997) );
  INV_X1 U17357 ( .A(n23996), .ZN(n23998) );
  CLKBUF_X1 U17358 ( .A(n24000), .Z(n23999) );
  CLKBUF_X1 U17359 ( .A(n21004), .Z(n24000) );
  INV_X1 U17360 ( .A(n26633), .ZN(n24001) );
  INV_X1 U17361 ( .A(n24001), .ZN(n24002) );
  INV_X1 U17362 ( .A(n24001), .ZN(n24003) );
  INV_X1 U17363 ( .A(n24000), .ZN(n24004) );
  INV_X1 U17364 ( .A(n24004), .ZN(n24005) );
  INV_X1 U17365 ( .A(n24004), .ZN(n24006) );
  CLKBUF_X1 U17366 ( .A(n24008), .Z(n24007) );
  CLKBUF_X1 U17367 ( .A(n21059), .Z(n24008) );
  INV_X1 U17368 ( .A(n26635), .ZN(n24009) );
  INV_X1 U17369 ( .A(n24009), .ZN(n24010) );
  INV_X1 U17370 ( .A(n24009), .ZN(n24011) );
  INV_X1 U17371 ( .A(n24008), .ZN(n24012) );
  INV_X1 U17372 ( .A(n24012), .ZN(n24013) );
  INV_X1 U17373 ( .A(n24012), .ZN(n24014) );
  CLKBUF_X1 U17374 ( .A(r899_B_9_), .Z(n24015) );
  CLKBUF_X1 U17375 ( .A(n24017), .Z(n24016) );
  CLKBUF_X1 U17376 ( .A(n45500), .Z(n24017) );
  NOR2_X1 U17377 ( .A1(n24220), .A2(n4567), .ZN(n45500) );
  INV_X1 U17378 ( .A(n19279), .ZN(n24018) );
  INV_X1 U17379 ( .A(n24018), .ZN(n24019) );
  INV_X1 U17380 ( .A(n24018), .ZN(n24020) );
  INV_X1 U17381 ( .A(n24017), .ZN(n24021) );
  INV_X1 U17382 ( .A(n24021), .ZN(n24022) );
  INV_X1 U17383 ( .A(n24021), .ZN(n24023) );
  CLKBUF_X1 U17384 ( .A(n24025), .Z(n24024) );
  CLKBUF_X1 U17385 ( .A(n3079), .Z(n24025) );
  NOR2_X1 U17386 ( .A1(n25291), .A2(n3099), .ZN(n3079) );
  INV_X1 U17387 ( .A(n19280), .ZN(n24026) );
  INV_X1 U17388 ( .A(n24026), .ZN(n24027) );
  INV_X1 U17389 ( .A(n24026), .ZN(n24028) );
  INV_X1 U17390 ( .A(n24025), .ZN(n24029) );
  INV_X1 U17391 ( .A(n24029), .ZN(n24030) );
  INV_X1 U17392 ( .A(n24029), .ZN(n24031) );
  CLKBUF_X1 U17393 ( .A(n24033), .Z(n24032) );
  CLKBUF_X1 U17394 ( .A(n3078), .Z(n24033) );
  INV_X1 U17395 ( .A(n19281), .ZN(n24034) );
  INV_X1 U17396 ( .A(n24034), .ZN(n24035) );
  INV_X1 U17397 ( .A(n24034), .ZN(n24036) );
  INV_X1 U17398 ( .A(n24033), .ZN(n24037) );
  INV_X1 U17399 ( .A(n24037), .ZN(n24038) );
  INV_X1 U17400 ( .A(n24037), .ZN(n24039) );
  CLKBUF_X1 U17401 ( .A(n24041), .Z(n24040) );
  CLKBUF_X1 U17402 ( .A(n45490), .Z(n24041) );
  INV_X1 U17403 ( .A(n19282), .ZN(n24042) );
  INV_X1 U17404 ( .A(n24042), .ZN(n24043) );
  INV_X1 U17405 ( .A(n24042), .ZN(n24044) );
  INV_X1 U17406 ( .A(n24041), .ZN(n24045) );
  INV_X1 U17407 ( .A(n24045), .ZN(n24046) );
  INV_X1 U17408 ( .A(n24045), .ZN(n24047) );
  CLKBUF_X1 U17409 ( .A(n24049), .Z(n24048) );
  CLKBUF_X1 U17410 ( .A(n47060), .Z(n24049) );
  INV_X1 U17411 ( .A(n24049), .ZN(n24050) );
  INV_X1 U17412 ( .A(n24050), .ZN(n24051) );
  INV_X1 U17413 ( .A(n24050), .ZN(n24052) );
  INV_X1 U17414 ( .A(n19283), .ZN(n24053) );
  INV_X1 U17415 ( .A(n24053), .ZN(n24054) );
  INV_X1 U17416 ( .A(n24053), .ZN(n24055) );
  CLKBUF_X1 U17417 ( .A(n24057), .Z(n24056) );
  CLKBUF_X1 U17418 ( .A(n20922), .Z(n24057) );
  INV_X1 U17419 ( .A(n22717), .ZN(n24058) );
  INV_X1 U17420 ( .A(n24058), .ZN(n24059) );
  INV_X1 U17421 ( .A(n24058), .ZN(n24060) );
  CLKBUF_X1 U17422 ( .A(n24062), .Z(n24061) );
  CLKBUF_X1 U17423 ( .A(n21407), .Z(n24062) );
  INV_X1 U17424 ( .A(n22720), .ZN(n24063) );
  INV_X1 U17425 ( .A(n24063), .ZN(n24064) );
  INV_X1 U17426 ( .A(n24063), .ZN(n24065) );
  CLKBUF_X1 U17427 ( .A(n24067), .Z(n24066) );
  CLKBUF_X1 U17428 ( .A(n20927), .Z(n24067) );
  INV_X1 U17429 ( .A(n22723), .ZN(n24068) );
  INV_X1 U17430 ( .A(n24068), .ZN(n24069) );
  INV_X1 U17431 ( .A(n24068), .ZN(n24070) );
  CLKBUF_X1 U17432 ( .A(n22725), .Z(n24071) );
  INV_X1 U17433 ( .A(n24071), .ZN(n24072) );
  INV_X1 U17434 ( .A(n24072), .ZN(n24073) );
  INV_X1 U17435 ( .A(n24072), .ZN(n24074) );
  CLKBUF_X1 U17436 ( .A(n24076), .Z(n24075) );
  CLKBUF_X1 U17437 ( .A(n21413), .Z(n24076) );
  INV_X1 U17438 ( .A(n22730), .ZN(n24077) );
  INV_X1 U17439 ( .A(n24077), .ZN(n24078) );
  INV_X1 U17440 ( .A(n24077), .ZN(n24079) );
  INV_X1 U17441 ( .A(n18824), .ZN(n24080) );
  INV_X1 U17442 ( .A(n18824), .ZN(n24081) );
  INV_X1 U17443 ( .A(n18825), .ZN(n24082) );
  INV_X1 U17444 ( .A(n18825), .ZN(n24083) );
  INV_X1 U17445 ( .A(n18826), .ZN(n24084) );
  INV_X1 U17446 ( .A(n18826), .ZN(n24085) );
  INV_X1 U17447 ( .A(n18827), .ZN(n24086) );
  INV_X1 U17448 ( .A(n18827), .ZN(n24087) );
  CLKBUF_X1 U17449 ( .A(n4818), .Z(n24088) );
  INV_X1 U17450 ( .A(n24088), .ZN(n24089) );
  INV_X1 U17451 ( .A(n24089), .ZN(n24090) );
  INV_X1 U17452 ( .A(n24089), .ZN(n24091) );
  CLKBUF_X1 U17453 ( .A(n4819), .Z(n24092) );
  INV_X1 U17454 ( .A(n24092), .ZN(n24093) );
  INV_X1 U17455 ( .A(n24093), .ZN(n24094) );
  INV_X1 U17456 ( .A(n24093), .ZN(n24095) );
  CLKBUF_X1 U17457 ( .A(n47050), .Z(n24096) );
  INV_X1 U17458 ( .A(n24096), .ZN(n24097) );
  INV_X1 U17459 ( .A(n24097), .ZN(n24098) );
  INV_X1 U17460 ( .A(n24097), .ZN(n24099) );
  CLKBUF_X1 U17461 ( .A(n24101), .Z(n24100) );
  CLKBUF_X1 U17462 ( .A(n27796), .Z(n24101) );
  CLKBUF_X1 U17463 ( .A(n24103), .Z(n24102) );
  CLKBUF_X1 U17464 ( .A(n27804), .Z(n24103) );
  INV_X1 U17465 ( .A(n26583), .ZN(n24104) );
  INV_X1 U17466 ( .A(n24104), .ZN(n24105) );
  INV_X1 U17467 ( .A(n24104), .ZN(n24106) );
  INV_X1 U17468 ( .A(n18828), .ZN(n24107) );
  INV_X1 U17469 ( .A(n18828), .ZN(n24108) );
  INV_X1 U17470 ( .A(n18829), .ZN(n24109) );
  INV_X1 U17471 ( .A(n18829), .ZN(n24110) );
  INV_X1 U17472 ( .A(n18830), .ZN(n24111) );
  INV_X1 U17473 ( .A(n18830), .ZN(n24112) );
  INV_X1 U17474 ( .A(n18831), .ZN(n24113) );
  INV_X1 U17475 ( .A(n18831), .ZN(n24114) );
  INV_X1 U17476 ( .A(n18832), .ZN(n24115) );
  INV_X1 U17477 ( .A(n18832), .ZN(n24116) );
  INV_X1 U17478 ( .A(n18833), .ZN(n24117) );
  INV_X1 U17479 ( .A(n18833), .ZN(n24118) );
  INV_X1 U17480 ( .A(n18834), .ZN(n24119) );
  INV_X1 U17481 ( .A(n18834), .ZN(n24120) );
  INV_X1 U17482 ( .A(n18835), .ZN(n24121) );
  INV_X1 U17483 ( .A(n18835), .ZN(n24122) );
  INV_X1 U17484 ( .A(n18836), .ZN(n24123) );
  INV_X1 U17485 ( .A(n18836), .ZN(n24124) );
  INV_X1 U17486 ( .A(n18837), .ZN(n24125) );
  INV_X1 U17487 ( .A(n18837), .ZN(n24126) );
  INV_X1 U17488 ( .A(n18838), .ZN(n24127) );
  INV_X1 U17489 ( .A(n18838), .ZN(n24128) );
  INV_X1 U17490 ( .A(n18839), .ZN(n24129) );
  INV_X1 U17491 ( .A(n18839), .ZN(n24130) );
  INV_X1 U17492 ( .A(n18840), .ZN(n24131) );
  INV_X1 U17493 ( .A(n18840), .ZN(n24132) );
  INV_X1 U17494 ( .A(n18841), .ZN(n24133) );
  INV_X1 U17495 ( .A(n18841), .ZN(n24134) );
  INV_X1 U17496 ( .A(n18842), .ZN(n24135) );
  INV_X1 U17497 ( .A(n18842), .ZN(n24136) );
  INV_X1 U17498 ( .A(n18843), .ZN(n24137) );
  INV_X1 U17499 ( .A(n18843), .ZN(n24138) );
  INV_X1 U17500 ( .A(n18844), .ZN(n24139) );
  INV_X1 U17501 ( .A(n18844), .ZN(n24140) );
  CLKBUF_X1 U17502 ( .A(n51360), .Z(n24141) );
  INV_X1 U17503 ( .A(n18845), .ZN(n24142) );
  INV_X1 U17504 ( .A(n18845), .ZN(n24143) );
  INV_X1 U17505 ( .A(n18846), .ZN(n24144) );
  INV_X1 U17506 ( .A(n18846), .ZN(n24145) );
  INV_X1 U17507 ( .A(n18847), .ZN(n24146) );
  INV_X1 U17508 ( .A(n18847), .ZN(n24147) );
  INV_X1 U17509 ( .A(n18848), .ZN(n24148) );
  INV_X1 U17510 ( .A(n18848), .ZN(n24149) );
  CLKBUF_X1 U17511 ( .A(n27789), .Z(n24150) );
  INV_X1 U17512 ( .A(n24150), .ZN(n24151) );
  INV_X1 U17513 ( .A(n24151), .ZN(n24152) );
  INV_X1 U17514 ( .A(n24151), .ZN(n24153) );
  INV_X1 U17515 ( .A(n19298), .ZN(n24154) );
  INV_X1 U17516 ( .A(n24154), .ZN(n24155) );
  INV_X1 U17517 ( .A(n24154), .ZN(n24156) );
  CLKBUF_X1 U17518 ( .A(n27726), .Z(n24157) );
  INV_X1 U17519 ( .A(n19299), .ZN(n24158) );
  INV_X1 U17520 ( .A(n24158), .ZN(n24159) );
  INV_X1 U17521 ( .A(n24158), .ZN(n24160) );
  CLKBUF_X1 U17522 ( .A(n4714), .Z(n24161) );
  INV_X1 U17523 ( .A(n26710), .ZN(n24162) );
  INV_X1 U17524 ( .A(n24162), .ZN(n24163) );
  INV_X1 U17525 ( .A(n24162), .ZN(n24164) );
  CLKBUF_X1 U17526 ( .A(n4713), .Z(n24165) );
  INV_X1 U17527 ( .A(n26714), .ZN(n24166) );
  INV_X1 U17528 ( .A(n24166), .ZN(n24167) );
  INV_X1 U17529 ( .A(n24166), .ZN(n24168) );
  INV_X1 U17530 ( .A(n18849), .ZN(n24169) );
  INV_X1 U17531 ( .A(n18849), .ZN(n24170) );
  INV_X1 U17532 ( .A(n54230), .ZN(n24171) );
  INV_X1 U17533 ( .A(n24171), .ZN(n24172) );
  INV_X1 U17534 ( .A(n24171), .ZN(n24173) );
  INV_X1 U17535 ( .A(n27797), .ZN(n24174) );
  INV_X1 U17536 ( .A(n27797), .ZN(n24175) );
  INV_X1 U17537 ( .A(n26719), .ZN(n24176) );
  INV_X1 U17538 ( .A(n24176), .ZN(n24177) );
  INV_X1 U17539 ( .A(n24176), .ZN(n24178) );
  INV_X1 U17540 ( .A(n18850), .ZN(n24179) );
  INV_X1 U17541 ( .A(n18850), .ZN(n24180) );
  INV_X1 U17542 ( .A(n26722), .ZN(n24181) );
  INV_X1 U17543 ( .A(n24181), .ZN(n24182) );
  INV_X1 U17544 ( .A(n24181), .ZN(n24183) );
  INV_X1 U17545 ( .A(n18851), .ZN(n24184) );
  INV_X1 U17546 ( .A(n18851), .ZN(n24185) );
  INV_X1 U17547 ( .A(n26727), .ZN(n24186) );
  INV_X1 U17548 ( .A(n24186), .ZN(n24187) );
  INV_X1 U17549 ( .A(n24186), .ZN(n24188) );
  INV_X1 U17550 ( .A(n26728), .ZN(n24189) );
  INV_X1 U17551 ( .A(n24189), .ZN(n24190) );
  INV_X1 U17552 ( .A(n24189), .ZN(n24191) );
  INV_X1 U17553 ( .A(n18854), .ZN(n24192) );
  INV_X1 U17554 ( .A(n18854), .ZN(n24193) );
  INV_X1 U17555 ( .A(n26730), .ZN(n24194) );
  INV_X1 U17556 ( .A(n24194), .ZN(n24195) );
  INV_X1 U17557 ( .A(n24194), .ZN(n24196) );
  INV_X1 U17558 ( .A(n26731), .ZN(n24197) );
  INV_X1 U17559 ( .A(n24197), .ZN(n24198) );
  INV_X1 U17560 ( .A(n24197), .ZN(n24199) );
  INV_X1 U17561 ( .A(n3236), .ZN(n24200) );
  INV_X1 U17562 ( .A(n24200), .ZN(n24201) );
  INV_X1 U17563 ( .A(n24200), .ZN(n24202) );
  INV_X1 U17564 ( .A(n26733), .ZN(n24203) );
  INV_X1 U17565 ( .A(n24203), .ZN(n24204) );
  INV_X1 U17566 ( .A(n24203), .ZN(n24205) );
  INV_X1 U17567 ( .A(n3443), .ZN(n24206) );
  INV_X1 U17568 ( .A(n24206), .ZN(n24207) );
  INV_X1 U17569 ( .A(n24206), .ZN(n24208) );
  INV_X1 U17570 ( .A(n267401), .ZN(n24209) );
  INV_X1 U17571 ( .A(n24209), .ZN(n24210) );
  INV_X1 U17572 ( .A(n24209), .ZN(n24211) );
  INV_X1 U17573 ( .A(n18855), .ZN(n24212) );
  INV_X1 U17574 ( .A(n18855), .ZN(n24213) );
  INV_X1 U17575 ( .A(n18856), .ZN(n24214) );
  INV_X1 U17576 ( .A(n18856), .ZN(n24215) );
  INV_X1 U17577 ( .A(n18857), .ZN(n24216) );
  INV_X1 U17578 ( .A(n18857), .ZN(n24217) );
  INV_X1 U17579 ( .A(n18858), .ZN(n24218) );
  INV_X1 U17580 ( .A(n18858), .ZN(n24219) );
  INV_X1 U17581 ( .A(n18859), .ZN(n24220) );
  INV_X1 U17582 ( .A(n18859), .ZN(n24221) );
  CLKBUF_X1 U17583 ( .A(n27802), .Z(n24222) );
  INV_X1 U17584 ( .A(n21326), .ZN(n27802) );
  INV_X1 U17585 ( .A(n26748), .ZN(n24223) );
  INV_X1 U17586 ( .A(n24223), .ZN(n24224) );
  INV_X1 U17587 ( .A(n24223), .ZN(n24225) );
  CLKBUF_X1 U17588 ( .A(n27798), .Z(n24226) );
  INV_X1 U17589 ( .A(n21337), .ZN(n27798) );
  INV_X1 U17590 ( .A(n26751), .ZN(n24227) );
  INV_X1 U17591 ( .A(n24227), .ZN(n24228) );
  INV_X1 U17592 ( .A(n24227), .ZN(n24229) );
  INV_X1 U17593 ( .A(n22832), .ZN(n24230) );
  INV_X1 U17594 ( .A(n24230), .ZN(n24231) );
  INV_X1 U17595 ( .A(n24230), .ZN(n24232) );
  INV_X1 U17596 ( .A(n22840), .ZN(n24233) );
  INV_X1 U17597 ( .A(n24233), .ZN(n24234) );
  INV_X1 U17598 ( .A(n24233), .ZN(n24235) );
  INV_X1 U17599 ( .A(n22842), .ZN(n24236) );
  INV_X1 U17600 ( .A(n24236), .ZN(n24237) );
  INV_X1 U17601 ( .A(n24236), .ZN(n24238) );
  INV_X1 U17602 ( .A(n22844), .ZN(n24239) );
  INV_X1 U17603 ( .A(n24239), .ZN(n24240) );
  INV_X1 U17604 ( .A(n24239), .ZN(n24241) );
  INV_X1 U17605 ( .A(n22849), .ZN(n24242) );
  INV_X1 U17606 ( .A(n24242), .ZN(n24243) );
  INV_X1 U17607 ( .A(n24242), .ZN(n24244) );
  INV_X1 U17608 ( .A(n22851), .ZN(n24245) );
  INV_X1 U17609 ( .A(n24245), .ZN(n24246) );
  INV_X1 U17610 ( .A(n24245), .ZN(n24247) );
  INV_X1 U17611 ( .A(n22856), .ZN(n24248) );
  INV_X1 U17612 ( .A(n24248), .ZN(n24249) );
  INV_X1 U17613 ( .A(n24248), .ZN(n24250) );
  INV_X1 U17614 ( .A(n22861), .ZN(n24251) );
  INV_X1 U17615 ( .A(n24251), .ZN(n24252) );
  INV_X1 U17616 ( .A(n24251), .ZN(n24253) );
  INV_X1 U17617 ( .A(n22866), .ZN(n24254) );
  INV_X1 U17618 ( .A(n24254), .ZN(n24255) );
  INV_X1 U17619 ( .A(n24254), .ZN(n24256) );
  INV_X1 U17620 ( .A(n26779), .ZN(n24257) );
  INV_X1 U17621 ( .A(n24257), .ZN(n24258) );
  INV_X1 U17622 ( .A(n24257), .ZN(n24259) );
  INV_X1 U17623 ( .A(n22871), .ZN(n24260) );
  INV_X1 U17624 ( .A(n24260), .ZN(n24261) );
  INV_X1 U17625 ( .A(n24260), .ZN(n24262) );
  INV_X1 U17626 ( .A(n22872), .ZN(n24263) );
  INV_X1 U17627 ( .A(n24263), .ZN(n24264) );
  INV_X1 U17628 ( .A(n24263), .ZN(n24265) );
  INV_X1 U17629 ( .A(n20505), .ZN(n24266) );
  INV_X1 U17630 ( .A(n24266), .ZN(n24267) );
  INV_X1 U17631 ( .A(n24266), .ZN(n24268) );
  INV_X1 U17632 ( .A(n26784), .ZN(n24269) );
  INV_X1 U17633 ( .A(n24269), .ZN(n24270) );
  INV_X1 U17634 ( .A(n24269), .ZN(n24271) );
  INV_X1 U17635 ( .A(n19265), .ZN(n24272) );
  INV_X1 U17636 ( .A(n24272), .ZN(n24273) );
  INV_X1 U17637 ( .A(n24272), .ZN(n24274) );
  INV_X1 U17638 ( .A(n26788), .ZN(n24275) );
  INV_X1 U17639 ( .A(n24275), .ZN(n24276) );
  INV_X1 U17640 ( .A(n24275), .ZN(n24277) );
  INV_X1 U17641 ( .A(n267901), .ZN(n24278) );
  INV_X1 U17642 ( .A(n24278), .ZN(n24279) );
  INV_X1 U17643 ( .A(n24278), .ZN(n24280) );
  INV_X1 U17644 ( .A(n26791), .ZN(n24281) );
  INV_X1 U17645 ( .A(n24281), .ZN(n24282) );
  INV_X1 U17646 ( .A(n24281), .ZN(n24283) );
  INV_X1 U17647 ( .A(n19264), .ZN(n24284) );
  INV_X1 U17648 ( .A(n24284), .ZN(n24285) );
  INV_X1 U17649 ( .A(n24284), .ZN(n24286) );
  INV_X1 U17650 ( .A(n26795), .ZN(n24287) );
  INV_X1 U17651 ( .A(n24287), .ZN(n24288) );
  INV_X1 U17652 ( .A(n24287), .ZN(n24289) );
  INV_X1 U17653 ( .A(n26798), .ZN(n24290) );
  INV_X1 U17654 ( .A(n24290), .ZN(n24291) );
  INV_X1 U17655 ( .A(n24290), .ZN(n24292) );
  INV_X1 U17656 ( .A(n27259), .ZN(n24293) );
  INV_X1 U17657 ( .A(n24293), .ZN(n24294) );
  INV_X1 U17658 ( .A(n24293), .ZN(n24295) );
  INV_X1 U17659 ( .A(n268001), .ZN(n24296) );
  INV_X1 U17660 ( .A(n24296), .ZN(n24297) );
  INV_X1 U17661 ( .A(n24296), .ZN(n24298) );
  INV_X1 U17662 ( .A(n26801), .ZN(n24299) );
  INV_X1 U17663 ( .A(n24299), .ZN(n24300) );
  INV_X1 U17664 ( .A(n24299), .ZN(n24301) );
  INV_X1 U17665 ( .A(n26804), .ZN(n24302) );
  INV_X1 U17666 ( .A(n24302), .ZN(n24303) );
  INV_X1 U17667 ( .A(n24302), .ZN(n24304) );
  INV_X1 U17668 ( .A(n27171), .ZN(n24305) );
  INV_X1 U17669 ( .A(n24305), .ZN(n24306) );
  INV_X1 U17670 ( .A(n24305), .ZN(n24307) );
  INV_X1 U17671 ( .A(n26807), .ZN(n24308) );
  INV_X1 U17672 ( .A(n24308), .ZN(n24309) );
  INV_X1 U17673 ( .A(n24308), .ZN(n24310) );
  INV_X1 U17674 ( .A(n26808), .ZN(n24311) );
  INV_X1 U17675 ( .A(n24311), .ZN(n24312) );
  INV_X1 U17676 ( .A(n24311), .ZN(n24313) );
  INV_X1 U17677 ( .A(n18921), .ZN(n24314) );
  INV_X1 U17678 ( .A(n24314), .ZN(n24315) );
  INV_X1 U17679 ( .A(n24314), .ZN(n24316) );
  INV_X1 U17680 ( .A(n18920), .ZN(n24317) );
  INV_X1 U17681 ( .A(n24317), .ZN(n24318) );
  INV_X1 U17682 ( .A(n24317), .ZN(n24319) );
  INV_X1 U17683 ( .A(n18921), .ZN(n24320) );
  INV_X1 U17684 ( .A(n24320), .ZN(n24321) );
  INV_X1 U17685 ( .A(n24320), .ZN(n24322) );
  INV_X1 U17686 ( .A(n18920), .ZN(n24323) );
  INV_X1 U17687 ( .A(n24323), .ZN(n24324) );
  INV_X1 U17688 ( .A(n24323), .ZN(n24325) );
  INV_X1 U17689 ( .A(n18919), .ZN(n24326) );
  INV_X1 U17690 ( .A(n24326), .ZN(n24327) );
  INV_X1 U17691 ( .A(n24326), .ZN(n24328) );
  INV_X1 U17692 ( .A(n18918), .ZN(n24329) );
  INV_X1 U17693 ( .A(n24329), .ZN(n24330) );
  INV_X1 U17694 ( .A(n24329), .ZN(n24331) );
  INV_X1 U17695 ( .A(n18919), .ZN(n24332) );
  INV_X1 U17696 ( .A(n24332), .ZN(n24333) );
  INV_X1 U17697 ( .A(n24332), .ZN(n24334) );
  INV_X1 U17698 ( .A(n18918), .ZN(n24335) );
  INV_X1 U17699 ( .A(n24335), .ZN(n24336) );
  INV_X1 U17700 ( .A(n24335), .ZN(n24337) );
  INV_X1 U17701 ( .A(n26842), .ZN(n24338) );
  INV_X1 U17702 ( .A(n24338), .ZN(n24339) );
  INV_X1 U17703 ( .A(n24338), .ZN(n24340) );
  INV_X1 U17704 ( .A(n19261), .ZN(n24341) );
  INV_X1 U17705 ( .A(n24341), .ZN(n24342) );
  INV_X1 U17706 ( .A(n24341), .ZN(n24343) );
  INV_X1 U17707 ( .A(n26846), .ZN(n24344) );
  INV_X1 U17708 ( .A(n24344), .ZN(n24345) );
  INV_X1 U17709 ( .A(n24344), .ZN(n24346) );
  INV_X1 U17710 ( .A(n19260), .ZN(n24347) );
  INV_X1 U17711 ( .A(n24347), .ZN(n24348) );
  INV_X1 U17712 ( .A(n24347), .ZN(n24349) );
  INV_X1 U17713 ( .A(n26849), .ZN(n24350) );
  INV_X1 U17714 ( .A(n24350), .ZN(n24351) );
  INV_X1 U17715 ( .A(n24350), .ZN(n24352) );
  INV_X1 U17716 ( .A(n19259), .ZN(n24353) );
  INV_X1 U17717 ( .A(n24353), .ZN(n24354) );
  INV_X1 U17718 ( .A(n24353), .ZN(n24355) );
  INV_X1 U17719 ( .A(n19258), .ZN(n24356) );
  INV_X1 U17720 ( .A(n24356), .ZN(n24357) );
  INV_X1 U17721 ( .A(n24356), .ZN(n24358) );
  INV_X1 U17722 ( .A(n26853), .ZN(n24359) );
  INV_X1 U17723 ( .A(n24359), .ZN(n24360) );
  INV_X1 U17724 ( .A(n24359), .ZN(n24361) );
  INV_X1 U17725 ( .A(n18860), .ZN(n24362) );
  INV_X1 U17726 ( .A(n18860), .ZN(n24363) );
  INV_X1 U17727 ( .A(n18861), .ZN(n24364) );
  INV_X1 U17728 ( .A(n24364), .ZN(n24365) );
  INV_X1 U17729 ( .A(n24364), .ZN(n24366) );
  INV_X1 U17730 ( .A(n26855), .ZN(n24367) );
  INV_X1 U17731 ( .A(n24367), .ZN(n24368) );
  INV_X1 U17732 ( .A(n24367), .ZN(n24369) );
  INV_X1 U17733 ( .A(n27116), .ZN(n24370) );
  INV_X1 U17734 ( .A(n27116), .ZN(n24371) );
  INV_X1 U17735 ( .A(n27115), .ZN(n24372) );
  INV_X1 U17736 ( .A(n27115), .ZN(n24373) );
  INV_X1 U17737 ( .A(n26866), .ZN(n24374) );
  INV_X1 U17738 ( .A(n24374), .ZN(n24375) );
  INV_X1 U17739 ( .A(n27114), .ZN(n24376) );
  INV_X1 U17740 ( .A(n18862), .ZN(n24377) );
  INV_X1 U17741 ( .A(n18864), .ZN(n24378) );
  INV_X1 U17742 ( .A(n18864), .ZN(n24379) );
  INV_X1 U17743 ( .A(n18865), .ZN(n24380) );
  INV_X1 U17744 ( .A(n18865), .ZN(n24381) );
  INV_X1 U17745 ( .A(n18866), .ZN(n24382) );
  INV_X1 U17746 ( .A(n18866), .ZN(n24383) );
  INV_X1 U17747 ( .A(n18867), .ZN(n24384) );
  INV_X1 U17748 ( .A(n18867), .ZN(n24385) );
  INV_X1 U17749 ( .A(n27120), .ZN(n24386) );
  INV_X1 U17750 ( .A(n27120), .ZN(n24387) );
  INV_X1 U17751 ( .A(n27119), .ZN(n24388) );
  INV_X1 U17752 ( .A(n27119), .ZN(n24389) );
  INV_X1 U17753 ( .A(n27118), .ZN(n24390) );
  INV_X1 U17754 ( .A(n27118), .ZN(n24391) );
  INV_X1 U17755 ( .A(n27117), .ZN(n24392) );
  INV_X1 U17756 ( .A(n27117), .ZN(n24393) );
  INV_X1 U17757 ( .A(n26902), .ZN(n24394) );
  INV_X1 U17758 ( .A(n24394), .ZN(n24395) );
  INV_X1 U17759 ( .A(n24394), .ZN(n24396) );
  INV_X1 U17760 ( .A(n18868), .ZN(n24397) );
  INV_X1 U17761 ( .A(n18868), .ZN(n24398) );
  INV_X1 U17762 ( .A(n18869), .ZN(n24399) );
  INV_X1 U17763 ( .A(n18869), .ZN(n24400) );
  INV_X1 U17764 ( .A(n18870), .ZN(n24401) );
  INV_X1 U17765 ( .A(n18870), .ZN(n24402) );
  INV_X1 U17766 ( .A(n18871), .ZN(n24403) );
  INV_X1 U17767 ( .A(n18871), .ZN(n24404) );
  INV_X1 U17768 ( .A(n18872), .ZN(n24405) );
  INV_X1 U17769 ( .A(n18872), .ZN(n24406) );
  INV_X1 U17770 ( .A(n18873), .ZN(n24407) );
  INV_X1 U17771 ( .A(n18873), .ZN(n24408) );
  INV_X1 U17772 ( .A(n18874), .ZN(n24409) );
  INV_X1 U17773 ( .A(n18874), .ZN(n24410) );
  INV_X1 U17774 ( .A(n18875), .ZN(n24411) );
  INV_X1 U17775 ( .A(n18875), .ZN(n24412) );
  INV_X1 U17776 ( .A(n18876), .ZN(n24413) );
  INV_X1 U17777 ( .A(n18876), .ZN(n24414) );
  INV_X1 U17778 ( .A(n18877), .ZN(n24415) );
  INV_X1 U17779 ( .A(n18877), .ZN(n24416) );
  CLKBUF_X1 U17780 ( .A(n26923), .Z(n24417) );
  INV_X1 U17781 ( .A(n18878), .ZN(n24418) );
  INV_X1 U17782 ( .A(n18878), .ZN(n24419) );
  INV_X1 U17783 ( .A(n26925), .ZN(n24420) );
  INV_X1 U17784 ( .A(n24420), .ZN(n24421) );
  INV_X1 U17785 ( .A(n24420), .ZN(n24422) );
  INV_X1 U17786 ( .A(n19272), .ZN(n24423) );
  INV_X1 U17787 ( .A(n24423), .ZN(n24424) );
  INV_X1 U17788 ( .A(n24423), .ZN(n24425) );
  INV_X1 U17789 ( .A(n18879), .ZN(n24426) );
  INV_X1 U17790 ( .A(n18879), .ZN(n24427) );
  INV_X1 U17791 ( .A(n27110), .ZN(n24428) );
  INV_X1 U17792 ( .A(n27110), .ZN(n24429) );
  INV_X1 U17793 ( .A(n18880), .ZN(n24430) );
  INV_X1 U17794 ( .A(n18880), .ZN(n24431) );
  INV_X1 U17795 ( .A(n26948), .ZN(n24432) );
  INV_X1 U17796 ( .A(n24432), .ZN(n24433) );
  INV_X1 U17797 ( .A(n24432), .ZN(n24434) );
  INV_X1 U17798 ( .A(n18881), .ZN(n24435) );
  INV_X1 U17799 ( .A(n18881), .ZN(n24436) );
  INV_X1 U17800 ( .A(n26965), .ZN(n24437) );
  INV_X1 U17801 ( .A(n26965), .ZN(n24438) );
  INV_X1 U17802 ( .A(n18882), .ZN(n24439) );
  INV_X1 U17803 ( .A(n18882), .ZN(n24440) );
  INV_X1 U17804 ( .A(n18883), .ZN(n24441) );
  INV_X1 U17805 ( .A(n18883), .ZN(n24442) );
  INV_X1 U17806 ( .A(n18945), .ZN(n24443) );
  INV_X1 U17807 ( .A(n24443), .ZN(n24444) );
  INV_X1 U17808 ( .A(n24443), .ZN(n24445) );
  INV_X1 U17809 ( .A(n18945), .ZN(n24446) );
  INV_X1 U17810 ( .A(n24446), .ZN(n24447) );
  INV_X1 U17811 ( .A(n24446), .ZN(n24448) );
  INV_X1 U17812 ( .A(n18884), .ZN(n24449) );
  INV_X1 U17813 ( .A(n18884), .ZN(n24450) );
  INV_X1 U17814 ( .A(n18885), .ZN(n24451) );
  INV_X1 U17815 ( .A(n18885), .ZN(n24452) );
  INV_X1 U17816 ( .A(n18886), .ZN(n24453) );
  INV_X1 U17817 ( .A(n18886), .ZN(n24454) );
  INV_X1 U17818 ( .A(n18887), .ZN(n24455) );
  INV_X1 U17819 ( .A(n18887), .ZN(n24456) );
  INV_X1 U17820 ( .A(n18888), .ZN(n24457) );
  INV_X1 U17821 ( .A(n18888), .ZN(n24458) );
  INV_X1 U17822 ( .A(n18889), .ZN(n24459) );
  INV_X1 U17823 ( .A(n18889), .ZN(n24460) );
  INV_X1 U17824 ( .A(n18890), .ZN(n24461) );
  INV_X1 U17825 ( .A(n18890), .ZN(n24462) );
  INV_X1 U17826 ( .A(n18891), .ZN(n24463) );
  INV_X1 U17827 ( .A(n18891), .ZN(n24464) );
  INV_X1 U17828 ( .A(n18892), .ZN(n24465) );
  INV_X1 U17829 ( .A(n18892), .ZN(n24466) );
  INV_X1 U17830 ( .A(n18893), .ZN(n24467) );
  INV_X1 U17831 ( .A(n18893), .ZN(n24468) );
  INV_X1 U17832 ( .A(n27207), .ZN(n24469) );
  INV_X1 U17833 ( .A(n24469), .ZN(n24470) );
  INV_X1 U17834 ( .A(n24469), .ZN(n24471) );
  INV_X1 U17835 ( .A(n26142), .ZN(n24472) );
  INV_X1 U17836 ( .A(n24472), .ZN(n24473) );
  INV_X1 U17837 ( .A(n24472), .ZN(n24474) );
  INV_X1 U17838 ( .A(n26138), .ZN(n24475) );
  INV_X1 U17839 ( .A(n24475), .ZN(n24476) );
  INV_X1 U17840 ( .A(n24475), .ZN(n24477) );
  INV_X1 U17841 ( .A(n27150), .ZN(n24478) );
  INV_X1 U17842 ( .A(n24478), .ZN(n24479) );
  INV_X1 U17843 ( .A(n24478), .ZN(n24480) );
  INV_X1 U17844 ( .A(n27272), .ZN(n24481) );
  INV_X1 U17845 ( .A(n24481), .ZN(n24482) );
  INV_X1 U17846 ( .A(n24481), .ZN(n24483) );
  INV_X1 U17847 ( .A(n18894), .ZN(n24484) );
  INV_X1 U17848 ( .A(n18894), .ZN(n24485) );
  INV_X1 U17849 ( .A(n18895), .ZN(n24486) );
  INV_X1 U17850 ( .A(n18895), .ZN(n24487) );
  INV_X1 U17851 ( .A(n18896), .ZN(n24488) );
  INV_X1 U17852 ( .A(n18896), .ZN(n24489) );
  INV_X1 U17853 ( .A(n18897), .ZN(n24490) );
  INV_X1 U17854 ( .A(n18897), .ZN(n24491) );
  INV_X1 U17855 ( .A(n18898), .ZN(n24492) );
  INV_X1 U17856 ( .A(n18898), .ZN(n24493) );
  INV_X1 U17857 ( .A(n18899), .ZN(n24494) );
  INV_X1 U17858 ( .A(n18899), .ZN(n24495) );
  INV_X1 U17859 ( .A(n18900), .ZN(n24496) );
  INV_X1 U17860 ( .A(n18900), .ZN(n24497) );
  INV_X1 U17861 ( .A(n27086), .ZN(n24498) );
  INV_X1 U17862 ( .A(n24498), .ZN(n24499) );
  INV_X1 U17863 ( .A(n24498), .ZN(n24500) );
  INV_X1 U17864 ( .A(n18901), .ZN(n24501) );
  INV_X1 U17865 ( .A(n18901), .ZN(n24502) );
  INV_X1 U17866 ( .A(n27002), .ZN(n24503) );
  INV_X1 U17867 ( .A(n24503), .ZN(n24504) );
  INV_X1 U17868 ( .A(n24503), .ZN(n24505) );
  INV_X1 U17869 ( .A(n18902), .ZN(n24506) );
  INV_X1 U17870 ( .A(n18902), .ZN(n24507) );
  INV_X1 U17871 ( .A(n27014), .ZN(n24508) );
  INV_X1 U17872 ( .A(n24508), .ZN(n24509) );
  INV_X1 U17873 ( .A(n24508), .ZN(n24510) );
  INV_X1 U17874 ( .A(n18903), .ZN(n24511) );
  INV_X1 U17875 ( .A(n19028), .ZN(n24512) );
  INV_X1 U17876 ( .A(n24512), .ZN(n24513) );
  INV_X1 U17877 ( .A(n24512), .ZN(n24514) );
  INV_X1 U17878 ( .A(n18904), .ZN(n24515) );
  INV_X1 U17879 ( .A(n18904), .ZN(n24516) );
  INV_X1 U17880 ( .A(n18905), .ZN(n24517) );
  INV_X1 U17881 ( .A(n18905), .ZN(n24518) );
  INV_X1 U17882 ( .A(n19024), .ZN(n24519) );
  INV_X1 U17883 ( .A(n24519), .ZN(n24520) );
  INV_X1 U17884 ( .A(n24519), .ZN(n24521) );
  INV_X1 U17885 ( .A(n18906), .ZN(n24522) );
  INV_X1 U17886 ( .A(n18906), .ZN(n24523) );
  INV_X1 U17887 ( .A(n18907), .ZN(n24524) );
  INV_X1 U17888 ( .A(n18907), .ZN(n24525) );
  INV_X1 U17889 ( .A(n18908), .ZN(n24526) );
  INV_X1 U17890 ( .A(n18908), .ZN(n24527) );
  INV_X1 U17891 ( .A(n18909), .ZN(n24528) );
  INV_X1 U17892 ( .A(n18909), .ZN(n24529) );
  INV_X1 U17893 ( .A(n18917), .ZN(n24530) );
  INV_X1 U17894 ( .A(n24530), .ZN(n24531) );
  INV_X1 U17895 ( .A(n24530), .ZN(n24532) );
  INV_X1 U17896 ( .A(n27242), .ZN(n24533) );
  INV_X1 U17897 ( .A(n24533), .ZN(n24534) );
  INV_X1 U17898 ( .A(n24533), .ZN(n24535) );
  INV_X1 U17899 ( .A(n18910), .ZN(n24536) );
  INV_X1 U17900 ( .A(n18910), .ZN(n24537) );
  INV_X1 U17901 ( .A(n27161), .ZN(n24538) );
  INV_X1 U17902 ( .A(n24538), .ZN(n24539) );
  INV_X1 U17903 ( .A(n24538), .ZN(n24540) );
  INV_X1 U17904 ( .A(n18911), .ZN(n24541) );
  INV_X1 U17905 ( .A(n18911), .ZN(n24542) );
  INV_X1 U17906 ( .A(n27249), .ZN(n24543) );
  INV_X1 U17907 ( .A(n24543), .ZN(n24544) );
  INV_X1 U17908 ( .A(n24543), .ZN(n24545) );
  INV_X1 U17909 ( .A(n27165), .ZN(n24546) );
  INV_X1 U17910 ( .A(n24546), .ZN(n24547) );
  INV_X1 U17911 ( .A(n24546), .ZN(n24548) );
  INV_X1 U17912 ( .A(n27164), .ZN(n24549) );
  INV_X1 U17913 ( .A(n24549), .ZN(n24550) );
  INV_X1 U17914 ( .A(n24549), .ZN(n24551) );
  INV_X1 U17915 ( .A(n18912), .ZN(n24552) );
  INV_X1 U17916 ( .A(n18912), .ZN(n24553) );
  INV_X1 U17917 ( .A(n27162), .ZN(n24554) );
  INV_X1 U17918 ( .A(n24554), .ZN(n24555) );
  INV_X1 U17919 ( .A(n24554), .ZN(n24556) );
  INV_X1 U17920 ( .A(n27161), .ZN(n24557) );
  INV_X1 U17921 ( .A(n24557), .ZN(n24558) );
  INV_X1 U17922 ( .A(n24557), .ZN(n24559) );
  INV_X1 U17923 ( .A(n27242), .ZN(n24560) );
  INV_X1 U17924 ( .A(n24560), .ZN(n24561) );
  INV_X1 U17925 ( .A(n24560), .ZN(n24562) );
  INV_X1 U17926 ( .A(n27253), .ZN(n24563) );
  INV_X1 U17927 ( .A(n24563), .ZN(n24564) );
  INV_X1 U17928 ( .A(n24563), .ZN(n24565) );
  INV_X1 U17929 ( .A(n27252), .ZN(n24566) );
  INV_X1 U17930 ( .A(n24566), .ZN(n24567) );
  INV_X1 U17931 ( .A(n24566), .ZN(n24568) );
  INV_X1 U17932 ( .A(n18913), .ZN(n24569) );
  INV_X1 U17933 ( .A(n18913), .ZN(n24570) );
  INV_X1 U17934 ( .A(n27250), .ZN(n24571) );
  INV_X1 U17935 ( .A(n24571), .ZN(n24572) );
  INV_X1 U17936 ( .A(n24571), .ZN(n24573) );
  INV_X1 U17937 ( .A(n27249), .ZN(n24574) );
  INV_X1 U17938 ( .A(n24574), .ZN(n24575) );
  INV_X1 U17939 ( .A(n24574), .ZN(n24576) );
  INV_X1 U17940 ( .A(n27170), .ZN(n24577) );
  INV_X1 U17941 ( .A(n24577), .ZN(n24578) );
  INV_X1 U17942 ( .A(n24577), .ZN(n24579) );
  INV_X1 U17943 ( .A(n27258), .ZN(n24580) );
  INV_X1 U17944 ( .A(n24580), .ZN(n24581) );
  INV_X1 U17945 ( .A(n24580), .ZN(n24582) );
  INV_X1 U17946 ( .A(n20493), .ZN(n24583) );
  INV_X1 U17947 ( .A(n20494), .ZN(n24584) );
  INV_X1 U17948 ( .A(n20488), .ZN(n24585) );
  INV_X1 U17949 ( .A(n20489), .ZN(n24586) );
  INV_X1 U17950 ( .A(n20494), .ZN(n24587) );
  INV_X1 U17951 ( .A(n27109), .ZN(n24588) );
  INV_X1 U17952 ( .A(n20489), .ZN(n24589) );
  INV_X1 U17953 ( .A(n27072), .ZN(n24590) );
  INV_X1 U17954 ( .A(n18914), .ZN(n24591) );
  INV_X1 U17955 ( .A(n18914), .ZN(n24592) );
  INV_X1 U17956 ( .A(n27049), .ZN(n24593) );
  INV_X1 U17957 ( .A(n24593), .ZN(n24594) );
  INV_X1 U17958 ( .A(n24593), .ZN(n24595) );
  INV_X1 U17959 ( .A(n18915), .ZN(n24596) );
  INV_X1 U17960 ( .A(n18915), .ZN(n24597) );
  INV_X1 U17961 ( .A(n27031), .ZN(n24598) );
  INV_X1 U17962 ( .A(n24598), .ZN(n24599) );
  INV_X1 U17963 ( .A(n24598), .ZN(n24600) );
  INV_X1 U17964 ( .A(n26939), .ZN(n24601) );
  INV_X1 U17965 ( .A(n24601), .ZN(n24602) );
  INV_X1 U17966 ( .A(n24601), .ZN(n24603) );
  INV_X1 U17967 ( .A(n27160), .ZN(n24604) );
  INV_X1 U17968 ( .A(n24604), .ZN(n24605) );
  INV_X1 U17969 ( .A(n24604), .ZN(n24606) );
  INV_X1 U17970 ( .A(n27160), .ZN(n24607) );
  INV_X1 U17971 ( .A(n24607), .ZN(n24608) );
  INV_X1 U17972 ( .A(n24607), .ZN(n24609) );
  INV_X1 U17973 ( .A(n27159), .ZN(n24610) );
  INV_X1 U17974 ( .A(n24610), .ZN(n24611) );
  INV_X1 U17975 ( .A(n24610), .ZN(n24612) );
  INV_X1 U17976 ( .A(n27159), .ZN(n24613) );
  INV_X1 U17977 ( .A(n24613), .ZN(n24614) );
  INV_X1 U17978 ( .A(n24613), .ZN(n24615) );
  INV_X1 U17979 ( .A(n18916), .ZN(n24616) );
  INV_X1 U17980 ( .A(n18916), .ZN(n24617) );
  INV_X1 U17981 ( .A(n18917), .ZN(n24618) );
  INV_X1 U17982 ( .A(n27248), .ZN(n24619) );
  INV_X1 U17983 ( .A(n24619), .ZN(n24620) );
  INV_X1 U17984 ( .A(n24619), .ZN(n24621) );
  INV_X1 U17985 ( .A(n27248), .ZN(n24622) );
  INV_X1 U17986 ( .A(n24622), .ZN(n24623) );
  INV_X1 U17987 ( .A(n24622), .ZN(n24624) );
  INV_X1 U17988 ( .A(n27247), .ZN(n24625) );
  INV_X1 U17989 ( .A(n24625), .ZN(n24626) );
  INV_X1 U17990 ( .A(n24625), .ZN(n24627) );
  INV_X1 U17991 ( .A(n27247), .ZN(n24628) );
  INV_X1 U17992 ( .A(n24628), .ZN(n24629) );
  INV_X1 U17993 ( .A(n24628), .ZN(n24630) );
  INV_X1 U17994 ( .A(n20889), .ZN(n24631) );
  INV_X1 U17995 ( .A(n24631), .ZN(n24632) );
  INV_X1 U17996 ( .A(n24631), .ZN(n24633) );
  INV_X1 U17997 ( .A(n26998), .ZN(n24634) );
  INV_X1 U17998 ( .A(n24634), .ZN(n24635) );
  INV_X1 U17999 ( .A(n24634), .ZN(n24636) );
  INV_X1 U18000 ( .A(n26999), .ZN(n24637) );
  INV_X1 U18001 ( .A(n24637), .ZN(n24638) );
  INV_X1 U18002 ( .A(n24637), .ZN(n24639) );
  INV_X1 U18003 ( .A(n27112), .ZN(n24640) );
  INV_X1 U18004 ( .A(n24640), .ZN(n24641) );
  INV_X1 U18005 ( .A(n24640), .ZN(n24642) );
  INV_X1 U18006 ( .A(n19108), .ZN(n24643) );
  INV_X1 U18007 ( .A(n24643), .ZN(n24644) );
  INV_X1 U18008 ( .A(n24643), .ZN(n24645) );
  INV_X1 U18009 ( .A(n19108), .ZN(n24646) );
  INV_X1 U18010 ( .A(n24646), .ZN(n24647) );
  INV_X1 U18011 ( .A(n24646), .ZN(n24648) );
  INV_X1 U18012 ( .A(n27111), .ZN(n24649) );
  INV_X1 U18013 ( .A(n24649), .ZN(n24650) );
  INV_X1 U18014 ( .A(n25378), .ZN(n24651) );
  INV_X1 U18015 ( .A(n25378), .ZN(n24652) );
  INV_X1 U18016 ( .A(n5133), .ZN(n24653) );
  INV_X1 U18017 ( .A(n24653), .ZN(n24654) );
  INV_X1 U18018 ( .A(n24653), .ZN(n24655) );
  INV_X1 U18019 ( .A(n18922), .ZN(n24656) );
  INV_X1 U18020 ( .A(n18922), .ZN(n24657) );
  INV_X1 U18021 ( .A(n19757), .ZN(n24658) );
  INV_X1 U18022 ( .A(n19318), .ZN(n24659) );
  INV_X1 U18023 ( .A(n26329), .ZN(n24660) );
  INV_X1 U18024 ( .A(n24660), .ZN(n24661) );
  INV_X1 U18025 ( .A(n24660), .ZN(n24662) );
  INV_X1 U18026 ( .A(n25646), .ZN(n24663) );
  INV_X1 U18027 ( .A(n24663), .ZN(n24664) );
  INV_X1 U18028 ( .A(n24663), .ZN(n24665) );
  INV_X1 U18029 ( .A(n26994), .ZN(n24666) );
  INV_X1 U18030 ( .A(n24666), .ZN(n24667) );
  INV_X1 U18031 ( .A(n24666), .ZN(n24668) );
  INV_X1 U18032 ( .A(n22969), .ZN(n24669) );
  INV_X1 U18033 ( .A(n24669), .ZN(n24670) );
  INV_X1 U18034 ( .A(n24669), .ZN(n24671) );
  INV_X1 U18035 ( .A(n22972), .ZN(n24672) );
  INV_X1 U18036 ( .A(n24672), .ZN(n24673) );
  INV_X1 U18037 ( .A(n24672), .ZN(n24674) );
  INV_X1 U18038 ( .A(n18923), .ZN(n24675) );
  INV_X1 U18039 ( .A(n18923), .ZN(n24676) );
  INV_X1 U18040 ( .A(n18924), .ZN(n24677) );
  INV_X1 U18041 ( .A(n18924), .ZN(n24678) );
  INV_X1 U18042 ( .A(n18925), .ZN(n24679) );
  INV_X1 U18043 ( .A(n18925), .ZN(n24680) );
  INV_X1 U18044 ( .A(n18926), .ZN(n24681) );
  INV_X1 U18045 ( .A(n18926), .ZN(n24682) );
  INV_X1 U18046 ( .A(n18927), .ZN(n24683) );
  INV_X1 U18047 ( .A(n18927), .ZN(n24684) );
  INV_X1 U18048 ( .A(n18928), .ZN(n24685) );
  INV_X1 U18049 ( .A(n18928), .ZN(n24686) );
  INV_X1 U18050 ( .A(n18929), .ZN(n24687) );
  INV_X1 U18051 ( .A(n18929), .ZN(n24688) );
  INV_X1 U18052 ( .A(n18930), .ZN(n24689) );
  INV_X1 U18053 ( .A(n18930), .ZN(n24690) );
  INV_X1 U18054 ( .A(n18931), .ZN(n24691) );
  INV_X1 U18055 ( .A(n18931), .ZN(n24692) );
  INV_X1 U18056 ( .A(n18932), .ZN(n24693) );
  INV_X1 U18057 ( .A(n18932), .ZN(n24694) );
  INV_X1 U18058 ( .A(n18933), .ZN(n24695) );
  INV_X1 U18059 ( .A(n18933), .ZN(n24696) );
  INV_X1 U18060 ( .A(n18934), .ZN(n24697) );
  INV_X1 U18061 ( .A(n18934), .ZN(n24698) );
  INV_X1 U18062 ( .A(n18935), .ZN(n24699) );
  INV_X1 U18063 ( .A(n18935), .ZN(n24700) );
  INV_X1 U18064 ( .A(n18936), .ZN(n24701) );
  INV_X1 U18065 ( .A(n18936), .ZN(n24702) );
  INV_X1 U18066 ( .A(n18937), .ZN(n24703) );
  INV_X1 U18067 ( .A(n18937), .ZN(n24704) );
  INV_X1 U18068 ( .A(n18938), .ZN(n24705) );
  INV_X1 U18069 ( .A(n18938), .ZN(n24706) );
  INV_X1 U18070 ( .A(n18939), .ZN(n24707) );
  INV_X1 U18071 ( .A(n18939), .ZN(n24708) );
  INV_X1 U18072 ( .A(n18940), .ZN(n24709) );
  INV_X1 U18073 ( .A(n18940), .ZN(n24710) );
  INV_X1 U18074 ( .A(n18941), .ZN(n24711) );
  INV_X1 U18075 ( .A(n18941), .ZN(n24712) );
  INV_X1 U18076 ( .A(n50780), .ZN(n24713) );
  INV_X1 U18077 ( .A(n24713), .ZN(n24714) );
  INV_X1 U18078 ( .A(n24713), .ZN(n24715) );
  INV_X1 U18079 ( .A(n44680), .ZN(n24716) );
  INV_X1 U18080 ( .A(n24716), .ZN(n24717) );
  INV_X1 U18081 ( .A(n24716), .ZN(n24718) );
  INV_X1 U18082 ( .A(n3483), .ZN(n24719) );
  INV_X1 U18083 ( .A(n24719), .ZN(n24720) );
  INV_X1 U18084 ( .A(n24719), .ZN(n24721) );
  INV_X1 U18085 ( .A(n18942), .ZN(n24722) );
  INV_X1 U18086 ( .A(n18942), .ZN(n24723) );
  INV_X1 U18087 ( .A(n18943), .ZN(n24724) );
  INV_X1 U18088 ( .A(n18943), .ZN(n24725) );
  INV_X1 U18089 ( .A(n18944), .ZN(n24726) );
  INV_X1 U18090 ( .A(n18944), .ZN(n24727) );
  INV_X1 U18091 ( .A(n4542), .ZN(n24728) );
  INV_X1 U18092 ( .A(n24728), .ZN(n24729) );
  INV_X1 U18093 ( .A(n21417), .ZN(n24730) );
  INV_X1 U18094 ( .A(n21420), .ZN(n24731) );
  INV_X1 U18095 ( .A(n27262), .ZN(n24732) );
  INV_X1 U18096 ( .A(n24732), .ZN(n24733) );
  INV_X1 U18097 ( .A(n27151), .ZN(n24734) );
  INV_X1 U18098 ( .A(n24734), .ZN(n24735) );
  INV_X1 U18099 ( .A(n26651), .ZN(n24736) );
  INV_X1 U18100 ( .A(n24736), .ZN(n24737) );
  INV_X1 U18101 ( .A(n24740), .ZN(n24738) );
  INV_X1 U18102 ( .A(n24742), .ZN(n24739) );
  INV_X1 U18103 ( .A(n27126), .ZN(n24740) );
  INV_X1 U18104 ( .A(n24740), .ZN(n24741) );
  INV_X1 U18105 ( .A(n27274), .ZN(n24742) );
  INV_X1 U18106 ( .A(n24742), .ZN(n24743) );
  INV_X1 U18107 ( .A(n18946), .ZN(n24744) );
  INV_X1 U18108 ( .A(n27028), .ZN(n24745) );
  INV_X1 U18109 ( .A(n24745), .ZN(n24746) );
  INV_X1 U18110 ( .A(n24745), .ZN(n24747) );
  INV_X1 U18111 ( .A(n18947), .ZN(n24748) );
  INV_X1 U18112 ( .A(n18948), .ZN(n24749) );
  INV_X1 U18113 ( .A(n24700), .ZN(n24750) );
  INV_X1 U18114 ( .A(n24750), .ZN(n24751) );
  CLKBUF_X1 U18115 ( .A(n22891), .Z(n24752) );
  INV_X1 U18116 ( .A(n24486), .ZN(n24753) );
  INV_X1 U18117 ( .A(n24753), .ZN(n24754) );
  CLKBUF_X1 U18118 ( .A(n24744), .Z(n27220) );
  INV_X1 U18119 ( .A(n27220), .ZN(n24755) );
  INV_X1 U18120 ( .A(n27220), .ZN(n24756) );
  INV_X1 U18121 ( .A(n24707), .ZN(n24757) );
  INV_X1 U18122 ( .A(n24759), .ZN(n24758) );
  INV_X1 U18123 ( .A(n27197), .ZN(n24759) );
  INV_X1 U18124 ( .A(n24759), .ZN(n24760) );
  INV_X1 U18125 ( .A(n19236), .ZN(n24761) );
  INV_X1 U18126 ( .A(n24761), .ZN(n24762) );
  INV_X1 U18127 ( .A(n19235), .ZN(n24763) );
  INV_X1 U18128 ( .A(n24763), .ZN(n24764) );
  INV_X1 U18129 ( .A(n27265), .ZN(n24765) );
  INV_X1 U18130 ( .A(n24765), .ZN(n24766) );
  INV_X1 U18131 ( .A(n27264), .ZN(n24767) );
  INV_X1 U18132 ( .A(n24767), .ZN(n24768) );
  INV_X1 U18133 ( .A(n24767), .ZN(n24769) );
  INV_X1 U18134 ( .A(n27155), .ZN(n24770) );
  INV_X1 U18135 ( .A(n24770), .ZN(n24771) );
  INV_X1 U18136 ( .A(n27154), .ZN(n24772) );
  INV_X1 U18137 ( .A(n24772), .ZN(n24773) );
  INV_X1 U18138 ( .A(n24772), .ZN(n24774) );
  INV_X1 U18139 ( .A(n27209), .ZN(n24775) );
  INV_X1 U18140 ( .A(n24775), .ZN(n24776) );
  INV_X1 U18141 ( .A(n25875), .ZN(n24777) );
  INV_X1 U18142 ( .A(n24777), .ZN(n24778) );
  INV_X1 U18143 ( .A(n25873), .ZN(n24779) );
  INV_X1 U18144 ( .A(n24779), .ZN(n24780) );
  INV_X1 U18145 ( .A(n27208), .ZN(n24781) );
  INV_X1 U18146 ( .A(n24781), .ZN(n24782) );
  INV_X1 U18147 ( .A(n24781), .ZN(n24783) );
  INV_X1 U18148 ( .A(n22883), .ZN(n24784) );
  INV_X1 U18149 ( .A(n24784), .ZN(n24785) );
  CLKBUF_X1 U18150 ( .A(n19313), .Z(n24786) );
  INV_X1 U18151 ( .A(n24790), .ZN(n24787) );
  INV_X1 U18152 ( .A(n24787), .ZN(n24788) );
  CLKBUF_X1 U18153 ( .A(n24790), .Z(n24789) );
  CLKBUF_X1 U18154 ( .A(n24708), .Z(n24790) );
  CLKBUF_X1 U18155 ( .A(n24758), .Z(n27198) );
  INV_X1 U18156 ( .A(n27198), .ZN(n24791) );
  INV_X1 U18157 ( .A(n27198), .ZN(n24792) );
  INV_X1 U18158 ( .A(n18951), .ZN(n24793) );
  INV_X1 U18159 ( .A(n18951), .ZN(n24794) );
  INV_X1 U18160 ( .A(n259901), .ZN(n24795) );
  INV_X1 U18161 ( .A(n24795), .ZN(n24796) );
  INV_X1 U18162 ( .A(n24704), .ZN(n24797) );
  INV_X1 U18163 ( .A(n24797), .ZN(n24798) );
  INV_X1 U18164 ( .A(n24710), .ZN(n24799) );
  INV_X1 U18165 ( .A(n24799), .ZN(n24800) );
  INV_X1 U18166 ( .A(n18952), .ZN(n24801) );
  INV_X1 U18167 ( .A(n18953), .ZN(n24802) );
  INV_X1 U18168 ( .A(n25994), .ZN(n24803) );
  INV_X1 U18169 ( .A(n24803), .ZN(n24804) );
  INV_X1 U18170 ( .A(n26158), .ZN(n24805) );
  INV_X1 U18171 ( .A(n24805), .ZN(n24806) );
  INV_X1 U18172 ( .A(n26149), .ZN(n24807) );
  INV_X1 U18173 ( .A(n24807), .ZN(n24808) );
  INV_X1 U18174 ( .A(n18954), .ZN(n24809) );
  INV_X1 U18175 ( .A(n4542), .ZN(n24810) );
  INV_X1 U18176 ( .A(n24729), .ZN(n24811) );
  INV_X1 U18177 ( .A(n26939), .ZN(n24812) );
  INV_X1 U18178 ( .A(n24812), .ZN(n24813) );
  INV_X1 U18179 ( .A(n18955), .ZN(n24814) );
  INV_X1 U18180 ( .A(n18956), .ZN(n24815) );
  INV_X1 U18181 ( .A(n26937), .ZN(n24816) );
  INV_X1 U18182 ( .A(n24816), .ZN(n24817) );
  INV_X1 U18183 ( .A(n18957), .ZN(n24818) );
  INV_X1 U18184 ( .A(n18958), .ZN(n24819) );
  INV_X1 U18185 ( .A(n22877), .ZN(n24820) );
  INV_X1 U18186 ( .A(n24820), .ZN(n24821) );
  INV_X1 U18187 ( .A(n18959), .ZN(n24822) );
  INV_X1 U18188 ( .A(n17094), .ZN(n24823) );
  INV_X1 U18189 ( .A(n18960), .ZN(n24824) );
  INV_X1 U18190 ( .A(n18961), .ZN(n24825) );
  INV_X1 U18191 ( .A(n18962), .ZN(n24826) );
  INV_X1 U18192 ( .A(n17093), .ZN(n24827) );
  INV_X1 U18193 ( .A(n18963), .ZN(n24828) );
  INV_X1 U18194 ( .A(n18964), .ZN(n24829) );
  INV_X1 U18195 ( .A(n17092), .ZN(n24830) );
  INV_X1 U18196 ( .A(n18965), .ZN(n24831) );
  INV_X1 U18197 ( .A(n18966), .ZN(n24832) );
  INV_X1 U18198 ( .A(n18966), .ZN(n24833) );
  INV_X1 U18199 ( .A(n18967), .ZN(n24834) );
  INV_X1 U18200 ( .A(n17091), .ZN(n24835) );
  INV_X1 U18201 ( .A(n18968), .ZN(n24836) );
  INV_X1 U18202 ( .A(n18969), .ZN(n24837) );
  INV_X1 U18203 ( .A(n18970), .ZN(n24838) );
  INV_X1 U18204 ( .A(n79), .ZN(n24839) );
  INV_X1 U18205 ( .A(n78), .ZN(n24840) );
  INV_X1 U18206 ( .A(n18971), .ZN(n24841) );
  INV_X1 U18207 ( .A(n18972), .ZN(n24842) );
  INV_X1 U18208 ( .A(n18973), .ZN(n24843) );
  INV_X1 U18209 ( .A(n77), .ZN(n24844) );
  INV_X1 U18210 ( .A(n18974), .ZN(n24845) );
  INV_X1 U18211 ( .A(n18975), .ZN(n24846) );
  INV_X1 U18212 ( .A(n76), .ZN(n24847) );
  INV_X1 U18213 ( .A(n18976), .ZN(n24848) );
  INV_X1 U18214 ( .A(n75), .ZN(n24849) );
  INV_X1 U18215 ( .A(n18977), .ZN(n24850) );
  INV_X1 U18216 ( .A(n74), .ZN(n24851) );
  INV_X1 U18217 ( .A(n18978), .ZN(n24852) );
  INV_X1 U18218 ( .A(n18979), .ZN(n24853) );
  INV_X1 U18219 ( .A(n18980), .ZN(n24854) );
  INV_X1 U18220 ( .A(n73), .ZN(n24855) );
  INV_X1 U18221 ( .A(n18981), .ZN(n24856) );
  INV_X1 U18222 ( .A(n18982), .ZN(n24857) );
  INV_X1 U18223 ( .A(n26992), .ZN(n24858) );
  INV_X1 U18224 ( .A(n18983), .ZN(n24859) );
  INV_X1 U18225 ( .A(n26866), .ZN(n24860) );
  INV_X1 U18226 ( .A(n24860), .ZN(n24861) );
  INV_X1 U18227 ( .A(n26903), .ZN(n24862) );
  INV_X1 U18228 ( .A(n24862), .ZN(n24863) );
  INV_X1 U18229 ( .A(n24862), .ZN(n24864) );
  INV_X1 U18230 ( .A(n26841), .ZN(n24865) );
  INV_X1 U18231 ( .A(n24865), .ZN(n24866) );
  INV_X1 U18232 ( .A(n26845), .ZN(n24867) );
  INV_X1 U18233 ( .A(n24867), .ZN(n24868) );
  INV_X1 U18234 ( .A(n26841), .ZN(n24869) );
  INV_X1 U18235 ( .A(n24869), .ZN(n24870) );
  INV_X1 U18236 ( .A(n26845), .ZN(n24871) );
  INV_X1 U18237 ( .A(n24871), .ZN(n24872) );
  INV_X1 U18238 ( .A(n26803), .ZN(n24873) );
  INV_X1 U18239 ( .A(n24873), .ZN(n24874) );
  INV_X1 U18240 ( .A(n24873), .ZN(n24875) );
  INV_X1 U18241 ( .A(n26806), .ZN(n24876) );
  INV_X1 U18242 ( .A(n24876), .ZN(n24877) );
  INV_X1 U18243 ( .A(n26797), .ZN(n24878) );
  INV_X1 U18244 ( .A(n24878), .ZN(n24879) );
  INV_X1 U18245 ( .A(n24878), .ZN(n24880) );
  INV_X1 U18246 ( .A(n26803), .ZN(n24881) );
  INV_X1 U18247 ( .A(n24881), .ZN(n24882) );
  INV_X1 U18248 ( .A(n24881), .ZN(n24883) );
  INV_X1 U18249 ( .A(n26797), .ZN(n24884) );
  INV_X1 U18250 ( .A(n24884), .ZN(n24885) );
  INV_X1 U18251 ( .A(n24884), .ZN(n24886) );
  INV_X1 U18252 ( .A(n26793), .ZN(n24887) );
  INV_X1 U18253 ( .A(n24887), .ZN(n24888) );
  INV_X1 U18254 ( .A(n26782), .ZN(n24889) );
  INV_X1 U18255 ( .A(n24889), .ZN(n24890) );
  INV_X1 U18256 ( .A(n24889), .ZN(n24891) );
  INV_X1 U18257 ( .A(n26786), .ZN(n24892) );
  INV_X1 U18258 ( .A(n24892), .ZN(n24893) );
  INV_X1 U18259 ( .A(n18984), .ZN(n24894) );
  INV_X1 U18260 ( .A(n26765), .ZN(n24895) );
  INV_X1 U18261 ( .A(n24895), .ZN(n24896) );
  INV_X1 U18262 ( .A(n26767), .ZN(n24897) );
  INV_X1 U18263 ( .A(n24897), .ZN(n24898) );
  INV_X1 U18264 ( .A(n26771), .ZN(n24899) );
  INV_X1 U18265 ( .A(n24899), .ZN(n24900) );
  INV_X1 U18266 ( .A(n26771), .ZN(n24901) );
  INV_X1 U18267 ( .A(n24901), .ZN(n24902) );
  INV_X1 U18268 ( .A(n26759), .ZN(n24903) );
  INV_X1 U18269 ( .A(n24903), .ZN(n24904) );
  INV_X1 U18270 ( .A(n26767), .ZN(n24905) );
  INV_X1 U18271 ( .A(n24905), .ZN(n24906) );
  INV_X1 U18272 ( .A(n25160), .ZN(n24907) );
  INV_X1 U18273 ( .A(n25142), .ZN(n24908) );
  INV_X1 U18274 ( .A(n26765), .ZN(n24909) );
  INV_X1 U18275 ( .A(n24909), .ZN(n24910) );
  INV_X1 U18276 ( .A(n26759), .ZN(n24911) );
  INV_X1 U18277 ( .A(n24911), .ZN(n24912) );
  INV_X1 U18278 ( .A(n26988), .ZN(n24913) );
  INV_X1 U18279 ( .A(n24913), .ZN(n24914) );
  INV_X1 U18280 ( .A(n24913), .ZN(n24915) );
  INV_X1 U18281 ( .A(n19016), .ZN(n24916) );
  INV_X1 U18282 ( .A(n24916), .ZN(n24917) );
  INV_X1 U18283 ( .A(n18988), .ZN(n24918) );
  INV_X1 U18284 ( .A(n18989), .ZN(n24919) );
  INV_X1 U18285 ( .A(n18989), .ZN(n24920) );
  CLKBUF_X1 U18286 ( .A(n26715), .Z(n24921) );
  INV_X1 U18287 ( .A(n18990), .ZN(n24922) );
  INV_X1 U18288 ( .A(n18990), .ZN(n24923) );
  CLKBUF_X1 U18289 ( .A(n22789), .Z(n26713) );
  INV_X1 U18290 ( .A(n26713), .ZN(n24924) );
  INV_X1 U18291 ( .A(n26713), .ZN(n24925) );
  INV_X1 U18292 ( .A(n24165), .ZN(n24926) );
  INV_X1 U18293 ( .A(n24926), .ZN(n24927) );
  INV_X1 U18294 ( .A(n24926), .ZN(n24928) );
  CLKBUF_X1 U18295 ( .A(n24932), .Z(n24929) );
  INV_X1 U18296 ( .A(n19301), .ZN(n24930) );
  INV_X1 U18297 ( .A(n24930), .ZN(n24931) );
  INV_X1 U18298 ( .A(n24930), .ZN(n24932) );
  CLKBUF_X1 U18299 ( .A(n22783), .Z(n26709) );
  INV_X1 U18300 ( .A(n26709), .ZN(n24933) );
  INV_X1 U18301 ( .A(n26709), .ZN(n24934) );
  INV_X1 U18302 ( .A(n24161), .ZN(n24935) );
  INV_X1 U18303 ( .A(n24935), .ZN(n24936) );
  INV_X1 U18304 ( .A(n24935), .ZN(n24937) );
  CLKBUF_X1 U18305 ( .A(n22781), .Z(n26706) );
  INV_X1 U18306 ( .A(n26706), .ZN(n24938) );
  INV_X1 U18307 ( .A(n26706), .ZN(n24939) );
  INV_X1 U18308 ( .A(n24157), .ZN(n24940) );
  INV_X1 U18309 ( .A(n24940), .ZN(n24941) );
  INV_X1 U18310 ( .A(n24940), .ZN(n24942) );
  CLKBUF_X1 U18311 ( .A(n26700), .Z(n24943) );
  CLKBUF_X1 U18312 ( .A(n22779), .Z(n26703) );
  INV_X1 U18313 ( .A(n26703), .ZN(n24944) );
  INV_X1 U18314 ( .A(n26703), .ZN(n24945) );
  INV_X1 U18315 ( .A(n22776), .ZN(n24946) );
  INV_X1 U18316 ( .A(n24946), .ZN(n24947) );
  INV_X1 U18317 ( .A(n26700), .ZN(n24948) );
  INV_X1 U18318 ( .A(n24948), .ZN(n24949) );
  INV_X1 U18319 ( .A(n22773), .ZN(n24950) );
  INV_X1 U18320 ( .A(n24950), .ZN(n24951) );
  CLKBUF_X1 U18321 ( .A(n26694), .Z(n24952) );
  INV_X1 U18322 ( .A(n26691), .ZN(n24953) );
  INV_X1 U18323 ( .A(n24953), .ZN(n24954) );
  INV_X1 U18324 ( .A(n22769), .ZN(n24955) );
  INV_X1 U18325 ( .A(n24955), .ZN(n24956) );
  INV_X1 U18326 ( .A(n26694), .ZN(n24957) );
  INV_X1 U18327 ( .A(n24957), .ZN(n24958) );
  CLKBUF_X1 U18328 ( .A(n26684), .Z(n24959) );
  INV_X1 U18329 ( .A(n26682), .ZN(n24960) );
  INV_X1 U18330 ( .A(n24960), .ZN(n24961) );
  INV_X1 U18331 ( .A(n26684), .ZN(n24962) );
  INV_X1 U18332 ( .A(n24962), .ZN(n24963) );
  INV_X1 U18333 ( .A(n22759), .ZN(n24964) );
  INV_X1 U18334 ( .A(n24964), .ZN(n24965) );
  CLKBUF_X1 U18335 ( .A(n26680), .Z(n24966) );
  INV_X1 U18336 ( .A(n22756), .ZN(n24967) );
  INV_X1 U18337 ( .A(n24967), .ZN(n24968) );
  INV_X1 U18338 ( .A(n26680), .ZN(n24969) );
  INV_X1 U18339 ( .A(n24969), .ZN(n24970) );
  INV_X1 U18340 ( .A(n72), .ZN(n24971) );
  INV_X1 U18341 ( .A(n26676), .ZN(n24972) );
  INV_X1 U18342 ( .A(n24972), .ZN(n24973) );
  INV_X1 U18343 ( .A(n71), .ZN(n24974) );
  INV_X1 U18344 ( .A(n18991), .ZN(n24975) );
  INV_X1 U18345 ( .A(n18992), .ZN(n24976) );
  INV_X1 U18346 ( .A(n18993), .ZN(n24977) );
  INV_X1 U18347 ( .A(n18994), .ZN(n24978) );
  INV_X1 U18348 ( .A(n18995), .ZN(n24979) );
  INV_X1 U18349 ( .A(n18996), .ZN(n24980) );
  INV_X1 U18350 ( .A(n18997), .ZN(n24981) );
  INV_X1 U18351 ( .A(n18998), .ZN(n24982) );
  INV_X1 U18352 ( .A(n18999), .ZN(n24983) );
  INV_X1 U18353 ( .A(n24103), .ZN(n24984) );
  INV_X1 U18354 ( .A(n24984), .ZN(n24985) );
  INV_X1 U18355 ( .A(n26670), .ZN(n24986) );
  INV_X1 U18356 ( .A(n24986), .ZN(n24987) );
  INV_X1 U18357 ( .A(n22748), .ZN(n24988) );
  INV_X1 U18358 ( .A(n24988), .ZN(n24989) );
  INV_X1 U18359 ( .A(n26664), .ZN(n24990) );
  INV_X1 U18360 ( .A(n24990), .ZN(n24991) );
  INV_X1 U18361 ( .A(n19291), .ZN(n24992) );
  INV_X1 U18362 ( .A(n24992), .ZN(n24993) );
  INV_X1 U18363 ( .A(n24992), .ZN(n24994) );
  INV_X1 U18364 ( .A(n24076), .ZN(n24995) );
  INV_X1 U18365 ( .A(n24995), .ZN(n24996) );
  INV_X1 U18366 ( .A(n19000), .ZN(n24997) );
  INV_X1 U18367 ( .A(n21403), .ZN(n24998) );
  INV_X1 U18368 ( .A(n24998), .ZN(n24999) );
  INV_X1 U18369 ( .A(n22725), .ZN(n25000) );
  INV_X1 U18370 ( .A(n25000), .ZN(n25001) );
  INV_X1 U18371 ( .A(n25000), .ZN(n25002) );
  INV_X1 U18372 ( .A(n24067), .ZN(n25003) );
  INV_X1 U18373 ( .A(n25003), .ZN(n25004) );
  INV_X1 U18374 ( .A(n26651), .ZN(n25005) );
  INV_X1 U18375 ( .A(n25005), .ZN(n25006) );
  INV_X1 U18376 ( .A(n24057), .ZN(n25007) );
  INV_X1 U18377 ( .A(n25007), .ZN(n25008) );
  INV_X1 U18378 ( .A(n24062), .ZN(n25009) );
  INV_X1 U18379 ( .A(n25009), .ZN(n25010) );
  INV_X1 U18380 ( .A(n27262), .ZN(n25011) );
  INV_X1 U18381 ( .A(n25011), .ZN(n25012) );
  INV_X1 U18382 ( .A(n25304), .ZN(n25013) );
  CLKBUF_X1 U18383 ( .A(n22691), .Z(n25014) );
  INV_X1 U18384 ( .A(n26923), .ZN(n25015) );
  INV_X1 U18385 ( .A(n25015), .ZN(n25016) );
  INV_X1 U18386 ( .A(n25015), .ZN(n25017) );
  INV_X1 U18387 ( .A(n25296), .ZN(n25018) );
  CLKBUF_X1 U18388 ( .A(n22685), .Z(n25019) );
  INV_X1 U18389 ( .A(n26924), .ZN(n25020) );
  INV_X1 U18390 ( .A(n25020), .ZN(n25021) );
  INV_X1 U18391 ( .A(n25020), .ZN(n25022) );
  INV_X1 U18392 ( .A(n19001), .ZN(n25023) );
  CLKBUF_X1 U18393 ( .A(n24822), .Z(n26617) );
  INV_X1 U18394 ( .A(n26617), .ZN(n25024) );
  INV_X1 U18395 ( .A(n26617), .ZN(n25025) );
  CLKBUF_X1 U18396 ( .A(n25023), .Z(n26615) );
  INV_X1 U18397 ( .A(n26615), .ZN(n25026) );
  INV_X1 U18398 ( .A(n26615), .ZN(n25027) );
  INV_X1 U18399 ( .A(n26616), .ZN(n25028) );
  INV_X1 U18400 ( .A(n25028), .ZN(n25029) );
  INV_X1 U18401 ( .A(n26603), .ZN(n25030) );
  INV_X1 U18402 ( .A(n25030), .ZN(n25031) );
  INV_X1 U18403 ( .A(n25026), .ZN(n25032) );
  INV_X1 U18404 ( .A(n25032), .ZN(n25033) );
  INV_X1 U18405 ( .A(n19002), .ZN(n25034) );
  INV_X1 U18406 ( .A(n19003), .ZN(n25035) );
  INV_X1 U18407 ( .A(n19004), .ZN(n25036) );
  INV_X1 U18408 ( .A(n26602), .ZN(n25037) );
  INV_X1 U18409 ( .A(n25037), .ZN(n25038) );
  INV_X1 U18410 ( .A(n26601), .ZN(n25039) );
  INV_X1 U18411 ( .A(n25039), .ZN(n25040) );
  INV_X1 U18412 ( .A(n19005), .ZN(n25041) );
  INV_X1 U18413 ( .A(n19006), .ZN(n25042) );
  INV_X1 U18414 ( .A(n19007), .ZN(n25043) );
  INV_X1 U18415 ( .A(n19008), .ZN(n25044) );
  INV_X1 U18416 ( .A(n26600), .ZN(n25045) );
  INV_X1 U18417 ( .A(n25045), .ZN(n25046) );
  INV_X1 U18418 ( .A(n26599), .ZN(n25047) );
  INV_X1 U18419 ( .A(n25047), .ZN(n25048) );
  INV_X1 U18420 ( .A(n19009), .ZN(n25049) );
  INV_X1 U18421 ( .A(n19010), .ZN(n25050) );
  INV_X1 U18422 ( .A(n19011), .ZN(n25051) );
  INV_X1 U18423 ( .A(n19012), .ZN(n25052) );
  INV_X1 U18424 ( .A(n26598), .ZN(n25053) );
  INV_X1 U18425 ( .A(n25053), .ZN(n25054) );
  INV_X1 U18426 ( .A(n26597), .ZN(n25055) );
  INV_X1 U18427 ( .A(n25055), .ZN(n25056) );
  INV_X1 U18428 ( .A(n19013), .ZN(n25057) );
  INV_X1 U18429 ( .A(n19014), .ZN(n25058) );
  INV_X1 U18430 ( .A(n19015), .ZN(n25059) );
  INV_X1 U18431 ( .A(n25285), .ZN(n25060) );
  INV_X1 U18432 ( .A(n22531), .ZN(n25061) );
  INV_X1 U18433 ( .A(n26596), .ZN(n25062) );
  INV_X1 U18434 ( .A(n25062), .ZN(n25063) );
  INV_X1 U18435 ( .A(n26590), .ZN(n25064) );
  INV_X1 U18436 ( .A(n25064), .ZN(n25065) );
  INV_X1 U18437 ( .A(n18853), .ZN(n25066) );
  INV_X1 U18438 ( .A(n26385), .ZN(n25067) );
  INV_X1 U18439 ( .A(n25067), .ZN(n25068) );
  INV_X1 U18440 ( .A(n26942), .ZN(n25069) );
  INV_X1 U18441 ( .A(n25069), .ZN(n25070) );
  INV_X1 U18442 ( .A(n26384), .ZN(n25071) );
  INV_X1 U18443 ( .A(n25071), .ZN(n25072) );
  INV_X1 U18444 ( .A(n26385), .ZN(n25073) );
  INV_X1 U18445 ( .A(n25073), .ZN(n25074) );
  INV_X1 U18446 ( .A(n26158), .ZN(n25075) );
  INV_X1 U18447 ( .A(n25075), .ZN(n25076) );
  INV_X1 U18448 ( .A(n26384), .ZN(n25077) );
  INV_X1 U18449 ( .A(n25077), .ZN(n25078) );
  INV_X1 U18450 ( .A(n25978), .ZN(n25079) );
  INV_X1 U18451 ( .A(n25079), .ZN(n25080) );
  INV_X1 U18452 ( .A(n26149), .ZN(n25081) );
  INV_X1 U18453 ( .A(n25081), .ZN(n25082) );
  INV_X1 U18454 ( .A(n259701), .ZN(n25083) );
  INV_X1 U18455 ( .A(n25083), .ZN(n25084) );
  INV_X1 U18456 ( .A(n19017), .ZN(n25085) );
  INV_X1 U18457 ( .A(n19017), .ZN(n25086) );
  INV_X1 U18458 ( .A(n19018), .ZN(n25087) );
  INV_X1 U18459 ( .A(n19019), .ZN(n25088) );
  INV_X1 U18460 ( .A(n19019), .ZN(n25089) );
  XNOR2_X1 U18461 ( .A(n539), .B(n24679), .ZN(r899_B_7_) );
  NOR3_X1 U18462 ( .A1(n539), .A2(n465), .A3(n24679), .ZN(r899_B_9_) );
  INV_X1 U18463 ( .A(n20909), .ZN(n25090) );
  INV_X1 U18464 ( .A(n20909), .ZN(n25091) );
  INV_X1 U18465 ( .A(n26992), .ZN(n25092) );
  INV_X1 U18466 ( .A(n20911), .ZN(n25093) );
  INV_X1 U18467 ( .A(n20911), .ZN(n25094) );
  INV_X1 U18468 ( .A(n20912), .ZN(n25095) );
  INV_X1 U18469 ( .A(n20912), .ZN(n25096) );
  INV_X1 U18470 ( .A(n20913), .ZN(n25097) );
  INV_X1 U18471 ( .A(n20913), .ZN(n25098) );
  INV_X1 U18472 ( .A(n20915), .ZN(n25099) );
  INV_X1 U18473 ( .A(n20915), .ZN(n25100) );
  INV_X1 U18474 ( .A(n20916), .ZN(n25101) );
  INV_X1 U18475 ( .A(n20916), .ZN(n25102) );
  INV_X1 U18476 ( .A(n20917), .ZN(n25103) );
  INV_X1 U18477 ( .A(n20917), .ZN(n25104) );
  INV_X1 U18478 ( .A(n20919), .ZN(n25105) );
  INV_X1 U18479 ( .A(n20919), .ZN(n25106) );
  INV_X1 U18480 ( .A(n22945), .ZN(n25107) );
  INV_X1 U18481 ( .A(n21410), .ZN(n25108) );
  INV_X1 U18482 ( .A(n25107), .ZN(n25109) );
  INV_X1 U18483 ( .A(n25107), .ZN(n25110) );
  INV_X1 U18484 ( .A(n20920), .ZN(n25111) );
  INV_X1 U18485 ( .A(n20924), .ZN(n25112) );
  INV_X1 U18486 ( .A(n20924), .ZN(n25113) );
  INV_X1 U18487 ( .A(n20925), .ZN(n25114) );
  INV_X1 U18488 ( .A(n20928), .ZN(n25115) );
  INV_X1 U18489 ( .A(n20928), .ZN(n25116) );
  INV_X1 U18490 ( .A(n20929), .ZN(n25117) );
  INV_X1 U18491 ( .A(n20929), .ZN(n25118) );
  INV_X1 U18492 ( .A(n20930), .ZN(n25119) );
  INV_X1 U18493 ( .A(n20930), .ZN(n25120) );
  INV_X1 U18494 ( .A(n20931), .ZN(n25121) );
  INV_X1 U18495 ( .A(n20931), .ZN(n25122) );
  INV_X1 U18496 ( .A(n20932), .ZN(n25123) );
  INV_X1 U18497 ( .A(n20932), .ZN(n25124) );
  INV_X1 U18498 ( .A(n20933), .ZN(n25125) );
  INV_X1 U18499 ( .A(n20933), .ZN(n25126) );
  INV_X1 U18500 ( .A(n27228), .ZN(n25127) );
  INV_X1 U18501 ( .A(n20940), .ZN(n25128) );
  INV_X1 U18502 ( .A(n25127), .ZN(n25129) );
  INV_X1 U18503 ( .A(n20937), .ZN(n25130) );
  INV_X1 U18504 ( .A(n20934), .ZN(n25131) );
  INV_X1 U18505 ( .A(n20934), .ZN(n25132) );
  INV_X1 U18506 ( .A(n26320), .ZN(n25133) );
  INV_X1 U18507 ( .A(n20936), .ZN(n25134) );
  INV_X1 U18508 ( .A(n20936), .ZN(n25135) );
  INV_X1 U18509 ( .A(n20937), .ZN(n25136) );
  INV_X1 U18510 ( .A(n20939), .ZN(n25137) );
  INV_X1 U18511 ( .A(n20939), .ZN(n25138) );
  INV_X1 U18512 ( .A(n20940), .ZN(n25139) );
  INV_X1 U18513 ( .A(n20941), .ZN(n25140) );
  INV_X1 U18514 ( .A(n20941), .ZN(n25141) );
  INV_X1 U18515 ( .A(n27225), .ZN(n25142) );
  INV_X1 U18516 ( .A(n20943), .ZN(n25143) );
  INV_X1 U18517 ( .A(n20943), .ZN(n25144) );
  INV_X1 U18518 ( .A(n27174), .ZN(n25145) );
  INV_X1 U18519 ( .A(n20950), .ZN(n25146) );
  INV_X1 U18520 ( .A(n25145), .ZN(n25147) );
  INV_X1 U18521 ( .A(n20947), .ZN(n25148) );
  INV_X1 U18522 ( .A(n20944), .ZN(n25149) );
  INV_X1 U18523 ( .A(n20944), .ZN(n25150) );
  INV_X1 U18524 ( .A(n26319), .ZN(n25151) );
  INV_X1 U18525 ( .A(n20946), .ZN(n25152) );
  INV_X1 U18526 ( .A(n20946), .ZN(n25153) );
  INV_X1 U18527 ( .A(n20947), .ZN(n25154) );
  INV_X1 U18528 ( .A(n20949), .ZN(n25155) );
  INV_X1 U18529 ( .A(n20949), .ZN(n25156) );
  INV_X1 U18530 ( .A(n20950), .ZN(n25157) );
  INV_X1 U18531 ( .A(n20951), .ZN(n25158) );
  INV_X1 U18532 ( .A(n20951), .ZN(n25159) );
  INV_X1 U18533 ( .A(n27172), .ZN(n25160) );
  INV_X1 U18534 ( .A(n20953), .ZN(n25161) );
  INV_X1 U18535 ( .A(n20953), .ZN(n25162) );
  INV_X1 U18536 ( .A(n20954), .ZN(n25163) );
  INV_X1 U18537 ( .A(n20954), .ZN(n25164) );
  CLKBUF_X1 U18538 ( .A(n24620), .Z(n27257) );
  INV_X1 U18539 ( .A(n27257), .ZN(n25165) );
  INV_X1 U18540 ( .A(n27257), .ZN(n25166) );
  INV_X1 U18541 ( .A(n20955), .ZN(n25167) );
  INV_X1 U18542 ( .A(n20955), .ZN(n25168) );
  CLKBUF_X1 U18543 ( .A(n24605), .Z(n27169) );
  INV_X1 U18544 ( .A(n27169), .ZN(n25169) );
  INV_X1 U18545 ( .A(n27169), .ZN(n25170) );
  INV_X1 U18546 ( .A(n20956), .ZN(n25171) );
  INV_X1 U18547 ( .A(n20956), .ZN(n25172) );
  CLKBUF_X1 U18548 ( .A(n24623), .Z(n27254) );
  INV_X1 U18549 ( .A(n27254), .ZN(n25173) );
  INV_X1 U18550 ( .A(n27254), .ZN(n25174) );
  CLKBUF_X1 U18551 ( .A(n24608), .Z(n27166) );
  INV_X1 U18552 ( .A(n27166), .ZN(n25175) );
  INV_X1 U18553 ( .A(n27166), .ZN(n25176) );
  INV_X1 U18554 ( .A(n20957), .ZN(n25177) );
  INV_X1 U18555 ( .A(n20957), .ZN(n25178) );
  INV_X1 U18556 ( .A(n20958), .ZN(n25179) );
  INV_X1 U18557 ( .A(n20958), .ZN(n25180) );
  INV_X1 U18558 ( .A(n20959), .ZN(n25181) );
  INV_X1 U18559 ( .A(n20959), .ZN(n25182) );
  INV_X1 U18560 ( .A(n20960), .ZN(n25183) );
  INV_X1 U18561 ( .A(n20961), .ZN(n25184) );
  INV_X1 U18562 ( .A(n20960), .ZN(n25185) );
  INV_X1 U18563 ( .A(n20962), .ZN(n25186) );
  INV_X1 U18564 ( .A(n20962), .ZN(n25187) );
  INV_X1 U18565 ( .A(n20964), .ZN(n25188) );
  INV_X1 U18566 ( .A(n20964), .ZN(n25189) );
  INV_X1 U18567 ( .A(n20966), .ZN(n25190) );
  INV_X1 U18568 ( .A(n20966), .ZN(n25191) );
  INV_X1 U18569 ( .A(n20967), .ZN(n25192) );
  INV_X1 U18570 ( .A(n20967), .ZN(n25193) );
  INV_X1 U18571 ( .A(n20968), .ZN(n25194) );
  INV_X1 U18572 ( .A(n20969), .ZN(n25195) );
  INV_X1 U18573 ( .A(n20969), .ZN(n25196) );
  INV_X1 U18574 ( .A(n20970), .ZN(n25197) );
  INV_X1 U18575 ( .A(n20972), .ZN(n25198) );
  INV_X1 U18576 ( .A(n20972), .ZN(n25199) );
  INV_X1 U18577 ( .A(n20973), .ZN(n25200) );
  INV_X1 U18578 ( .A(n20974), .ZN(n25201) );
  INV_X1 U18579 ( .A(n20974), .ZN(n25202) );
  INV_X1 U18580 ( .A(n20975), .ZN(n25203) );
  INV_X1 U18581 ( .A(n20977), .ZN(n25204) );
  INV_X1 U18582 ( .A(n20977), .ZN(n25205) );
  INV_X1 U18583 ( .A(n20978), .ZN(n25206) );
  INV_X1 U18584 ( .A(n27263), .ZN(n25207) );
  INV_X1 U18585 ( .A(n20980), .ZN(n25208) );
  INV_X1 U18586 ( .A(n20980), .ZN(n25209) );
  INV_X1 U18587 ( .A(n20981), .ZN(n25210) );
  INV_X1 U18588 ( .A(n20982), .ZN(n25211) );
  INV_X1 U18589 ( .A(n20982), .ZN(n25212) );
  INV_X1 U18590 ( .A(n20983), .ZN(n25213) );
  INV_X1 U18591 ( .A(n20984), .ZN(n25214) );
  INV_X1 U18592 ( .A(n20984), .ZN(n25215) );
  INV_X1 U18593 ( .A(n20985), .ZN(n25216) );
  INV_X1 U18594 ( .A(n20986), .ZN(n25217) );
  INV_X1 U18595 ( .A(n20986), .ZN(n25218) );
  INV_X1 U18596 ( .A(n27153), .ZN(n25219) );
  INV_X1 U18597 ( .A(n20988), .ZN(n25220) );
  INV_X1 U18598 ( .A(n20988), .ZN(n25221) );
  INV_X1 U18599 ( .A(n20989), .ZN(n25222) );
  INV_X1 U18600 ( .A(n20990), .ZN(n25223) );
  INV_X1 U18601 ( .A(n20990), .ZN(n25224) );
  INV_X1 U18602 ( .A(n20991), .ZN(n25225) );
  INV_X1 U18603 ( .A(n20991), .ZN(n25226) );
  INV_X1 U18604 ( .A(n20992), .ZN(n25227) );
  INV_X1 U18605 ( .A(n20992), .ZN(n25228) );
  INV_X1 U18606 ( .A(n20993), .ZN(n25229) );
  INV_X1 U18607 ( .A(n20993), .ZN(n25230) );
  INV_X1 U18608 ( .A(n20994), .ZN(n25231) );
  INV_X1 U18609 ( .A(n20994), .ZN(n25232) );
  INV_X1 U18610 ( .A(n20995), .ZN(n25233) );
  INV_X1 U18611 ( .A(n20995), .ZN(n25234) );
  INV_X1 U18612 ( .A(n20996), .ZN(n25235) );
  INV_X1 U18613 ( .A(n20996), .ZN(n25236) );
  INV_X1 U18614 ( .A(n20997), .ZN(n25237) );
  INV_X1 U18615 ( .A(n20997), .ZN(n25238) );
  INV_X1 U18616 ( .A(n20999), .ZN(n25239) );
  INV_X1 U18617 ( .A(n21002), .ZN(n25240) );
  INV_X1 U18618 ( .A(n21002), .ZN(n25241) );
  INV_X1 U18619 ( .A(n20619), .ZN(n25242) );
  INV_X1 U18620 ( .A(n25242), .ZN(n25243) );
  INV_X1 U18621 ( .A(n25242), .ZN(n25244) );
  INV_X1 U18622 ( .A(n21006), .ZN(n25245) );
  INV_X1 U18623 ( .A(n21006), .ZN(n25246) );
  INV_X1 U18624 ( .A(n21007), .ZN(n25247) );
  INV_X1 U18625 ( .A(n21007), .ZN(n25248) );
  INV_X1 U18626 ( .A(n21008), .ZN(n25249) );
  INV_X1 U18627 ( .A(n21008), .ZN(n25250) );
  INV_X1 U18628 ( .A(n24213), .ZN(n25251) );
  CLKBUF_X1 U18629 ( .A(n21424), .Z(n25252) );
  INV_X1 U18630 ( .A(n26747), .ZN(n25253) );
  INV_X1 U18631 ( .A(n25253), .ZN(n25254) );
  INV_X1 U18632 ( .A(n25253), .ZN(n25255) );
  INV_X1 U18633 ( .A(n24919), .ZN(n25256) );
  INV_X1 U18634 ( .A(n26745), .ZN(n25257) );
  INV_X1 U18635 ( .A(n25257), .ZN(n25258) );
  INV_X1 U18636 ( .A(n25257), .ZN(n25259) );
  CLKBUF_X1 U18637 ( .A(n24207), .Z(n26741) );
  INV_X1 U18638 ( .A(n26741), .ZN(n25260) );
  INV_X1 U18639 ( .A(n26741), .ZN(n25261) );
  INV_X1 U18640 ( .A(n26742), .ZN(n25262) );
  INV_X1 U18641 ( .A(n25262), .ZN(n25263) );
  INV_X1 U18642 ( .A(n25262), .ZN(n25264) );
  INV_X1 U18643 ( .A(n20722), .ZN(n25265) );
  INV_X1 U18644 ( .A(n19306), .ZN(n25266) );
  INV_X1 U18645 ( .A(n25266), .ZN(n25267) );
  INV_X1 U18646 ( .A(n25266), .ZN(n25268) );
  CLKBUF_X1 U18647 ( .A(n24201), .Z(n26734) );
  INV_X1 U18648 ( .A(n26734), .ZN(n25269) );
  INV_X1 U18649 ( .A(n26734), .ZN(n25270) );
  INV_X1 U18650 ( .A(n26735), .ZN(n25271) );
  INV_X1 U18651 ( .A(n25271), .ZN(n25272) );
  INV_X1 U18652 ( .A(n25271), .ZN(n25273) );
  CLKBUF_X1 U18653 ( .A(n26742), .Z(n25274) );
  INV_X1 U18654 ( .A(n19305), .ZN(n25275) );
  INV_X1 U18655 ( .A(n25275), .ZN(n25276) );
  INV_X1 U18656 ( .A(n25275), .ZN(n25277) );
  CLKBUF_X1 U18657 ( .A(n26735), .Z(n25278) );
  INV_X1 U18658 ( .A(n19304), .ZN(n25279) );
  INV_X1 U18659 ( .A(n25279), .ZN(n25280) );
  INV_X1 U18660 ( .A(n25279), .ZN(n25281) );
  INV_X1 U18661 ( .A(n21012), .ZN(n25282) );
  INV_X1 U18662 ( .A(n21012), .ZN(n25283) );
  INV_X1 U18663 ( .A(n24193), .ZN(n25284) );
  CLKBUF_X1 U18664 ( .A(n26943), .Z(n25285) );
  CLKBUF_X1 U18665 ( .A(n24185), .Z(n26725) );
  INV_X1 U18666 ( .A(n26725), .ZN(n25286) );
  INV_X1 U18667 ( .A(n26725), .ZN(n25287) );
  INV_X1 U18668 ( .A(n26950), .ZN(n25288) );
  INV_X1 U18669 ( .A(n21016), .ZN(n25289) );
  INV_X1 U18670 ( .A(n21016), .ZN(n25290) );
  INV_X1 U18671 ( .A(n21017), .ZN(n25291) );
  INV_X1 U18672 ( .A(n21017), .ZN(n25292) );
  CLKBUF_X1 U18673 ( .A(n24179), .Z(n26723) );
  INV_X1 U18674 ( .A(n26723), .ZN(n25293) );
  INV_X1 U18675 ( .A(n26723), .ZN(n25294) );
  INV_X1 U18676 ( .A(n19072), .ZN(n25295) );
  INV_X1 U18677 ( .A(n19072), .ZN(n25296) );
  INV_X1 U18678 ( .A(n21018), .ZN(n25297) );
  INV_X1 U18679 ( .A(n21018), .ZN(n25298) );
  INV_X1 U18680 ( .A(n21019), .ZN(n25299) );
  INV_X1 U18681 ( .A(n21019), .ZN(n25300) );
  CLKBUF_X1 U18682 ( .A(n24174), .Z(n26720) );
  INV_X1 U18683 ( .A(n26720), .ZN(n25301) );
  INV_X1 U18684 ( .A(n26720), .ZN(n25302) );
  INV_X1 U18685 ( .A(n19075), .ZN(n25303) );
  INV_X1 U18686 ( .A(n19075), .ZN(n25304) );
  INV_X1 U18687 ( .A(n21020), .ZN(n25305) );
  INV_X1 U18688 ( .A(n21020), .ZN(n25306) );
  INV_X1 U18689 ( .A(n21021), .ZN(n25307) );
  INV_X1 U18690 ( .A(n21021), .ZN(n25308) );
  INV_X1 U18691 ( .A(n24173), .ZN(n25309) );
  INV_X1 U18692 ( .A(n26717), .ZN(n25310) );
  INV_X1 U18693 ( .A(n25310), .ZN(n25311) );
  INV_X1 U18694 ( .A(n21025), .ZN(n25312) );
  INV_X1 U18695 ( .A(n21025), .ZN(n25313) );
  INV_X1 U18696 ( .A(n18149), .ZN(n25314) );
  INV_X1 U18697 ( .A(n18149), .ZN(n25315) );
  INV_X1 U18698 ( .A(n21026), .ZN(n25316) );
  INV_X1 U18699 ( .A(n21026), .ZN(n25317) );
  INV_X1 U18700 ( .A(n21027), .ZN(n25318) );
  INV_X1 U18701 ( .A(n21027), .ZN(n25319) );
  INV_X1 U18702 ( .A(n21028), .ZN(n25320) );
  INV_X1 U18703 ( .A(n21028), .ZN(n25321) );
  INV_X1 U18704 ( .A(n21030), .ZN(n25322) );
  INV_X1 U18705 ( .A(n21030), .ZN(n25323) );
  INV_X1 U18706 ( .A(n21032), .ZN(n25324) );
  INV_X1 U18707 ( .A(n21032), .ZN(n25325) );
  INV_X1 U18708 ( .A(n21033), .ZN(n25326) );
  INV_X1 U18709 ( .A(n21033), .ZN(n25327) );
  INV_X1 U18710 ( .A(n21035), .ZN(n25328) );
  INV_X1 U18711 ( .A(n21035), .ZN(n25329) );
  INV_X1 U18712 ( .A(n21037), .ZN(n25330) );
  INV_X1 U18713 ( .A(n21037), .ZN(n25331) );
  INV_X1 U18714 ( .A(n26690), .ZN(n25332) );
  INV_X1 U18715 ( .A(n21039), .ZN(n25333) );
  INV_X1 U18716 ( .A(n21039), .ZN(n25334) );
  INV_X1 U18717 ( .A(n21040), .ZN(n25335) );
  INV_X1 U18718 ( .A(n21040), .ZN(n25336) );
  INV_X1 U18719 ( .A(n26688), .ZN(n25337) );
  INV_X1 U18720 ( .A(n21042), .ZN(n25338) );
  INV_X1 U18721 ( .A(n21042), .ZN(n25339) );
  INV_X1 U18722 ( .A(n26689), .ZN(n25340) );
  INV_X1 U18723 ( .A(n21044), .ZN(n25341) );
  INV_X1 U18724 ( .A(n21044), .ZN(n25342) );
  INV_X1 U18725 ( .A(n26675), .ZN(n25343) );
  INV_X1 U18726 ( .A(n21046), .ZN(n25344) );
  INV_X1 U18727 ( .A(n21046), .ZN(n25345) );
  INV_X1 U18728 ( .A(n21048), .ZN(n25346) );
  INV_X1 U18729 ( .A(n21048), .ZN(n25347) );
  INV_X1 U18730 ( .A(n21049), .ZN(n25348) );
  INV_X1 U18731 ( .A(n21049), .ZN(n25349) );
  INV_X1 U18732 ( .A(n21050), .ZN(n25350) );
  INV_X1 U18733 ( .A(n21050), .ZN(n25351) );
  INV_X1 U18734 ( .A(n21051), .ZN(n25352) );
  INV_X1 U18735 ( .A(n21051), .ZN(n25353) );
  INV_X1 U18736 ( .A(n21052), .ZN(n25354) );
  INV_X1 U18737 ( .A(n21052), .ZN(n25355) );
  INV_X1 U18738 ( .A(n21053), .ZN(n25356) );
  INV_X1 U18739 ( .A(n21053), .ZN(n25357) );
  INV_X1 U18740 ( .A(n21054), .ZN(n25358) );
  INV_X1 U18741 ( .A(n21054), .ZN(n25359) );
  INV_X1 U18742 ( .A(n21055), .ZN(n25360) );
  INV_X1 U18743 ( .A(n21055), .ZN(n25361) );
  INV_X1 U18744 ( .A(n21056), .ZN(n25362) );
  INV_X1 U18745 ( .A(n21057), .ZN(n25363) );
  INV_X1 U18746 ( .A(n21060), .ZN(n25364) );
  INV_X1 U18747 ( .A(n21060), .ZN(n25365) );
  INV_X1 U18748 ( .A(n21061), .ZN(n25366) );
  INV_X1 U18749 ( .A(n21064), .ZN(n25367) );
  INV_X1 U18750 ( .A(n21067), .ZN(n25368) );
  INV_X1 U18751 ( .A(n21067), .ZN(n25369) );
  INV_X1 U18752 ( .A(n21068), .ZN(n25370) );
  INV_X1 U18753 ( .A(n21068), .ZN(n25371) );
  INV_X1 U18754 ( .A(n21069), .ZN(n25372) );
  INV_X1 U18755 ( .A(n21069), .ZN(n25373) );
  INV_X1 U18756 ( .A(n21070), .ZN(n25374) );
  INV_X1 U18757 ( .A(n21070), .ZN(n25375) );
  INV_X1 U18758 ( .A(n4571), .ZN(n25376) );
  INV_X1 U18759 ( .A(n25376), .ZN(n25377) );
  INV_X1 U18760 ( .A(n25376), .ZN(n25378) );
  INV_X1 U18761 ( .A(n21071), .ZN(n25379) );
  INV_X1 U18762 ( .A(n21071), .ZN(n25380) );
  INV_X1 U18763 ( .A(n21072), .ZN(n25381) );
  INV_X1 U18764 ( .A(n21072), .ZN(n25382) );
  INV_X1 U18765 ( .A(n21073), .ZN(n25383) );
  INV_X1 U18766 ( .A(n21073), .ZN(n25384) );
  INV_X1 U18767 ( .A(n21074), .ZN(n25385) );
  INV_X1 U18768 ( .A(n21074), .ZN(n25386) );
  INV_X1 U18769 ( .A(n21075), .ZN(n25387) );
  INV_X1 U18770 ( .A(n21075), .ZN(n25388) );
  INV_X1 U18771 ( .A(n21076), .ZN(n25389) );
  INV_X1 U18772 ( .A(n21076), .ZN(n25390) );
  INV_X1 U18773 ( .A(n21077), .ZN(n25391) );
  INV_X1 U18774 ( .A(n21077), .ZN(n25392) );
  INV_X1 U18775 ( .A(n21078), .ZN(n25393) );
  INV_X1 U18776 ( .A(n21078), .ZN(n25394) );
  INV_X1 U18777 ( .A(n21079), .ZN(n25395) );
  INV_X1 U18778 ( .A(n21079), .ZN(n25396) );
  INV_X1 U18779 ( .A(n21080), .ZN(n25397) );
  INV_X1 U18780 ( .A(n21080), .ZN(n25398) );
  INV_X1 U18781 ( .A(n21081), .ZN(n25399) );
  INV_X1 U18782 ( .A(n21081), .ZN(n25400) );
  INV_X1 U18783 ( .A(n21082), .ZN(n25401) );
  INV_X1 U18784 ( .A(n21082), .ZN(n25402) );
  INV_X1 U18785 ( .A(n21083), .ZN(n25403) );
  INV_X1 U18786 ( .A(n21083), .ZN(n25404) );
  INV_X1 U18787 ( .A(n21084), .ZN(n25405) );
  INV_X1 U18788 ( .A(n21084), .ZN(n25406) );
  INV_X1 U18789 ( .A(n21085), .ZN(n25407) );
  INV_X1 U18790 ( .A(n21085), .ZN(n25408) );
  INV_X1 U18791 ( .A(n21086), .ZN(n25409) );
  INV_X1 U18792 ( .A(n21086), .ZN(n25410) );
  INV_X1 U18793 ( .A(n21087), .ZN(n25411) );
  INV_X1 U18794 ( .A(n21087), .ZN(n25412) );
  INV_X1 U18795 ( .A(n21088), .ZN(n25413) );
  INV_X1 U18796 ( .A(n21088), .ZN(n25414) );
  INV_X1 U18797 ( .A(n21089), .ZN(n25415) );
  INV_X1 U18798 ( .A(n21089), .ZN(n25416) );
  INV_X1 U18799 ( .A(n21090), .ZN(n25417) );
  INV_X1 U18800 ( .A(n21090), .ZN(n25418) );
  INV_X1 U18801 ( .A(n21091), .ZN(n25419) );
  INV_X1 U18802 ( .A(n21091), .ZN(n25420) );
  INV_X1 U18803 ( .A(n21092), .ZN(n25421) );
  INV_X1 U18804 ( .A(n21092), .ZN(n25422) );
  INV_X1 U18805 ( .A(n21093), .ZN(n25423) );
  INV_X1 U18806 ( .A(n21093), .ZN(n25424) );
  INV_X1 U18807 ( .A(n21094), .ZN(n25425) );
  INV_X1 U18808 ( .A(n21094), .ZN(n25426) );
  INV_X1 U18809 ( .A(n21095), .ZN(n25427) );
  INV_X1 U18810 ( .A(n21095), .ZN(n25428) );
  INV_X1 U18811 ( .A(n21096), .ZN(n25429) );
  INV_X1 U18812 ( .A(n21096), .ZN(n25430) );
  INV_X1 U18813 ( .A(n21097), .ZN(n25431) );
  INV_X1 U18814 ( .A(n21097), .ZN(n25432) );
  INV_X1 U18815 ( .A(n21098), .ZN(n25433) );
  INV_X1 U18816 ( .A(n21098), .ZN(n25434) );
  INV_X1 U18817 ( .A(n21099), .ZN(n25435) );
  INV_X1 U18818 ( .A(n21099), .ZN(n25436) );
  INV_X1 U18819 ( .A(n21100), .ZN(n25437) );
  INV_X1 U18820 ( .A(n21100), .ZN(n25438) );
  INV_X1 U18821 ( .A(n21101), .ZN(n25439) );
  INV_X1 U18822 ( .A(n21101), .ZN(n25440) );
  INV_X1 U18823 ( .A(n21102), .ZN(n25441) );
  INV_X1 U18824 ( .A(n21102), .ZN(n25442) );
  INV_X1 U18825 ( .A(n21103), .ZN(n25443) );
  INV_X1 U18826 ( .A(n21103), .ZN(n25444) );
  INV_X1 U18827 ( .A(n21104), .ZN(n25445) );
  INV_X1 U18828 ( .A(n21104), .ZN(n25446) );
  INV_X1 U18829 ( .A(n21105), .ZN(n25447) );
  INV_X1 U18830 ( .A(n21105), .ZN(n25448) );
  INV_X1 U18831 ( .A(n21106), .ZN(n25449) );
  INV_X1 U18832 ( .A(n21106), .ZN(n25450) );
  INV_X1 U18833 ( .A(n21107), .ZN(n25451) );
  INV_X1 U18834 ( .A(n21107), .ZN(n25452) );
  INV_X1 U18835 ( .A(n21108), .ZN(n25453) );
  INV_X1 U18836 ( .A(n21108), .ZN(n25454) );
  INV_X1 U18837 ( .A(n21109), .ZN(n25455) );
  INV_X1 U18838 ( .A(n21109), .ZN(n25456) );
  INV_X1 U18839 ( .A(n21110), .ZN(n25457) );
  INV_X1 U18840 ( .A(n21110), .ZN(n25458) );
  INV_X1 U18841 ( .A(n21111), .ZN(n25459) );
  INV_X1 U18842 ( .A(n21111), .ZN(n25460) );
  INV_X1 U18843 ( .A(n21112), .ZN(n25461) );
  INV_X1 U18844 ( .A(n21112), .ZN(n25462) );
  INV_X1 U18845 ( .A(n21113), .ZN(n25463) );
  INV_X1 U18846 ( .A(n21113), .ZN(n25464) );
  INV_X1 U18847 ( .A(n40530), .ZN(n25465) );
  INV_X1 U18848 ( .A(n25465), .ZN(n25466) );
  INV_X1 U18849 ( .A(n25465), .ZN(n25467) );
  INV_X1 U18850 ( .A(n21114), .ZN(n25468) );
  INV_X1 U18851 ( .A(n21114), .ZN(n25469) );
  INV_X1 U18852 ( .A(n21115), .ZN(n25470) );
  INV_X1 U18853 ( .A(n21115), .ZN(n25471) );
  INV_X1 U18854 ( .A(n21116), .ZN(n25472) );
  INV_X1 U18855 ( .A(n21116), .ZN(n25473) );
  INV_X1 U18856 ( .A(n21117), .ZN(n25474) );
  INV_X1 U18857 ( .A(n21117), .ZN(n25475) );
  INV_X1 U18858 ( .A(n21118), .ZN(n25476) );
  INV_X1 U18859 ( .A(n21118), .ZN(n25477) );
  INV_X1 U18860 ( .A(n21119), .ZN(n25478) );
  INV_X1 U18861 ( .A(n21119), .ZN(n25479) );
  INV_X1 U18862 ( .A(n21120), .ZN(n25480) );
  INV_X1 U18863 ( .A(n21120), .ZN(n25481) );
  INV_X1 U18864 ( .A(n21121), .ZN(n25482) );
  INV_X1 U18865 ( .A(n21121), .ZN(n25483) );
  INV_X1 U18866 ( .A(n21122), .ZN(n25484) );
  INV_X1 U18867 ( .A(n21122), .ZN(n25485) );
  INV_X1 U18868 ( .A(n21123), .ZN(n25486) );
  INV_X1 U18869 ( .A(n21123), .ZN(n25487) );
  INV_X1 U18870 ( .A(n21124), .ZN(n25488) );
  INV_X1 U18871 ( .A(n21124), .ZN(n25489) );
  INV_X1 U18872 ( .A(n21125), .ZN(n25490) );
  INV_X1 U18873 ( .A(n21125), .ZN(n25491) );
  INV_X1 U18874 ( .A(n21126), .ZN(n25492) );
  INV_X1 U18875 ( .A(n21126), .ZN(n25493) );
  INV_X1 U18876 ( .A(n21127), .ZN(n25494) );
  INV_X1 U18877 ( .A(n21127), .ZN(n25495) );
  INV_X1 U18878 ( .A(n21128), .ZN(n25496) );
  INV_X1 U18879 ( .A(n21128), .ZN(n25497) );
  INV_X1 U18880 ( .A(n21129), .ZN(n25498) );
  INV_X1 U18881 ( .A(n21129), .ZN(n25499) );
  INV_X1 U18882 ( .A(n21130), .ZN(n25500) );
  INV_X1 U18883 ( .A(n21130), .ZN(n25501) );
  INV_X1 U18884 ( .A(n21131), .ZN(n25502) );
  INV_X1 U18885 ( .A(n21131), .ZN(n25503) );
  INV_X1 U18886 ( .A(n21132), .ZN(n25504) );
  INV_X1 U18887 ( .A(n21132), .ZN(n25505) );
  INV_X1 U18888 ( .A(n21133), .ZN(n25506) );
  INV_X1 U18889 ( .A(n21133), .ZN(n25507) );
  INV_X1 U18890 ( .A(n21134), .ZN(n25508) );
  INV_X1 U18891 ( .A(n21134), .ZN(n25509) );
  INV_X1 U18892 ( .A(n4029), .ZN(n25510) );
  INV_X1 U18893 ( .A(n21136), .ZN(n25511) );
  INV_X1 U18894 ( .A(n21136), .ZN(n25512) );
  INV_X1 U18895 ( .A(n21137), .ZN(n25513) );
  INV_X1 U18896 ( .A(n21137), .ZN(n25514) );
  INV_X1 U18897 ( .A(n25649), .ZN(n25515) );
  INV_X1 U18898 ( .A(n21139), .ZN(n25516) );
  INV_X1 U18899 ( .A(n21143), .ZN(n25517) );
  INV_X1 U18900 ( .A(n21143), .ZN(n25518) );
  INV_X1 U18901 ( .A(n25648), .ZN(n25519) );
  INV_X1 U18902 ( .A(n21145), .ZN(n25520) );
  INV_X1 U18903 ( .A(n21146), .ZN(n25521) );
  INV_X1 U18904 ( .A(n21149), .ZN(n25522) );
  INV_X1 U18905 ( .A(n21152), .ZN(n25523) );
  INV_X1 U18906 ( .A(n26999), .ZN(n27000) );
  INV_X1 U18907 ( .A(n27000), .ZN(n25524) );
  INV_X1 U18908 ( .A(n27000), .ZN(n25525) );
  INV_X1 U18909 ( .A(n21155), .ZN(n25526) );
  INV_X1 U18910 ( .A(n21158), .ZN(n25527) );
  INV_X1 U18911 ( .A(n27246), .ZN(n25528) );
  INV_X1 U18912 ( .A(n21162), .ZN(n25529) );
  INV_X1 U18913 ( .A(n21163), .ZN(n25530) );
  INV_X1 U18914 ( .A(n21166), .ZN(n25531) );
  INV_X1 U18915 ( .A(n21169), .ZN(n25532) );
  INV_X1 U18916 ( .A(n21170), .ZN(n25533) );
  INV_X1 U18917 ( .A(n21163), .ZN(n25534) );
  INV_X1 U18918 ( .A(n25337), .ZN(n25535) );
  INV_X1 U18919 ( .A(n21177), .ZN(n25536) );
  INV_X1 U18920 ( .A(n21170), .ZN(n25537) );
  INV_X1 U18921 ( .A(n25332), .ZN(n25538) );
  INV_X1 U18922 ( .A(n21184), .ZN(n25539) );
  INV_X1 U18923 ( .A(n17992), .ZN(n25540) );
  INV_X1 U18924 ( .A(n21188), .ZN(n25541) );
  INV_X1 U18925 ( .A(n21191), .ZN(n25542) );
  CLKBUF_X1 U18926 ( .A(n24626), .Z(n27251) );
  INV_X1 U18927 ( .A(n27251), .ZN(n25543) );
  INV_X1 U18928 ( .A(n27251), .ZN(n25544) );
  INV_X1 U18929 ( .A(n21194), .ZN(n25545) );
  INV_X1 U18930 ( .A(n21197), .ZN(n25546) );
  INV_X1 U18931 ( .A(n24620), .ZN(n25547) );
  INV_X1 U18932 ( .A(n24629), .ZN(n25548) );
  CLKBUF_X1 U18933 ( .A(n24618), .Z(n27243) );
  INV_X1 U18934 ( .A(n27243), .ZN(n25549) );
  INV_X1 U18935 ( .A(n27243), .ZN(n25550) );
  CLKBUF_X1 U18936 ( .A(n24616), .Z(n27187) );
  INV_X1 U18937 ( .A(n27187), .ZN(n25551) );
  INV_X1 U18938 ( .A(n27187), .ZN(n25552) );
  INV_X1 U18939 ( .A(n19189), .ZN(n25553) );
  INV_X1 U18940 ( .A(n19189), .ZN(n25554) );
  INV_X1 U18941 ( .A(n21200), .ZN(n25555) );
  CLKBUF_X1 U18942 ( .A(n24611), .Z(n27163) );
  INV_X1 U18943 ( .A(n27163), .ZN(n25556) );
  INV_X1 U18944 ( .A(n27163), .ZN(n25557) );
  INV_X1 U18945 ( .A(n21203), .ZN(n25558) );
  INV_X1 U18946 ( .A(n21206), .ZN(n25559) );
  INV_X1 U18947 ( .A(n21210), .ZN(n25560) );
  INV_X1 U18948 ( .A(n24605), .ZN(n25561) );
  INV_X1 U18949 ( .A(n24614), .ZN(n25562) );
  INV_X1 U18950 ( .A(n21214), .ZN(n25563) );
  INV_X1 U18951 ( .A(n21217), .ZN(n25564) );
  INV_X1 U18952 ( .A(n21220), .ZN(n25565) );
  INV_X1 U18953 ( .A(n21223), .ZN(n25566) );
  INV_X1 U18954 ( .A(n21226), .ZN(n25567) );
  INV_X1 U18955 ( .A(n21229), .ZN(n25568) );
  INV_X1 U18956 ( .A(n27047), .ZN(n25569) );
  INV_X1 U18957 ( .A(n21235), .ZN(n25570) );
  INV_X1 U18958 ( .A(n21238), .ZN(n25571) );
  INV_X1 U18959 ( .A(n17990), .ZN(n25572) );
  INV_X1 U18960 ( .A(n21242), .ZN(n25573) );
  INV_X1 U18961 ( .A(n21245), .ZN(n25574) );
  INV_X1 U18962 ( .A(n21248), .ZN(n25575) );
  CLKBUF_X1 U18963 ( .A(n20543), .Z(n27223) );
  INV_X1 U18964 ( .A(n27223), .ZN(n25576) );
  INV_X1 U18965 ( .A(n22892), .ZN(n25577) );
  INV_X1 U18966 ( .A(n25577), .ZN(n25578) );
  INV_X1 U18967 ( .A(n25577), .ZN(n25579) );
  INV_X1 U18968 ( .A(n21252), .ZN(n25580) );
  CLKBUF_X1 U18969 ( .A(n20542), .Z(n27224) );
  INV_X1 U18970 ( .A(n27224), .ZN(n25581) );
  INV_X1 U18971 ( .A(n21257), .ZN(n25582) );
  INV_X1 U18972 ( .A(n21260), .ZN(n25583) );
  INV_X1 U18973 ( .A(n21263), .ZN(n25584) );
  INV_X1 U18974 ( .A(n21266), .ZN(n25585) );
  CLKBUF_X1 U18975 ( .A(n24484), .Z(n27200) );
  INV_X1 U18976 ( .A(n27200), .ZN(n25586) );
  INV_X1 U18977 ( .A(n22887), .ZN(n25587) );
  INV_X1 U18978 ( .A(n25587), .ZN(n25588) );
  INV_X1 U18979 ( .A(n25587), .ZN(n25589) );
  CLKBUF_X1 U18980 ( .A(n24760), .Z(n27202) );
  INV_X1 U18981 ( .A(n27202), .ZN(n255901) );
  INV_X1 U18982 ( .A(n19313), .ZN(n25591) );
  INV_X1 U18983 ( .A(n25591), .ZN(n25592) );
  INV_X1 U18984 ( .A(n25591), .ZN(n25593) );
  INV_X1 U18985 ( .A(n21272), .ZN(n25594) );
  INV_X1 U18986 ( .A(n21275), .ZN(n25595) );
  CLKBUF_X1 U18987 ( .A(n22824), .Z(n26752) );
  INV_X1 U18988 ( .A(n26752), .ZN(n25596) );
  INV_X1 U18989 ( .A(n26752), .ZN(n25597) );
  INV_X1 U18990 ( .A(n24226), .ZN(n25598) );
  INV_X1 U18991 ( .A(n25598), .ZN(n25599) );
  INV_X1 U18992 ( .A(n25598), .ZN(n256001) );
  CLKBUF_X1 U18993 ( .A(n22821), .Z(n26749) );
  INV_X1 U18994 ( .A(n26749), .ZN(n25601) );
  INV_X1 U18995 ( .A(n26749), .ZN(n25602) );
  INV_X1 U18996 ( .A(n24222), .ZN(n25603) );
  INV_X1 U18997 ( .A(n25603), .ZN(n25604) );
  INV_X1 U18998 ( .A(n25603), .ZN(n25605) );
  INV_X1 U18999 ( .A(n21278), .ZN(n25606) );
  INV_X1 U19000 ( .A(n26976), .ZN(n25607) );
  INV_X1 U19001 ( .A(n24832), .ZN(n25608) );
  INV_X1 U19002 ( .A(n22817), .ZN(n25609) );
  INV_X1 U19003 ( .A(n25609), .ZN(n256101) );
  INV_X1 U19004 ( .A(n21281), .ZN(n25611) );
  INV_X1 U19005 ( .A(n21281), .ZN(n25612) );
  INV_X1 U19006 ( .A(n26746), .ZN(n25613) );
  INV_X1 U19007 ( .A(n25613), .ZN(n25614) );
  INV_X1 U19008 ( .A(n25613), .ZN(n25615) );
  INV_X1 U19009 ( .A(n21285), .ZN(n25616) );
  INV_X1 U19010 ( .A(n25883), .ZN(n25617) );
  INV_X1 U19011 ( .A(n21289), .ZN(n25618) );
  INV_X1 U19012 ( .A(n21292), .ZN(n25619) );
  INV_X1 U19013 ( .A(n21295), .ZN(n256201) );
  INV_X1 U19014 ( .A(n21298), .ZN(n25621) );
  INV_X1 U19015 ( .A(n21301), .ZN(n25622) );
  INV_X1 U19016 ( .A(n21304), .ZN(n25623) );
  INV_X1 U19017 ( .A(n21307), .ZN(n25624) );
  INV_X1 U19018 ( .A(n21310), .ZN(n25625) );
  INV_X1 U19019 ( .A(n21313), .ZN(n25626) );
  INV_X1 U19020 ( .A(n21316), .ZN(n25627) );
  INV_X1 U19021 ( .A(n21319), .ZN(n25628) );
  INV_X1 U19022 ( .A(n21322), .ZN(n25629) );
  INV_X1 U19023 ( .A(n25528), .ZN(n256301) );
  INV_X1 U19024 ( .A(n21329), .ZN(n25631) );
  INV_X1 U19025 ( .A(n21332), .ZN(n25632) );
  INV_X1 U19026 ( .A(n21335), .ZN(n25633) );
  INV_X1 U19027 ( .A(n21335), .ZN(n25634) );
  INV_X1 U19028 ( .A(n21339), .ZN(n25635) );
  INV_X1 U19029 ( .A(n21343), .ZN(n25636) );
  INV_X1 U19030 ( .A(n21346), .ZN(n25637) );
  INV_X1 U19031 ( .A(n21349), .ZN(n25638) );
  INV_X1 U19032 ( .A(n5205), .ZN(n25639) );
  INV_X1 U19033 ( .A(n21353), .ZN(n256401) );
  INV_X1 U19034 ( .A(n21357), .ZN(n25641) );
  INV_X1 U19035 ( .A(n21360), .ZN(n25642) );
  INV_X1 U19036 ( .A(n21364), .ZN(n25643) );
  INV_X1 U19037 ( .A(n5133), .ZN(n25644) );
  INV_X1 U19038 ( .A(n21374), .ZN(n25645) );
  INV_X1 U19039 ( .A(n21374), .ZN(n25646) );
  INV_X1 U19040 ( .A(n4721), .ZN(n25647) );
  INV_X1 U19041 ( .A(n25647), .ZN(n25648) );
  INV_X1 U19042 ( .A(n25647), .ZN(n25649) );
  INV_X1 U19043 ( .A(n21376), .ZN(n256501) );
  INV_X1 U19044 ( .A(n27043), .ZN(n25651) );
  INV_X1 U19045 ( .A(n21380), .ZN(n25652) );
  INV_X1 U19046 ( .A(n17132), .ZN(n25653) );
  INV_X1 U19047 ( .A(n21384), .ZN(n25654) );
  INV_X1 U19048 ( .A(n21388), .ZN(n25655) );
  INV_X1 U19049 ( .A(n21388), .ZN(n25656) );
  INV_X1 U19050 ( .A(n21391), .ZN(n25657) );
  INV_X1 U19051 ( .A(n21394), .ZN(n25658) );
  INV_X1 U19052 ( .A(n18277), .ZN(n25659) );
  INV_X1 U19053 ( .A(n21399), .ZN(n256601) );
  INV_X1 U19054 ( .A(n21400), .ZN(n25661) );
  INV_X1 U19055 ( .A(n22973), .ZN(n25662) );
  INV_X1 U19056 ( .A(n22974), .ZN(n25663) );
  INV_X1 U19057 ( .A(n22973), .ZN(n25664) );
  INV_X1 U19058 ( .A(n22974), .ZN(n25665) );
  INV_X1 U19059 ( .A(n22976), .ZN(n25666) );
  INV_X1 U19060 ( .A(n22975), .ZN(n25667) );
  INV_X1 U19061 ( .A(n22976), .ZN(n25668) );
  INV_X1 U19062 ( .A(n22975), .ZN(n25669) );
  INV_X1 U19063 ( .A(n22978), .ZN(n256701) );
  INV_X1 U19064 ( .A(n22977), .ZN(n25671) );
  INV_X1 U19065 ( .A(n22978), .ZN(n25672) );
  INV_X1 U19066 ( .A(n22977), .ZN(n25673) );
  INV_X1 U19067 ( .A(n21404), .ZN(n25674) );
  INV_X1 U19068 ( .A(n21404), .ZN(n25675) );
  INV_X1 U19069 ( .A(n21405), .ZN(n25676) );
  INV_X1 U19070 ( .A(n21405), .ZN(n25677) );
  INV_X1 U19071 ( .A(n22980), .ZN(n25678) );
  INV_X1 U19072 ( .A(n22979), .ZN(n25679) );
  INV_X1 U19073 ( .A(n22980), .ZN(n256801) );
  INV_X1 U19074 ( .A(n22979), .ZN(n25681) );
  INV_X1 U19075 ( .A(n25955), .ZN(n25682) );
  INV_X1 U19076 ( .A(n22983), .ZN(n25683) );
  INV_X1 U19077 ( .A(n22982), .ZN(n25684) );
  INV_X1 U19078 ( .A(n22983), .ZN(n25685) );
  INV_X1 U19079 ( .A(n22982), .ZN(n25686) );
  INV_X1 U19080 ( .A(n22985), .ZN(n25687) );
  INV_X1 U19081 ( .A(n22984), .ZN(n25688) );
  INV_X1 U19082 ( .A(n22985), .ZN(n25689) );
  INV_X1 U19083 ( .A(n22984), .ZN(n256901) );
  INV_X1 U19084 ( .A(n22987), .ZN(n25691) );
  INV_X1 U19085 ( .A(n22986), .ZN(n25692) );
  INV_X1 U19086 ( .A(n22987), .ZN(n25693) );
  INV_X1 U19087 ( .A(n22986), .ZN(n25694) );
  INV_X1 U19088 ( .A(n25947), .ZN(n25695) );
  INV_X1 U19089 ( .A(n22990), .ZN(n25696) );
  INV_X1 U19090 ( .A(n22989), .ZN(n25697) );
  INV_X1 U19091 ( .A(n22990), .ZN(n25698) );
  INV_X1 U19092 ( .A(n22989), .ZN(n25699) );
  INV_X1 U19093 ( .A(n22993), .ZN(n257001) );
  INV_X1 U19094 ( .A(n22992), .ZN(n25701) );
  INV_X1 U19095 ( .A(n22993), .ZN(n25702) );
  INV_X1 U19096 ( .A(n22992), .ZN(n25703) );
  INV_X1 U19097 ( .A(n22995), .ZN(n25704) );
  INV_X1 U19098 ( .A(n22994), .ZN(n25705) );
  INV_X1 U19099 ( .A(n22995), .ZN(n25706) );
  INV_X1 U19100 ( .A(n22994), .ZN(n25707) );
  INV_X1 U19101 ( .A(n22997), .ZN(n25708) );
  INV_X1 U19102 ( .A(n22996), .ZN(n25709) );
  INV_X1 U19103 ( .A(n22997), .ZN(n257101) );
  INV_X1 U19104 ( .A(n22996), .ZN(n25711) );
  INV_X1 U19105 ( .A(n23000), .ZN(n25712) );
  INV_X1 U19106 ( .A(n22999), .ZN(n25713) );
  INV_X1 U19107 ( .A(n23000), .ZN(n25714) );
  INV_X1 U19108 ( .A(n22999), .ZN(n25715) );
  INV_X1 U19109 ( .A(n23002), .ZN(n25716) );
  INV_X1 U19110 ( .A(n23001), .ZN(n25717) );
  INV_X1 U19111 ( .A(n23002), .ZN(n25718) );
  INV_X1 U19112 ( .A(n23001), .ZN(n25719) );
  INV_X1 U19113 ( .A(n23003), .ZN(n257201) );
  INV_X1 U19114 ( .A(n23004), .ZN(n25721) );
  INV_X1 U19115 ( .A(n23003), .ZN(n25722) );
  INV_X1 U19116 ( .A(n23004), .ZN(n25723) );
  INV_X1 U19117 ( .A(n23005), .ZN(n25724) );
  INV_X1 U19118 ( .A(n23006), .ZN(n25725) );
  INV_X1 U19119 ( .A(n23005), .ZN(n25726) );
  INV_X1 U19120 ( .A(n23006), .ZN(n25727) );
  INV_X1 U19121 ( .A(n23007), .ZN(n25728) );
  INV_X1 U19122 ( .A(n23008), .ZN(n25729) );
  INV_X1 U19123 ( .A(n23007), .ZN(n257301) );
  INV_X1 U19124 ( .A(n23008), .ZN(n25731) );
  INV_X1 U19125 ( .A(n23009), .ZN(n25732) );
  INV_X1 U19126 ( .A(n23010), .ZN(n25733) );
  INV_X1 U19127 ( .A(n23009), .ZN(n25734) );
  INV_X1 U19128 ( .A(n23010), .ZN(n25735) );
  INV_X1 U19129 ( .A(n23013), .ZN(n25736) );
  INV_X1 U19130 ( .A(n23012), .ZN(n25737) );
  INV_X1 U19131 ( .A(n23013), .ZN(n25738) );
  INV_X1 U19132 ( .A(n21409), .ZN(n25739) );
  INV_X1 U19133 ( .A(n21410), .ZN(n257401) );
  INV_X1 U19134 ( .A(n21409), .ZN(n25741) );
  INV_X1 U19135 ( .A(n23015), .ZN(n25742) );
  INV_X1 U19136 ( .A(n23015), .ZN(n25743) );
  INV_X1 U19137 ( .A(n21414), .ZN(n25744) );
  INV_X1 U19138 ( .A(n21414), .ZN(n25745) );
  INV_X1 U19139 ( .A(n23016), .ZN(n25746) );
  INV_X1 U19140 ( .A(n23017), .ZN(n25747) );
  INV_X1 U19141 ( .A(n23016), .ZN(n25748) );
  INV_X1 U19142 ( .A(n23017), .ZN(n25749) );
  INV_X1 U19143 ( .A(n23019), .ZN(n25750) );
  INV_X1 U19144 ( .A(n23018), .ZN(n25751) );
  INV_X1 U19145 ( .A(n23019), .ZN(n25752) );
  INV_X1 U19146 ( .A(n23018), .ZN(n25753) );
  INV_X1 U19147 ( .A(n23020), .ZN(n25754) );
  INV_X1 U19148 ( .A(n23021), .ZN(n25755) );
  INV_X1 U19149 ( .A(n23020), .ZN(n25756) );
  INV_X1 U19150 ( .A(n23021), .ZN(n25757) );
  INV_X1 U19151 ( .A(n23022), .ZN(n25758) );
  INV_X1 U19152 ( .A(n23023), .ZN(n25759) );
  INV_X1 U19153 ( .A(n23022), .ZN(n25760) );
  INV_X1 U19154 ( .A(n23023), .ZN(n25761) );
  INV_X1 U19155 ( .A(n25090), .ZN(n25762) );
  INV_X1 U19156 ( .A(n19020), .ZN(n25763) );
  INV_X1 U19157 ( .A(n27236), .ZN(n25764) );
  INV_X1 U19158 ( .A(n25764), .ZN(n25765) );
  INV_X1 U19159 ( .A(n25764), .ZN(n25766) );
  INV_X1 U19160 ( .A(n23025), .ZN(n25767) );
  INV_X1 U19161 ( .A(n23024), .ZN(n25768) );
  INV_X1 U19162 ( .A(n23025), .ZN(n25769) );
  INV_X1 U19163 ( .A(n23024), .ZN(n25770) );
  INV_X1 U19164 ( .A(n23027), .ZN(n25771) );
  INV_X1 U19165 ( .A(n23026), .ZN(n25772) );
  INV_X1 U19166 ( .A(n23026), .ZN(n25773) );
  INV_X1 U19167 ( .A(n23027), .ZN(n25774) );
  INV_X1 U19168 ( .A(n23029), .ZN(n25775) );
  INV_X1 U19169 ( .A(n23028), .ZN(n25776) );
  INV_X1 U19170 ( .A(n23028), .ZN(n25777) );
  INV_X1 U19171 ( .A(n23029), .ZN(n25778) );
  INV_X1 U19172 ( .A(n23031), .ZN(n25779) );
  INV_X1 U19173 ( .A(n23030), .ZN(n25780) );
  INV_X1 U19174 ( .A(n23031), .ZN(n25781) );
  INV_X1 U19175 ( .A(n23030), .ZN(n25782) );
  INV_X1 U19176 ( .A(n19023), .ZN(n25783) );
  INV_X1 U19177 ( .A(n25097), .ZN(n25784) );
  INV_X1 U19178 ( .A(n27240), .ZN(n25785) );
  INV_X1 U19179 ( .A(n25785), .ZN(n25786) );
  INV_X1 U19180 ( .A(n25785), .ZN(n25787) );
  INV_X1 U19181 ( .A(n23033), .ZN(n25788) );
  INV_X1 U19182 ( .A(n23032), .ZN(n25789) );
  INV_X1 U19183 ( .A(n23032), .ZN(n25790) );
  INV_X1 U19184 ( .A(n23033), .ZN(n25791) );
  INV_X1 U19185 ( .A(n23035), .ZN(n25792) );
  INV_X1 U19186 ( .A(n23034), .ZN(n25793) );
  INV_X1 U19187 ( .A(n23034), .ZN(n25794) );
  INV_X1 U19188 ( .A(n23035), .ZN(n25795) );
  INV_X1 U19189 ( .A(n25095), .ZN(n25796) );
  INV_X1 U19190 ( .A(n19022), .ZN(n25797) );
  INV_X1 U19191 ( .A(n27181), .ZN(n25798) );
  INV_X1 U19192 ( .A(n25798), .ZN(n25799) );
  INV_X1 U19193 ( .A(n25798), .ZN(n25800) );
  INV_X1 U19194 ( .A(n23037), .ZN(n25801) );
  INV_X1 U19195 ( .A(n23036), .ZN(n25802) );
  INV_X1 U19196 ( .A(n23036), .ZN(n25803) );
  INV_X1 U19197 ( .A(n23037), .ZN(n25804) );
  INV_X1 U19198 ( .A(n23039), .ZN(n25805) );
  INV_X1 U19199 ( .A(n23038), .ZN(n25806) );
  INV_X1 U19200 ( .A(n23038), .ZN(n25807) );
  INV_X1 U19201 ( .A(n23039), .ZN(n25808) );
  INV_X1 U19202 ( .A(n23041), .ZN(n25809) );
  INV_X1 U19203 ( .A(n23040), .ZN(n25810) );
  INV_X1 U19204 ( .A(n23041), .ZN(n25811) );
  INV_X1 U19205 ( .A(n23040), .ZN(n25812) );
  INV_X1 U19206 ( .A(n23043), .ZN(n25813) );
  INV_X1 U19207 ( .A(n23042), .ZN(n25814) );
  INV_X1 U19208 ( .A(n23043), .ZN(n25815) );
  INV_X1 U19209 ( .A(n23042), .ZN(n25816) );
  INV_X1 U19210 ( .A(n19026), .ZN(n25817) );
  INV_X1 U19211 ( .A(n25101), .ZN(n25818) );
  INV_X1 U19212 ( .A(n27185), .ZN(n25819) );
  INV_X1 U19213 ( .A(n25819), .ZN(n25820) );
  INV_X1 U19214 ( .A(n25819), .ZN(n25821) );
  INV_X1 U19215 ( .A(n23045), .ZN(n25822) );
  INV_X1 U19216 ( .A(n23044), .ZN(n25823) );
  INV_X1 U19217 ( .A(n23044), .ZN(n25824) );
  INV_X1 U19218 ( .A(n23045), .ZN(n25825) );
  INV_X1 U19219 ( .A(n23047), .ZN(n25826) );
  INV_X1 U19220 ( .A(n23046), .ZN(n25827) );
  INV_X1 U19221 ( .A(n23046), .ZN(n25828) );
  INV_X1 U19222 ( .A(n23047), .ZN(n25829) );
  INV_X1 U19223 ( .A(n20507), .ZN(n25830) );
  INV_X1 U19224 ( .A(n24730), .ZN(n25831) );
  CLKBUF_X1 U19225 ( .A(n20907), .Z(n25832) );
  INV_X1 U19226 ( .A(n25831), .ZN(n25833) );
  INV_X1 U19227 ( .A(n25833), .ZN(n25834) );
  INV_X1 U19228 ( .A(n25833), .ZN(n25835) );
  INV_X1 U19229 ( .A(n23048), .ZN(n25836) );
  INV_X1 U19230 ( .A(n23049), .ZN(n25837) );
  INV_X1 U19231 ( .A(n23048), .ZN(n25838) );
  INV_X1 U19232 ( .A(n23049), .ZN(n25839) );
  INV_X1 U19233 ( .A(n23050), .ZN(n25840) );
  INV_X1 U19234 ( .A(n23051), .ZN(n25841) );
  INV_X1 U19235 ( .A(n23050), .ZN(n25842) );
  INV_X1 U19236 ( .A(n23051), .ZN(n25843) );
  INV_X1 U19237 ( .A(n20511), .ZN(n25844) );
  INV_X1 U19238 ( .A(n24731), .ZN(n25845) );
  CLKBUF_X1 U19239 ( .A(n20902), .Z(n25846) );
  INV_X1 U19240 ( .A(n25845), .ZN(n25847) );
  INV_X1 U19241 ( .A(n25847), .ZN(n25848) );
  INV_X1 U19242 ( .A(n25847), .ZN(n25849) );
  INV_X1 U19243 ( .A(n23052), .ZN(n25850) );
  INV_X1 U19244 ( .A(n23053), .ZN(n25851) );
  INV_X1 U19245 ( .A(n23052), .ZN(n25852) );
  INV_X1 U19246 ( .A(n23053), .ZN(n25853) );
  INV_X1 U19247 ( .A(n23054), .ZN(n25854) );
  INV_X1 U19248 ( .A(n23055), .ZN(n25855) );
  INV_X1 U19249 ( .A(n23054), .ZN(n25856) );
  INV_X1 U19250 ( .A(n23055), .ZN(n25857) );
  INV_X1 U19251 ( .A(n23056), .ZN(n25858) );
  INV_X1 U19252 ( .A(n23057), .ZN(n25859) );
  INV_X1 U19253 ( .A(n23056), .ZN(n25860) );
  INV_X1 U19254 ( .A(n23057), .ZN(n25861) );
  INV_X1 U19255 ( .A(n23058), .ZN(n25862) );
  INV_X1 U19256 ( .A(n23059), .ZN(n25863) );
  INV_X1 U19257 ( .A(n23058), .ZN(n25864) );
  INV_X1 U19258 ( .A(n23059), .ZN(n25865) );
  INV_X1 U19259 ( .A(n23060), .ZN(n25866) );
  INV_X1 U19260 ( .A(n23061), .ZN(n25867) );
  INV_X1 U19261 ( .A(n23060), .ZN(n25868) );
  INV_X1 U19262 ( .A(n23061), .ZN(n25869) );
  CLKBUF_X1 U19263 ( .A(n20539), .Z(n27221) );
  INV_X1 U19264 ( .A(n21422), .ZN(n25870) );
  INV_X1 U19265 ( .A(n21422), .ZN(n25871) );
  INV_X1 U19266 ( .A(n23062), .ZN(n25872) );
  INV_X1 U19267 ( .A(n23062), .ZN(n25873) );
  INV_X1 U19268 ( .A(n23063), .ZN(n25874) );
  INV_X1 U19269 ( .A(n23063), .ZN(n25875) );
  INV_X1 U19270 ( .A(n23064), .ZN(n25876) );
  INV_X1 U19271 ( .A(n23065), .ZN(n25877) );
  INV_X1 U19272 ( .A(n23065), .ZN(n25878) );
  INV_X1 U19273 ( .A(n23064), .ZN(n25879) );
  INV_X1 U19274 ( .A(n23067), .ZN(n25880) );
  INV_X1 U19275 ( .A(n23067), .ZN(n25881) );
  INV_X1 U19276 ( .A(n23066), .ZN(n25882) );
  BUF_X1 U19277 ( .A(n25874), .Z(n25883) );
  INV_X1 U19278 ( .A(n23071), .ZN(n25884) );
  INV_X1 U19279 ( .A(n23072), .ZN(n25885) );
  INV_X1 U19280 ( .A(n23071), .ZN(n25886) );
  INV_X1 U19281 ( .A(n23072), .ZN(n25887) );
  INV_X1 U19282 ( .A(n23073), .ZN(n25888) );
  INV_X1 U19283 ( .A(n23074), .ZN(n25889) );
  INV_X1 U19284 ( .A(n23073), .ZN(n25890) );
  INV_X1 U19285 ( .A(n23074), .ZN(n25891) );
  INV_X1 U19286 ( .A(n21429), .ZN(n25892) );
  INV_X1 U19287 ( .A(n21429), .ZN(n25893) );
  INV_X1 U19288 ( .A(n24465), .ZN(n25894) );
  INV_X1 U19289 ( .A(n25894), .ZN(n25895) );
  INV_X1 U19290 ( .A(n23075), .ZN(n25896) );
  INV_X1 U19291 ( .A(n23076), .ZN(n25897) );
  INV_X1 U19292 ( .A(n23076), .ZN(n25898) );
  INV_X1 U19293 ( .A(n23075), .ZN(n25899) );
  INV_X1 U19294 ( .A(n23077), .ZN(n25900) );
  INV_X1 U19295 ( .A(n23078), .ZN(n25901) );
  INV_X1 U19296 ( .A(n23077), .ZN(n25902) );
  INV_X1 U19297 ( .A(n23078), .ZN(n25903) );
  CLKBUF_X1 U19298 ( .A(n26945), .Z(n25904) );
  INV_X1 U19299 ( .A(n26763), .ZN(n25905) );
  INV_X1 U19300 ( .A(n25905), .ZN(n25906) );
  INV_X1 U19301 ( .A(n25905), .ZN(n25907) );
  INV_X1 U19302 ( .A(n24430), .ZN(n26945) );
  INV_X1 U19303 ( .A(n24917), .ZN(n25908) );
  INV_X1 U19304 ( .A(n26758), .ZN(n25909) );
  INV_X1 U19305 ( .A(n25909), .ZN(n25910) );
  INV_X1 U19306 ( .A(n25909), .ZN(n25911) );
  INV_X1 U19307 ( .A(n20888), .ZN(n27739) );
  INV_X1 U19308 ( .A(n23080), .ZN(n25912) );
  INV_X1 U19309 ( .A(n23079), .ZN(n25913) );
  INV_X1 U19310 ( .A(n23080), .ZN(n25914) );
  INV_X1 U19311 ( .A(n23079), .ZN(n25915) );
  INV_X1 U19312 ( .A(n24915), .ZN(n25916) );
  INV_X1 U19313 ( .A(n24914), .ZN(n25917) );
  CLKBUF_X1 U19314 ( .A(n26947), .Z(n25918) );
  INV_X1 U19315 ( .A(n24431), .ZN(n26947) );
  INV_X1 U19316 ( .A(n23082), .ZN(n25919) );
  INV_X1 U19317 ( .A(n23081), .ZN(n259201) );
  INV_X1 U19318 ( .A(n23082), .ZN(n25921) );
  INV_X1 U19319 ( .A(n23081), .ZN(n25922) );
  INV_X1 U19320 ( .A(n23084), .ZN(n25923) );
  INV_X1 U19321 ( .A(n23083), .ZN(n25924) );
  INV_X1 U19322 ( .A(n23084), .ZN(n25925) );
  INV_X1 U19323 ( .A(n23083), .ZN(n25926) );
  INV_X1 U19324 ( .A(n23085), .ZN(n25927) );
  INV_X1 U19325 ( .A(n23086), .ZN(n25928) );
  INV_X1 U19326 ( .A(n23085), .ZN(n25929) );
  INV_X1 U19327 ( .A(n23086), .ZN(n259301) );
  INV_X1 U19328 ( .A(n23088), .ZN(n25931) );
  INV_X1 U19329 ( .A(n23087), .ZN(n25932) );
  INV_X1 U19330 ( .A(n23088), .ZN(n25933) );
  INV_X1 U19331 ( .A(n23087), .ZN(n25934) );
  INV_X1 U19332 ( .A(n23089), .ZN(n25935) );
  INV_X1 U19333 ( .A(n23090), .ZN(n25936) );
  INV_X1 U19334 ( .A(n23091), .ZN(n25937) );
  INV_X1 U19335 ( .A(n23092), .ZN(n25938) );
  INV_X1 U19336 ( .A(n23091), .ZN(n25939) );
  INV_X1 U19337 ( .A(n23092), .ZN(n259401) );
  INV_X1 U19338 ( .A(n17113), .ZN(n25941) );
  INV_X1 U19339 ( .A(n23093), .ZN(n25942) );
  INV_X1 U19340 ( .A(n17113), .ZN(n25943) );
  INV_X1 U19341 ( .A(n23093), .ZN(n25944) );
  INV_X1 U19342 ( .A(n23095), .ZN(n25945) );
  INV_X1 U19343 ( .A(n23094), .ZN(n25946) );
  INV_X1 U19344 ( .A(n23095), .ZN(n25947) );
  INV_X1 U19345 ( .A(n23094), .ZN(n25948) );
  INV_X1 U19346 ( .A(n23096), .ZN(n25949) );
  INV_X1 U19347 ( .A(n23097), .ZN(n259501) );
  INV_X1 U19348 ( .A(n23097), .ZN(n25951) );
  INV_X1 U19349 ( .A(n23096), .ZN(n25952) );
  INV_X1 U19350 ( .A(n23099), .ZN(n25953) );
  INV_X1 U19351 ( .A(n23098), .ZN(n25954) );
  INV_X1 U19352 ( .A(n23099), .ZN(n25955) );
  INV_X1 U19353 ( .A(n23098), .ZN(n25956) );
  INV_X1 U19354 ( .A(n23100), .ZN(n25957) );
  INV_X1 U19355 ( .A(n23102), .ZN(n25958) );
  INV_X1 U19356 ( .A(n23102), .ZN(n25959) );
  INV_X1 U19357 ( .A(n23101), .ZN(n259601) );
  INV_X1 U19358 ( .A(n23104), .ZN(n25961) );
  INV_X1 U19359 ( .A(n23104), .ZN(n25962) );
  INV_X1 U19360 ( .A(n23103), .ZN(n25963) );
  INV_X1 U19361 ( .A(n23105), .ZN(n25964) );
  INV_X1 U19362 ( .A(n23106), .ZN(n25965) );
  INV_X1 U19363 ( .A(n23106), .ZN(n25966) );
  INV_X1 U19364 ( .A(n23107), .ZN(n25967) );
  INV_X1 U19365 ( .A(n23108), .ZN(n25968) );
  INV_X1 U19366 ( .A(n23108), .ZN(n25969) );
  CLKBUF_X1 U19367 ( .A(n20495), .Z(n259701) );
  INV_X1 U19368 ( .A(n19250), .ZN(n25971) );
  INV_X1 U19369 ( .A(n19250), .ZN(n25972) );
  INV_X1 U19370 ( .A(n23113), .ZN(n25973) );
  INV_X1 U19371 ( .A(n23113), .ZN(n25974) );
  INV_X1 U19372 ( .A(n23116), .ZN(n25975) );
  INV_X1 U19373 ( .A(n23115), .ZN(n25976) );
  INV_X1 U19374 ( .A(n23116), .ZN(n25977) );
  CLKBUF_X1 U19375 ( .A(n20497), .Z(n25978) );
  INV_X1 U19376 ( .A(n19251), .ZN(n25979) );
  INV_X1 U19377 ( .A(n19251), .ZN(n259801) );
  INV_X1 U19378 ( .A(n23122), .ZN(n25981) );
  INV_X1 U19379 ( .A(n23121), .ZN(n25982) );
  INV_X1 U19380 ( .A(n23122), .ZN(n25983) );
  INV_X1 U19381 ( .A(n23124), .ZN(n25984) );
  INV_X1 U19382 ( .A(n23123), .ZN(n25985) );
  INV_X1 U19383 ( .A(n23124), .ZN(n25986) );
  INV_X1 U19384 ( .A(n23126), .ZN(n25987) );
  INV_X1 U19385 ( .A(n23125), .ZN(n25988) );
  INV_X1 U19386 ( .A(n23126), .ZN(n25989) );
  CLKBUF_X1 U19387 ( .A(n24704), .Z(n259901) );
  INV_X1 U19388 ( .A(n23134), .ZN(n25991) );
  INV_X1 U19389 ( .A(n23135), .ZN(n25992) );
  INV_X1 U19390 ( .A(n23135), .ZN(n25993) );
  CLKBUF_X1 U19391 ( .A(n24710), .Z(n25994) );
  INV_X1 U19392 ( .A(n23144), .ZN(n25995) );
  INV_X1 U19393 ( .A(n23144), .ZN(n25996) );
  INV_X1 U19394 ( .A(n23143), .ZN(n25997) );
  INV_X1 U19395 ( .A(n24896), .ZN(n25998) );
  CLKBUF_X1 U19396 ( .A(n24724), .Z(n25999) );
  INV_X1 U19397 ( .A(n23149), .ZN(n260001) );
  INV_X1 U19398 ( .A(n23148), .ZN(n26001) );
  INV_X1 U19399 ( .A(n23149), .ZN(n26002) );
  INV_X1 U19400 ( .A(n24894), .ZN(n26003) );
  INV_X1 U19401 ( .A(n24431), .ZN(n26946) );
  INV_X1 U19402 ( .A(n23151), .ZN(n26004) );
  INV_X1 U19403 ( .A(n23151), .ZN(n26005) );
  INV_X1 U19404 ( .A(n23150), .ZN(n26006) );
  INV_X1 U19405 ( .A(n20710), .ZN(n26007) );
  INV_X1 U19406 ( .A(n24900), .ZN(n26008) );
  BUF_X1 U19407 ( .A(n24724), .Z(n27196) );
  INV_X1 U19408 ( .A(n23156), .ZN(n26009) );
  INV_X1 U19409 ( .A(n23155), .ZN(n260101) );
  INV_X1 U19410 ( .A(n23156), .ZN(n26011) );
  INV_X1 U19411 ( .A(n24898), .ZN(n26012) );
  CLKBUF_X1 U19412 ( .A(n27217), .Z(n26013) );
  BUF_X1 U19413 ( .A(n24723), .Z(n27217) );
  INV_X1 U19414 ( .A(n23161), .ZN(n26014) );
  INV_X1 U19415 ( .A(n23160), .ZN(n26015) );
  INV_X1 U19416 ( .A(n23161), .ZN(n26016) );
  INV_X1 U19417 ( .A(n24904), .ZN(n26017) );
  BUF_X1 U19418 ( .A(n24722), .Z(n27218) );
  INV_X1 U19419 ( .A(n23166), .ZN(n26018) );
  INV_X1 U19420 ( .A(n23165), .ZN(n26019) );
  INV_X1 U19421 ( .A(n23166), .ZN(n260201) );
  INV_X1 U19422 ( .A(n24902), .ZN(n26021) );
  INV_X1 U19423 ( .A(n24907), .ZN(n26022) );
  INV_X1 U19424 ( .A(n20715), .ZN(n26023) );
  INV_X1 U19425 ( .A(n27172), .ZN(n26024) );
  INV_X1 U19426 ( .A(n21859), .ZN(n27799) );
  INV_X1 U19427 ( .A(n23175), .ZN(n26025) );
  INV_X1 U19428 ( .A(n23174), .ZN(n26026) );
  INV_X1 U19429 ( .A(n23175), .ZN(n26027) );
  INV_X1 U19430 ( .A(n23177), .ZN(n26028) );
  INV_X1 U19431 ( .A(n23176), .ZN(n26029) );
  INV_X1 U19432 ( .A(n23177), .ZN(n260301) );
  INV_X1 U19433 ( .A(n23179), .ZN(n26031) );
  INV_X1 U19434 ( .A(n23178), .ZN(n26032) );
  INV_X1 U19435 ( .A(n23179), .ZN(n26033) );
  INV_X1 U19436 ( .A(n24906), .ZN(n26034) );
  INV_X1 U19437 ( .A(n24910), .ZN(n26035) );
  INV_X1 U19438 ( .A(n20718), .ZN(n26036) );
  INV_X1 U19439 ( .A(n26035), .ZN(n26037) );
  INV_X1 U19440 ( .A(n26037), .ZN(n26038) );
  INV_X1 U19441 ( .A(n26037), .ZN(n26039) );
  INV_X1 U19442 ( .A(n23187), .ZN(n260401) );
  INV_X1 U19443 ( .A(n23186), .ZN(n26041) );
  INV_X1 U19444 ( .A(n23187), .ZN(n26042) );
  INV_X1 U19445 ( .A(n23188), .ZN(n26043) );
  INV_X1 U19446 ( .A(n23189), .ZN(n26044) );
  INV_X1 U19447 ( .A(n23189), .ZN(n26045) );
  INV_X1 U19448 ( .A(n24908), .ZN(n26046) );
  INV_X1 U19449 ( .A(n20717), .ZN(n26047) );
  INV_X1 U19450 ( .A(n27225), .ZN(n26048) );
  INV_X1 U19451 ( .A(n21861), .ZN(n27801) );
  INV_X1 U19452 ( .A(n23195), .ZN(n26049) );
  INV_X1 U19453 ( .A(n23194), .ZN(n260501) );
  INV_X1 U19454 ( .A(n23195), .ZN(n26051) );
  INV_X1 U19455 ( .A(n17112), .ZN(n26052) );
  INV_X1 U19456 ( .A(n27227), .ZN(n26053) );
  INV_X1 U19457 ( .A(n17112), .ZN(n26054) );
  INV_X1 U19458 ( .A(n23197), .ZN(n26055) );
  INV_X1 U19459 ( .A(n23196), .ZN(n26056) );
  INV_X1 U19460 ( .A(n23197), .ZN(n26057) );
  INV_X1 U19461 ( .A(n23199), .ZN(n26058) );
  INV_X1 U19462 ( .A(n23198), .ZN(n26059) );
  INV_X1 U19463 ( .A(n23199), .ZN(n260601) );
  INV_X1 U19464 ( .A(n23200), .ZN(n26061) );
  INV_X1 U19465 ( .A(n23201), .ZN(n26062) );
  INV_X1 U19466 ( .A(n23201), .ZN(n26063) );
  INV_X1 U19467 ( .A(n24912), .ZN(n26064) );
  CLKBUF_X1 U19468 ( .A(n26013), .Z(n26065) );
  INV_X1 U19469 ( .A(n23206), .ZN(n26066) );
  INV_X1 U19470 ( .A(n23205), .ZN(n26067) );
  INV_X1 U19471 ( .A(n23206), .ZN(n26068) );
  INV_X1 U19472 ( .A(n23208), .ZN(n26069) );
  INV_X1 U19473 ( .A(n23208), .ZN(n260701) );
  INV_X1 U19474 ( .A(n23207), .ZN(n26071) );
  INV_X1 U19475 ( .A(n23209), .ZN(n26072) );
  INV_X1 U19476 ( .A(n23210), .ZN(n26073) );
  INV_X1 U19477 ( .A(n23210), .ZN(n26074) );
  INV_X1 U19478 ( .A(n23211), .ZN(n26075) );
  INV_X1 U19479 ( .A(n23211), .ZN(n26076) );
  INV_X1 U19480 ( .A(n26549), .ZN(n26077) );
  INV_X1 U19481 ( .A(n23214), .ZN(n26078) );
  INV_X1 U19482 ( .A(n23213), .ZN(n26079) );
  INV_X1 U19483 ( .A(n23214), .ZN(n260801) );
  INV_X1 U19484 ( .A(n23215), .ZN(n26081) );
  INV_X1 U19485 ( .A(n23215), .ZN(n26082) );
  INV_X1 U19486 ( .A(n23216), .ZN(n26083) );
  INV_X1 U19487 ( .A(n17111), .ZN(n26084) );
  INV_X1 U19488 ( .A(n23217), .ZN(n26085) );
  INV_X1 U19489 ( .A(n23218), .ZN(n26086) );
  INV_X1 U19490 ( .A(n23219), .ZN(n26087) );
  INV_X1 U19491 ( .A(n23218), .ZN(n26088) );
  INV_X1 U19492 ( .A(n23221), .ZN(n26089) );
  INV_X1 U19493 ( .A(n23222), .ZN(n260901) );
  INV_X1 U19494 ( .A(n24696), .ZN(n26091) );
  INV_X1 U19495 ( .A(n23225), .ZN(n26092) );
  INV_X1 U19496 ( .A(n23224), .ZN(n26093) );
  INV_X1 U19497 ( .A(n23226), .ZN(n26094) );
  INV_X1 U19498 ( .A(n23228), .ZN(n26095) );
  INV_X1 U19499 ( .A(n23227), .ZN(n26096) );
  INV_X1 U19500 ( .A(n23229), .ZN(n26097) );
  INV_X1 U19501 ( .A(n23230), .ZN(n26098) );
  INV_X1 U19502 ( .A(n23229), .ZN(n26099) );
  INV_X1 U19503 ( .A(n23231), .ZN(n261001) );
  INV_X1 U19504 ( .A(n23232), .ZN(n26101) );
  INV_X1 U19505 ( .A(n24694), .ZN(n26102) );
  INV_X1 U19506 ( .A(n23235), .ZN(n26103) );
  INV_X1 U19507 ( .A(n23234), .ZN(n26104) );
  INV_X1 U19508 ( .A(n23236), .ZN(n26105) );
  INV_X1 U19509 ( .A(n23237), .ZN(n26106) );
  INV_X1 U19510 ( .A(n23238), .ZN(n26107) );
  INV_X1 U19511 ( .A(n23239), .ZN(n26108) );
  INV_X1 U19512 ( .A(n23242), .ZN(n26109) );
  INV_X1 U19513 ( .A(n23241), .ZN(n261101) );
  INV_X1 U19514 ( .A(n23244), .ZN(n26111) );
  INV_X1 U19515 ( .A(n23243), .ZN(n26112) );
  INV_X1 U19516 ( .A(n23246), .ZN(n26113) );
  INV_X1 U19517 ( .A(n23245), .ZN(n26114) );
  INV_X1 U19518 ( .A(n23248), .ZN(n26115) );
  INV_X1 U19519 ( .A(n23247), .ZN(n26116) );
  INV_X1 U19520 ( .A(n23250), .ZN(n26117) );
  INV_X1 U19521 ( .A(n23249), .ZN(n26118) );
  INV_X1 U19522 ( .A(n23252), .ZN(n26119) );
  INV_X1 U19523 ( .A(n23251), .ZN(n261201) );
  INV_X1 U19524 ( .A(n23254), .ZN(n26121) );
  INV_X1 U19525 ( .A(n23253), .ZN(n26122) );
  INV_X1 U19526 ( .A(n23257), .ZN(n26123) );
  INV_X1 U19527 ( .A(n23256), .ZN(n26124) );
  INV_X1 U19528 ( .A(n23259), .ZN(n26125) );
  INV_X1 U19529 ( .A(n23258), .ZN(n26126) );
  INV_X1 U19530 ( .A(n23261), .ZN(n26127) );
  INV_X1 U19531 ( .A(n23260), .ZN(n26128) );
  INV_X1 U19532 ( .A(n21600), .ZN(n26129) );
  INV_X1 U19533 ( .A(n26129), .ZN(n26130) );
  INV_X1 U19534 ( .A(n26129), .ZN(n26131) );
  INV_X1 U19535 ( .A(n26368), .ZN(n26132) );
  INV_X1 U19536 ( .A(n26132), .ZN(n26133) );
  INV_X1 U19537 ( .A(n26132), .ZN(n26134) );
  INV_X1 U19538 ( .A(n23263), .ZN(n26135) );
  INV_X1 U19539 ( .A(n23262), .ZN(n26136) );
  BUF_X1 U19540 ( .A(n21372), .Z(n26137) );
  BUF_X1 U19541 ( .A(n19236), .Z(n26138) );
  INV_X1 U19542 ( .A(n23271), .ZN(n26139) );
  INV_X1 U19543 ( .A(n23270), .ZN(n26140) );
  BUF_X1 U19544 ( .A(n21369), .Z(n26141) );
  BUF_X1 U19545 ( .A(n19235), .Z(n26142) );
  INV_X1 U19546 ( .A(n23278), .ZN(n26143) );
  INV_X1 U19547 ( .A(n23279), .ZN(n26144) );
  INV_X1 U19548 ( .A(n23281), .ZN(n26145) );
  INV_X1 U19549 ( .A(n23280), .ZN(n26146) );
  INV_X1 U19550 ( .A(n23282), .ZN(n26147) );
  INV_X1 U19551 ( .A(n23283), .ZN(n26148) );
  CLKBUF_X1 U19552 ( .A(n24703), .Z(n26149) );
  INV_X1 U19553 ( .A(n23289), .ZN(n26150) );
  INV_X1 U19554 ( .A(n23288), .ZN(n26151) );
  INV_X1 U19555 ( .A(n23290), .ZN(n26152) );
  INV_X1 U19556 ( .A(n23291), .ZN(n26153) );
  INV_X1 U19557 ( .A(n23293), .ZN(n26154) );
  INV_X1 U19558 ( .A(n23292), .ZN(n26155) );
  INV_X1 U19559 ( .A(n23295), .ZN(n26156) );
  INV_X1 U19560 ( .A(n23294), .ZN(n26157) );
  CLKBUF_X1 U19561 ( .A(n24709), .Z(n26158) );
  INV_X1 U19562 ( .A(n23301), .ZN(n26159) );
  INV_X1 U19563 ( .A(n23300), .ZN(n26160) );
  INV_X1 U19564 ( .A(n23301), .ZN(n26161) );
  INV_X1 U19565 ( .A(n23303), .ZN(n26162) );
  INV_X1 U19566 ( .A(n23302), .ZN(n26163) );
  INV_X1 U19567 ( .A(n23304), .ZN(n26164) );
  INV_X1 U19568 ( .A(n23305), .ZN(n26165) );
  INV_X1 U19569 ( .A(n23307), .ZN(n26166) );
  INV_X1 U19570 ( .A(n23306), .ZN(n26167) );
  INV_X1 U19571 ( .A(n23308), .ZN(n26168) );
  INV_X1 U19572 ( .A(n23309), .ZN(n26169) );
  INV_X1 U19573 ( .A(n23311), .ZN(n26170) );
  INV_X1 U19574 ( .A(n23310), .ZN(n26171) );
  INV_X1 U19575 ( .A(n23312), .ZN(n26172) );
  INV_X1 U19576 ( .A(n23313), .ZN(n26173) );
  INV_X1 U19577 ( .A(n23315), .ZN(n26174) );
  INV_X1 U19578 ( .A(n23314), .ZN(n26175) );
  INV_X1 U19579 ( .A(n23317), .ZN(n26176) );
  INV_X1 U19580 ( .A(n23316), .ZN(n26177) );
  INV_X1 U19581 ( .A(n23319), .ZN(n26178) );
  INV_X1 U19582 ( .A(n23318), .ZN(n26179) );
  INV_X1 U19583 ( .A(n23321), .ZN(n26180) );
  INV_X1 U19584 ( .A(n23320), .ZN(n26181) );
  INV_X1 U19585 ( .A(n23322), .ZN(n26182) );
  INV_X1 U19586 ( .A(n23323), .ZN(n26183) );
  INV_X1 U19587 ( .A(n23325), .ZN(n26184) );
  INV_X1 U19588 ( .A(n23324), .ZN(n26185) );
  INV_X1 U19589 ( .A(n23326), .ZN(n26186) );
  INV_X1 U19590 ( .A(n23327), .ZN(n26187) );
  INV_X1 U19591 ( .A(n23329), .ZN(n26188) );
  INV_X1 U19592 ( .A(n23328), .ZN(n26189) );
  INV_X1 U19593 ( .A(n23330), .ZN(n26190) );
  INV_X1 U19594 ( .A(n23331), .ZN(n26191) );
  INV_X1 U19595 ( .A(n24868), .ZN(n26192) );
  INV_X1 U19596 ( .A(n26192), .ZN(n26193) );
  INV_X1 U19597 ( .A(n26193), .ZN(n26194) );
  INV_X1 U19598 ( .A(n26193), .ZN(n26195) );
  BUF_X1 U19599 ( .A(n24726), .Z(n27206) );
  INV_X1 U19600 ( .A(n24866), .ZN(n26196) );
  INV_X1 U19601 ( .A(n26196), .ZN(n26197) );
  INV_X1 U19602 ( .A(n26197), .ZN(n26198) );
  INV_X1 U19603 ( .A(n26197), .ZN(n26199) );
  BUF_X1 U19604 ( .A(n24727), .Z(n27205) );
  INV_X1 U19605 ( .A(n24872), .ZN(n26200) );
  INV_X1 U19606 ( .A(n26200), .ZN(n26201) );
  INV_X1 U19607 ( .A(n26201), .ZN(n26202) );
  INV_X1 U19608 ( .A(n26201), .ZN(n26203) );
  INV_X1 U19609 ( .A(n24870), .ZN(n26204) );
  INV_X1 U19610 ( .A(n26204), .ZN(n26205) );
  INV_X1 U19611 ( .A(n26205), .ZN(n26206) );
  INV_X1 U19612 ( .A(n26205), .ZN(n26207) );
  INV_X1 U19613 ( .A(n23345), .ZN(n26208) );
  INV_X1 U19614 ( .A(n23344), .ZN(n26209) );
  INV_X1 U19615 ( .A(n23347), .ZN(n26210) );
  INV_X1 U19616 ( .A(n23346), .ZN(n26211) );
  INV_X1 U19617 ( .A(n23349), .ZN(n26212) );
  INV_X1 U19618 ( .A(n23348), .ZN(n26213) );
  INV_X1 U19619 ( .A(n23351), .ZN(n26214) );
  INV_X1 U19620 ( .A(n23350), .ZN(n26215) );
  INV_X1 U19621 ( .A(n23353), .ZN(n26216) );
  INV_X1 U19622 ( .A(n23352), .ZN(n26217) );
  INV_X1 U19623 ( .A(n23355), .ZN(n26218) );
  INV_X1 U19624 ( .A(n23354), .ZN(n26219) );
  INV_X1 U19625 ( .A(n23357), .ZN(n26220) );
  INV_X1 U19626 ( .A(n23356), .ZN(n26221) );
  INV_X1 U19627 ( .A(n23359), .ZN(n26222) );
  INV_X1 U19628 ( .A(n23358), .ZN(n26223) );
  INV_X1 U19629 ( .A(n23361), .ZN(n26224) );
  INV_X1 U19630 ( .A(n23360), .ZN(n26225) );
  INV_X1 U19631 ( .A(n23363), .ZN(n26226) );
  INV_X1 U19632 ( .A(n23362), .ZN(n26227) );
  INV_X1 U19633 ( .A(n23365), .ZN(n26228) );
  INV_X1 U19634 ( .A(n23364), .ZN(n26229) );
  INV_X1 U19635 ( .A(n23367), .ZN(n26230) );
  INV_X1 U19636 ( .A(n23366), .ZN(n26231) );
  INV_X1 U19637 ( .A(n23369), .ZN(n26232) );
  INV_X1 U19638 ( .A(n23368), .ZN(n26233) );
  INV_X1 U19639 ( .A(n23371), .ZN(n26234) );
  INV_X1 U19640 ( .A(n23370), .ZN(n26235) );
  INV_X1 U19641 ( .A(n23373), .ZN(n26236) );
  INV_X1 U19642 ( .A(n23372), .ZN(n26237) );
  INV_X1 U19643 ( .A(n23375), .ZN(n26238) );
  INV_X1 U19644 ( .A(n23374), .ZN(n26239) );
  INV_X1 U19645 ( .A(n24877), .ZN(n26240) );
  INV_X1 U19646 ( .A(n20703), .ZN(n26241) );
  INV_X1 U19647 ( .A(n19311), .ZN(n26242) );
  INV_X1 U19648 ( .A(n26242), .ZN(n26243) );
  INV_X1 U19649 ( .A(n26242), .ZN(n26244) );
  INV_X1 U19650 ( .A(n5297), .ZN(n277401) );
  INV_X1 U19651 ( .A(n24875), .ZN(n26245) );
  CLKBUF_X1 U19652 ( .A(n23389), .Z(n26246) );
  INV_X1 U19653 ( .A(n19262), .ZN(n26247) );
  INV_X1 U19654 ( .A(n26247), .ZN(n26248) );
  INV_X1 U19655 ( .A(n26247), .ZN(n26249) );
  INV_X1 U19656 ( .A(n23384), .ZN(n26250) );
  INV_X1 U19657 ( .A(n23383), .ZN(n26251) );
  INV_X1 U19658 ( .A(n23386), .ZN(n26252) );
  INV_X1 U19659 ( .A(n23385), .ZN(n26253) );
  INV_X1 U19660 ( .A(n24883), .ZN(n26254) );
  INV_X1 U19661 ( .A(n26246), .ZN(n26255) );
  INV_X1 U19662 ( .A(n26255), .ZN(n26256) );
  INV_X1 U19663 ( .A(n26255), .ZN(n26257) );
  BUF_X1 U19664 ( .A(n38050), .Z(n27171) );
  INV_X1 U19665 ( .A(n23391), .ZN(n26258) );
  INV_X1 U19666 ( .A(n23390), .ZN(n26259) );
  INV_X1 U19667 ( .A(n23393), .ZN(n26260) );
  INV_X1 U19668 ( .A(n23392), .ZN(n26261) );
  INV_X1 U19669 ( .A(n24880), .ZN(n26262) );
  CLKBUF_X1 U19670 ( .A(n23411), .Z(n26263) );
  INV_X1 U19671 ( .A(n19263), .ZN(n26264) );
  INV_X1 U19672 ( .A(n26264), .ZN(n26265) );
  INV_X1 U19673 ( .A(n26264), .ZN(n26266) );
  INV_X1 U19674 ( .A(n23398), .ZN(n26267) );
  INV_X1 U19675 ( .A(n23399), .ZN(n26268) );
  INV_X1 U19676 ( .A(n23401), .ZN(n26269) );
  INV_X1 U19677 ( .A(n23400), .ZN(n26270) );
  INV_X1 U19678 ( .A(n24888), .ZN(n26271) );
  INV_X1 U19679 ( .A(n26271), .ZN(n26272) );
  INV_X1 U19680 ( .A(n26272), .ZN(n26273) );
  INV_X1 U19681 ( .A(n26272), .ZN(n26274) );
  INV_X1 U19682 ( .A(n23406), .ZN(n26275) );
  INV_X1 U19683 ( .A(n23405), .ZN(n26276) );
  INV_X1 U19684 ( .A(n23408), .ZN(n26277) );
  INV_X1 U19685 ( .A(n23407), .ZN(n26278) );
  INV_X1 U19686 ( .A(n24886), .ZN(n26279) );
  INV_X1 U19687 ( .A(n26263), .ZN(n26280) );
  INV_X1 U19688 ( .A(n26280), .ZN(n26281) );
  INV_X1 U19689 ( .A(n26280), .ZN(n26282) );
  BUF_X1 U19690 ( .A(n3185), .Z(n27259) );
  INV_X1 U19691 ( .A(n23413), .ZN(n26283) );
  INV_X1 U19692 ( .A(n23412), .ZN(n26284) );
  INV_X1 U19693 ( .A(n23415), .ZN(n26285) );
  INV_X1 U19694 ( .A(n23414), .ZN(n26286) );
  INV_X1 U19695 ( .A(n24893), .ZN(n26287) );
  CLKBUF_X1 U19696 ( .A(n22493), .Z(n26288) );
  INV_X1 U19697 ( .A(n26287), .ZN(n26289) );
  INV_X1 U19698 ( .A(n26289), .ZN(n26290) );
  INV_X1 U19699 ( .A(n26289), .ZN(n26291) );
  INV_X1 U19700 ( .A(n23419), .ZN(n26292) );
  INV_X1 U19701 ( .A(n23420), .ZN(n26293) );
  INV_X1 U19702 ( .A(n23422), .ZN(n26294) );
  INV_X1 U19703 ( .A(n23421), .ZN(n26295) );
  INV_X1 U19704 ( .A(n24891), .ZN(n26296) );
  CLKBUF_X1 U19705 ( .A(n22493), .Z(n26297) );
  INV_X1 U19706 ( .A(n26296), .ZN(n26298) );
  INV_X1 U19707 ( .A(n26298), .ZN(n26299) );
  INV_X1 U19708 ( .A(n26298), .ZN(n26300) );
  INV_X1 U19709 ( .A(n23426), .ZN(n26301) );
  INV_X1 U19710 ( .A(n23425), .ZN(n26302) );
  INV_X1 U19711 ( .A(n23428), .ZN(n26303) );
  INV_X1 U19712 ( .A(n23427), .ZN(n26304) );
  INV_X1 U19713 ( .A(n23429), .ZN(n26305) );
  INV_X1 U19714 ( .A(n23430), .ZN(n26306) );
  INV_X1 U19715 ( .A(n23431), .ZN(n26307) );
  INV_X1 U19716 ( .A(n23432), .ZN(n26308) );
  INV_X1 U19717 ( .A(n23433), .ZN(n26309) );
  INV_X1 U19718 ( .A(n23434), .ZN(n26310) );
  INV_X1 U19719 ( .A(n23435), .ZN(n26311) );
  INV_X1 U19720 ( .A(n23436), .ZN(n26312) );
  INV_X1 U19721 ( .A(n23437), .ZN(n26313) );
  INV_X1 U19722 ( .A(n23438), .ZN(n26314) );
  INV_X1 U19723 ( .A(n23439), .ZN(n26315) );
  INV_X1 U19724 ( .A(n23440), .ZN(n26316) );
  INV_X1 U19725 ( .A(n23441), .ZN(n26317) );
  INV_X1 U19726 ( .A(n23442), .ZN(n26318) );
  INV_X1 U19727 ( .A(n23443), .ZN(n26319) );
  INV_X1 U19728 ( .A(n23444), .ZN(n26320) );
  INV_X1 U19729 ( .A(n19751), .ZN(n26321) );
  INV_X1 U19730 ( .A(n26321), .ZN(n26322) );
  INV_X1 U19731 ( .A(n23447), .ZN(n26323) );
  INV_X1 U19732 ( .A(n23447), .ZN(n26324) );
  INV_X1 U19733 ( .A(n23446), .ZN(n26325) );
  INV_X1 U19734 ( .A(n17110), .ZN(n26326) );
  INV_X1 U19735 ( .A(n17110), .ZN(n26327) );
  INV_X1 U19736 ( .A(n23448), .ZN(n26328) );
  BUF_X1 U19737 ( .A(n25646), .Z(n26329) );
  INV_X1 U19738 ( .A(n23452), .ZN(n26330) );
  INV_X1 U19739 ( .A(n23452), .ZN(n26331) );
  INV_X1 U19740 ( .A(n23453), .ZN(n26332) );
  INV_X1 U19741 ( .A(n23454), .ZN(n26333) );
  INV_X1 U19742 ( .A(n23454), .ZN(n26334) );
  INV_X1 U19743 ( .A(n23455), .ZN(n26335) );
  INV_X1 U19744 ( .A(n23456), .ZN(n26336) );
  INV_X1 U19745 ( .A(n23456), .ZN(n26337) );
  INV_X1 U19746 ( .A(n23457), .ZN(n26338) );
  INV_X1 U19747 ( .A(n23458), .ZN(n26339) );
  INV_X1 U19748 ( .A(n23458), .ZN(n26340) );
  INV_X1 U19749 ( .A(n23459), .ZN(n26341) );
  INV_X1 U19750 ( .A(n23460), .ZN(n26342) );
  INV_X1 U19751 ( .A(n23460), .ZN(n26343) );
  INV_X1 U19752 ( .A(n23461), .ZN(n26344) );
  INV_X1 U19753 ( .A(n23462), .ZN(n26345) );
  INV_X1 U19754 ( .A(n23462), .ZN(n26346) );
  INV_X1 U19755 ( .A(n23463), .ZN(n26347) );
  INV_X1 U19756 ( .A(n23464), .ZN(n26348) );
  INV_X1 U19757 ( .A(n23464), .ZN(n26349) );
  INV_X1 U19758 ( .A(n23465), .ZN(n26350) );
  INV_X1 U19759 ( .A(n23466), .ZN(n26351) );
  INV_X1 U19760 ( .A(n23466), .ZN(n26352) );
  INV_X1 U19761 ( .A(n23467), .ZN(n26353) );
  INV_X1 U19762 ( .A(n23468), .ZN(n26354) );
  INV_X1 U19763 ( .A(n23468), .ZN(n26355) );
  INV_X1 U19764 ( .A(n23469), .ZN(n26356) );
  INV_X1 U19765 ( .A(n23470), .ZN(n26357) );
  INV_X1 U19766 ( .A(n23470), .ZN(n26358) );
  INV_X1 U19767 ( .A(n23471), .ZN(n26359) );
  INV_X1 U19768 ( .A(n23472), .ZN(n26360) );
  INV_X1 U19769 ( .A(n23472), .ZN(n26361) );
  INV_X1 U19770 ( .A(n23473), .ZN(n26362) );
  INV_X1 U19771 ( .A(n23474), .ZN(n26363) );
  INV_X1 U19772 ( .A(n23474), .ZN(n26364) );
  INV_X1 U19773 ( .A(n23475), .ZN(n26365) );
  INV_X1 U19774 ( .A(n23476), .ZN(n26366) );
  INV_X1 U19775 ( .A(n23477), .ZN(n26367) );
  INV_X1 U19776 ( .A(n23476), .ZN(n26368) );
  INV_X1 U19777 ( .A(n23477), .ZN(n26369) );
  INV_X1 U19778 ( .A(n23478), .ZN(n263701) );
  INV_X1 U19779 ( .A(n23478), .ZN(n26371) );
  INV_X1 U19780 ( .A(n23479), .ZN(n26372) );
  INV_X1 U19781 ( .A(n23480), .ZN(n26373) );
  INV_X1 U19782 ( .A(n23481), .ZN(n26374) );
  INV_X1 U19783 ( .A(n23480), .ZN(n26375) );
  INV_X1 U19784 ( .A(n23481), .ZN(n26376) );
  INV_X1 U19785 ( .A(n23482), .ZN(n26377) );
  INV_X1 U19786 ( .A(n23483), .ZN(n26378) );
  INV_X1 U19787 ( .A(n23482), .ZN(n26379) );
  INV_X1 U19788 ( .A(n23483), .ZN(n26380) );
  INV_X1 U19789 ( .A(n23485), .ZN(n26381) );
  INV_X1 U19790 ( .A(n23485), .ZN(n26382) );
  INV_X1 U19791 ( .A(n23486), .ZN(n26383) );
  BUF_X1 U19792 ( .A(n24768), .Z(n26384) );
  BUF_X1 U19793 ( .A(n24773), .Z(n26385) );
  INV_X1 U19794 ( .A(n21953), .ZN(n26386) );
  INV_X1 U19795 ( .A(n21954), .ZN(n26387) );
  INV_X1 U19796 ( .A(n21953), .ZN(n26388) );
  INV_X1 U19797 ( .A(n23487), .ZN(n26389) );
  INV_X1 U19798 ( .A(n23487), .ZN(n26390) );
  INV_X1 U19799 ( .A(n23488), .ZN(n26391) );
  INV_X1 U19800 ( .A(n23490), .ZN(n26392) );
  INV_X1 U19801 ( .A(n23490), .ZN(n26393) );
  INV_X1 U19802 ( .A(n23491), .ZN(n26394) );
  INV_X1 U19803 ( .A(n19067), .ZN(n26395) );
  INV_X1 U19804 ( .A(n23494), .ZN(n26396) );
  INV_X1 U19805 ( .A(n23494), .ZN(n26397) );
  INV_X1 U19806 ( .A(n23495), .ZN(n26398) );
  INV_X1 U19807 ( .A(n23496), .ZN(n26399) );
  INV_X1 U19808 ( .A(n23496), .ZN(n26400) );
  INV_X1 U19809 ( .A(n23497), .ZN(n26401) );
  INV_X1 U19810 ( .A(n23498), .ZN(n26402) );
  INV_X1 U19811 ( .A(n23498), .ZN(n26403) );
  INV_X1 U19812 ( .A(n23499), .ZN(n26404) );
  INV_X1 U19813 ( .A(n23501), .ZN(n26405) );
  INV_X1 U19814 ( .A(n23503), .ZN(n26406) );
  INV_X1 U19815 ( .A(n23505), .ZN(n26407) );
  INV_X1 U19816 ( .A(n23507), .ZN(n26408) );
  INV_X1 U19817 ( .A(n23509), .ZN(n26409) );
  INV_X1 U19818 ( .A(n23511), .ZN(n264101) );
  INV_X1 U19819 ( .A(n23513), .ZN(n26411) );
  INV_X1 U19820 ( .A(n23515), .ZN(n26412) );
  INV_X1 U19821 ( .A(n23517), .ZN(n26413) );
  INV_X1 U19822 ( .A(n23519), .ZN(n26414) );
  INV_X1 U19823 ( .A(n23521), .ZN(n26415) );
  INV_X1 U19824 ( .A(n23523), .ZN(n26416) );
  INV_X1 U19825 ( .A(n23525), .ZN(n26417) );
  INV_X1 U19826 ( .A(n23527), .ZN(n26418) );
  INV_X1 U19827 ( .A(n23529), .ZN(n26419) );
  INV_X1 U19828 ( .A(n23531), .ZN(n264201) );
  INV_X1 U19829 ( .A(n23533), .ZN(n26421) );
  INV_X1 U19830 ( .A(n23535), .ZN(n26422) );
  INV_X1 U19831 ( .A(n23537), .ZN(n26423) );
  INV_X1 U19832 ( .A(n23539), .ZN(n26424) );
  INV_X1 U19833 ( .A(n23541), .ZN(n26425) );
  INV_X1 U19834 ( .A(n23543), .ZN(n26426) );
  INV_X1 U19835 ( .A(n23545), .ZN(n26427) );
  INV_X1 U19836 ( .A(n23547), .ZN(n26428) );
  INV_X1 U19837 ( .A(n23549), .ZN(n26429) );
  INV_X1 U19838 ( .A(n23552), .ZN(n264301) );
  INV_X1 U19839 ( .A(n23552), .ZN(n26431) );
  INV_X1 U19840 ( .A(n23554), .ZN(n26432) );
  INV_X1 U19841 ( .A(n23555), .ZN(n26433) );
  INV_X1 U19842 ( .A(n23554), .ZN(n26434) );
  INV_X1 U19843 ( .A(n23555), .ZN(n26435) );
  INV_X1 U19844 ( .A(n23557), .ZN(n26436) );
  INV_X1 U19845 ( .A(n23557), .ZN(n26437) );
  INV_X1 U19846 ( .A(n23559), .ZN(n26438) );
  INV_X1 U19847 ( .A(n23560), .ZN(n26439) );
  INV_X1 U19848 ( .A(n23559), .ZN(n264401) );
  INV_X1 U19849 ( .A(n23560), .ZN(n26441) );
  INV_X1 U19850 ( .A(n23562), .ZN(n26442) );
  INV_X1 U19851 ( .A(n23563), .ZN(n26443) );
  INV_X1 U19852 ( .A(n23562), .ZN(n26444) );
  INV_X1 U19853 ( .A(n23563), .ZN(n26445) );
  INV_X1 U19854 ( .A(n23565), .ZN(n26446) );
  INV_X1 U19855 ( .A(n23567), .ZN(n26447) );
  INV_X1 U19856 ( .A(n23569), .ZN(n26448) );
  INV_X1 U19857 ( .A(n23571), .ZN(n26449) );
  INV_X1 U19858 ( .A(n23573), .ZN(n264501) );
  INV_X1 U19859 ( .A(n23575), .ZN(n26451) );
  INV_X1 U19860 ( .A(n23577), .ZN(n26452) );
  INV_X1 U19861 ( .A(n23579), .ZN(n26453) );
  INV_X1 U19862 ( .A(n23581), .ZN(n26454) );
  INV_X1 U19863 ( .A(n23588), .ZN(n26455) );
  INV_X1 U19864 ( .A(n23589), .ZN(n26456) );
  INV_X1 U19865 ( .A(n23589), .ZN(n26457) );
  INV_X1 U19866 ( .A(n23590), .ZN(n26458) );
  INV_X1 U19867 ( .A(n23591), .ZN(n26459) );
  INV_X1 U19868 ( .A(n23591), .ZN(n264601) );
  INV_X1 U19869 ( .A(n23592), .ZN(n26461) );
  INV_X1 U19870 ( .A(n23593), .ZN(n26462) );
  INV_X1 U19871 ( .A(n23593), .ZN(n26463) );
  INV_X1 U19872 ( .A(n23594), .ZN(n26464) );
  INV_X1 U19873 ( .A(n23595), .ZN(n26465) );
  INV_X1 U19874 ( .A(n23595), .ZN(n26466) );
  INV_X1 U19875 ( .A(n23596), .ZN(n26467) );
  INV_X1 U19876 ( .A(n23597), .ZN(n26468) );
  INV_X1 U19877 ( .A(n23597), .ZN(n26469) );
  INV_X1 U19878 ( .A(n23598), .ZN(n264701) );
  INV_X1 U19879 ( .A(n23599), .ZN(n26471) );
  INV_X1 U19880 ( .A(n23599), .ZN(n26472) );
  INV_X1 U19881 ( .A(n23600), .ZN(n26473) );
  INV_X1 U19882 ( .A(n23601), .ZN(n26474) );
  INV_X1 U19883 ( .A(n23601), .ZN(n26475) );
  INV_X1 U19884 ( .A(n23602), .ZN(n26476) );
  INV_X1 U19885 ( .A(n23603), .ZN(n26477) );
  INV_X1 U19886 ( .A(n23603), .ZN(n26478) );
  INV_X1 U19887 ( .A(n23604), .ZN(n26479) );
  INV_X1 U19888 ( .A(n23606), .ZN(n264801) );
  INV_X1 U19889 ( .A(n23608), .ZN(n26481) );
  INV_X1 U19890 ( .A(n23610), .ZN(n26482) );
  INV_X1 U19891 ( .A(n23612), .ZN(n26483) );
  INV_X1 U19892 ( .A(n23614), .ZN(n26484) );
  INV_X1 U19893 ( .A(n23616), .ZN(n26485) );
  INV_X1 U19894 ( .A(n23618), .ZN(n26486) );
  INV_X1 U19895 ( .A(n23620), .ZN(n26487) );
  INV_X1 U19896 ( .A(n23622), .ZN(n26488) );
  INV_X1 U19897 ( .A(n23624), .ZN(n26489) );
  INV_X1 U19898 ( .A(n23626), .ZN(n264901) );
  INV_X1 U19899 ( .A(n23628), .ZN(n26491) );
  INV_X1 U19900 ( .A(n23630), .ZN(n26492) );
  INV_X1 U19901 ( .A(n23632), .ZN(n26493) );
  INV_X1 U19902 ( .A(n23634), .ZN(n26494) );
  INV_X1 U19903 ( .A(n23636), .ZN(n26495) );
  INV_X1 U19904 ( .A(n23637), .ZN(n26496) );
  INV_X1 U19905 ( .A(n23637), .ZN(n26497) );
  INV_X1 U19906 ( .A(n23638), .ZN(n26498) );
  INV_X1 U19907 ( .A(n23639), .ZN(n26499) );
  INV_X1 U19908 ( .A(n23639), .ZN(n265001) );
  INV_X1 U19909 ( .A(n23640), .ZN(n26501) );
  INV_X1 U19910 ( .A(n23641), .ZN(n26502) );
  INV_X1 U19911 ( .A(n23641), .ZN(n26503) );
  INV_X1 U19912 ( .A(n23642), .ZN(n26504) );
  INV_X1 U19913 ( .A(n23644), .ZN(n26505) );
  INV_X1 U19914 ( .A(n23645), .ZN(n26506) );
  INV_X1 U19915 ( .A(n23646), .ZN(n26507) );
  INV_X1 U19916 ( .A(n23646), .ZN(n26508) );
  INV_X1 U19917 ( .A(n23647), .ZN(n26509) );
  INV_X1 U19918 ( .A(n23648), .ZN(n265101) );
  INV_X1 U19919 ( .A(n23648), .ZN(n26511) );
  INV_X1 U19920 ( .A(n23649), .ZN(n26512) );
  INV_X1 U19921 ( .A(n19751), .ZN(n26513) );
  INV_X1 U19922 ( .A(n23651), .ZN(n26514) );
  INV_X1 U19923 ( .A(n23651), .ZN(n26515) );
  INV_X1 U19924 ( .A(n23653), .ZN(n26516) );
  INV_X1 U19925 ( .A(n23653), .ZN(n26517) );
  INV_X1 U19926 ( .A(n23652), .ZN(n26518) );
  INV_X1 U19927 ( .A(n23652), .ZN(n26519) );
  INV_X1 U19928 ( .A(n26990), .ZN(n265201) );
  INV_X1 U19929 ( .A(n23656), .ZN(n26521) );
  INV_X1 U19930 ( .A(n23656), .ZN(n26522) );
  INV_X1 U19931 ( .A(n23655), .ZN(n26523) );
  INV_X1 U19932 ( .A(n23655), .ZN(n26524) );
  INV_X1 U19933 ( .A(n23658), .ZN(n26525) );
  INV_X1 U19934 ( .A(n30950), .ZN(n26526) );
  INV_X1 U19935 ( .A(n23660), .ZN(n26527) );
  INV_X1 U19936 ( .A(n23661), .ZN(n26528) );
  INV_X1 U19937 ( .A(n23661), .ZN(n26529) );
  INV_X1 U19938 ( .A(n23660), .ZN(n265301) );
  INV_X1 U19939 ( .A(n26989), .ZN(n26531) );
  INV_X1 U19940 ( .A(n23664), .ZN(n26532) );
  INV_X1 U19941 ( .A(n23664), .ZN(n26533) );
  INV_X1 U19942 ( .A(n23663), .ZN(n26534) );
  INV_X1 U19943 ( .A(n23663), .ZN(n26535) );
  INV_X1 U19944 ( .A(n23665), .ZN(n26536) );
  INV_X1 U19945 ( .A(n23665), .ZN(n26537) );
  INV_X1 U19946 ( .A(n23666), .ZN(n26538) );
  INV_X1 U19947 ( .A(n23666), .ZN(n26539) );
  INV_X1 U19948 ( .A(n19270), .ZN(n265401) );
  INV_X1 U19949 ( .A(n19270), .ZN(n26541) );
  BUF_X1 U19950 ( .A(n24698), .Z(n27204) );
  BUF_X1 U19951 ( .A(n24697), .Z(n27203) );
  INV_X1 U19952 ( .A(n23675), .ZN(n26542) );
  INV_X1 U19953 ( .A(n23674), .ZN(n26543) );
  INV_X1 U19954 ( .A(n23675), .ZN(n26544) );
  INV_X1 U19955 ( .A(n23674), .ZN(n26545) );
  INV_X1 U19956 ( .A(n22492), .ZN(n26546) );
  INV_X1 U19957 ( .A(n27204), .ZN(n26547) );
  INV_X1 U19958 ( .A(n23672), .ZN(n26548) );
  INV_X1 U19959 ( .A(n26988), .ZN(n26549) );
  INV_X1 U19960 ( .A(n23677), .ZN(n265501) );
  INV_X1 U19961 ( .A(n23677), .ZN(n26551) );
  INV_X1 U19962 ( .A(n17268), .ZN(n26552) );
  INV_X1 U19963 ( .A(n23682), .ZN(n26553) );
  INV_X1 U19964 ( .A(n23683), .ZN(n26554) );
  INV_X1 U19965 ( .A(n23682), .ZN(n26555) );
  INV_X1 U19966 ( .A(n23687), .ZN(n26556) );
  INV_X1 U19967 ( .A(n23688), .ZN(n26557) );
  INV_X1 U19968 ( .A(n23687), .ZN(n26558) );
  INV_X1 U19969 ( .A(n23688), .ZN(n26559) );
  BUF_X1 U19970 ( .A(n21863), .Z(n265601) );
  BUF_X1 U19971 ( .A(n21862), .Z(n26561) );
  INV_X1 U19972 ( .A(n23692), .ZN(n26562) );
  INV_X1 U19973 ( .A(n23693), .ZN(n26563) );
  INV_X1 U19974 ( .A(n23692), .ZN(n26564) );
  INV_X1 U19975 ( .A(n23693), .ZN(n26565) );
  INV_X1 U19976 ( .A(n23697), .ZN(n26566) );
  INV_X1 U19977 ( .A(n23698), .ZN(n26567) );
  INV_X1 U19978 ( .A(n23697), .ZN(n26568) );
  INV_X1 U19979 ( .A(n23698), .ZN(n26569) );
  INV_X1 U19980 ( .A(n23702), .ZN(n26570) );
  INV_X1 U19981 ( .A(n23703), .ZN(n26571) );
  INV_X1 U19982 ( .A(n23702), .ZN(n26572) );
  INV_X1 U19983 ( .A(n23703), .ZN(n26573) );
  BUF_X1 U19984 ( .A(n21860), .Z(n26574) );
  INV_X1 U19985 ( .A(n23707), .ZN(n26575) );
  INV_X1 U19986 ( .A(n23708), .ZN(n26576) );
  INV_X1 U19987 ( .A(n23707), .ZN(n26577) );
  INV_X1 U19988 ( .A(n23708), .ZN(n26578) );
  INV_X1 U19989 ( .A(n23712), .ZN(n26579) );
  INV_X1 U19990 ( .A(n23713), .ZN(n26580) );
  INV_X1 U19991 ( .A(n23712), .ZN(n26581) );
  INV_X1 U19992 ( .A(n23713), .ZN(n26582) );
  INV_X1 U19993 ( .A(n24813), .ZN(n26583) );
  INV_X1 U19994 ( .A(n269401), .ZN(n26584) );
  INV_X1 U19995 ( .A(n26584), .ZN(n26585) );
  INV_X1 U19996 ( .A(n23722), .ZN(n26586) );
  INV_X1 U19997 ( .A(n23723), .ZN(n26587) );
  INV_X1 U19998 ( .A(n23723), .ZN(n26588) );
  INV_X1 U19999 ( .A(n23722), .ZN(n26589) );
  CLKBUF_X1 U20000 ( .A(n277801), .Z(n26590) );
  INV_X1 U20001 ( .A(n4721), .ZN(n277801) );
  INV_X1 U20002 ( .A(n23731), .ZN(n26591) );
  INV_X1 U20003 ( .A(n23731), .ZN(n26592) );
  INV_X1 U20004 ( .A(n27296), .ZN(n26593) );
  INV_X1 U20005 ( .A(n18720), .ZN(n26594) );
  INV_X1 U20006 ( .A(n18720), .ZN(n26595) );
  CLKBUF_X1 U20007 ( .A(n26953), .Z(n26596) );
  INV_X1 U20008 ( .A(n24435), .ZN(n26953) );
  CLKBUF_X1 U20009 ( .A(n26954), .Z(n26597) );
  INV_X1 U20010 ( .A(n24436), .ZN(n26954) );
  CLKBUF_X1 U20011 ( .A(n26955), .Z(n26598) );
  INV_X1 U20012 ( .A(n24436), .ZN(n26955) );
  CLKBUF_X1 U20013 ( .A(n26956), .Z(n26599) );
  INV_X1 U20014 ( .A(n24435), .ZN(n26956) );
  CLKBUF_X1 U20015 ( .A(n26957), .Z(n26600) );
  INV_X1 U20016 ( .A(n24437), .ZN(n26957) );
  CLKBUF_X1 U20017 ( .A(n26958), .Z(n26601) );
  INV_X1 U20018 ( .A(n24438), .ZN(n26958) );
  CLKBUF_X1 U20019 ( .A(n26959), .Z(n26602) );
  INV_X1 U20020 ( .A(n24438), .ZN(n26959) );
  CLKBUF_X1 U20021 ( .A(n26960), .Z(n26603) );
  INV_X1 U20022 ( .A(n24437), .ZN(n26960) );
  INV_X1 U20023 ( .A(n23938), .ZN(n26604) );
  INV_X1 U20024 ( .A(n23942), .ZN(n26605) );
  INV_X1 U20025 ( .A(n23948), .ZN(n26606) );
  INV_X1 U20026 ( .A(n23947), .ZN(n26607) );
  INV_X1 U20027 ( .A(n23948), .ZN(n26608) );
  INV_X1 U20028 ( .A(n23947), .ZN(n26609) );
  INV_X1 U20029 ( .A(r899_B_4_), .ZN(n26610) );
  INV_X1 U20030 ( .A(n18819), .ZN(n26611) );
  INV_X1 U20031 ( .A(n18819), .ZN(n26612) );
  INV_X1 U20032 ( .A(n26610), .ZN(n26613) );
  INV_X1 U20033 ( .A(n26962), .ZN(n26614) );
  CLKBUF_X1 U20034 ( .A(n26975), .Z(n26616) );
  BUF_X1 U20035 ( .A(n27782), .Z(n26975) );
  CLKBUF_X1 U20036 ( .A(n27781), .Z(n26618) );
  INV_X1 U20037 ( .A(n25024), .ZN(n26619) );
  INV_X1 U20038 ( .A(n26619), .ZN(n26620) );
  INV_X1 U20039 ( .A(n19237), .ZN(n27781) );
  INV_X1 U20040 ( .A(n22680), .ZN(n26621) );
  INV_X1 U20041 ( .A(n22680), .ZN(n26622) );
  INV_X1 U20042 ( .A(n22681), .ZN(n26623) );
  INV_X1 U20043 ( .A(n22681), .ZN(n26624) );
  INV_X1 U20044 ( .A(n24419), .ZN(n26625) );
  INV_X1 U20045 ( .A(n25019), .ZN(n26626) );
  INV_X1 U20046 ( .A(n26626), .ZN(n26627) );
  BUF_X1 U20047 ( .A(n3161), .Z(n27260) );
  INV_X1 U20048 ( .A(n22687), .ZN(n26628) );
  INV_X1 U20049 ( .A(n22687), .ZN(n26629) );
  INV_X1 U20050 ( .A(n22688), .ZN(n26630) );
  INV_X1 U20051 ( .A(n22688), .ZN(n26631) );
  INV_X1 U20052 ( .A(n22689), .ZN(n26632) );
  INV_X1 U20053 ( .A(n22689), .ZN(n26633) );
  INV_X1 U20054 ( .A(n24415), .ZN(n26634) );
  INV_X1 U20055 ( .A(n22693), .ZN(n26635) );
  INV_X1 U20056 ( .A(n22693), .ZN(n26636) );
  INV_X1 U20057 ( .A(r899_B_9_), .ZN(n26637) );
  INV_X1 U20058 ( .A(n45500), .ZN(n26638) );
  INV_X1 U20059 ( .A(n22696), .ZN(n26639) );
  INV_X1 U20060 ( .A(n3079), .ZN(n26640) );
  INV_X1 U20061 ( .A(n22700), .ZN(n26641) );
  INV_X1 U20062 ( .A(n22703), .ZN(n26642) );
  INV_X1 U20063 ( .A(n22706), .ZN(n26643) );
  INV_X1 U20064 ( .A(n47060), .ZN(n26644) );
  INV_X1 U20065 ( .A(n22710), .ZN(n26645) );
  BUF_X1 U20066 ( .A(n21398), .Z(n26646) );
  INV_X1 U20067 ( .A(n22713), .ZN(n26647) );
  INV_X1 U20068 ( .A(n22716), .ZN(n26648) );
  INV_X1 U20069 ( .A(n22719), .ZN(n26649) );
  INV_X1 U20070 ( .A(n22722), .ZN(n26650) );
  BUF_X1 U20071 ( .A(n25661), .Z(n26651) );
  INV_X1 U20072 ( .A(n19288), .ZN(n26652) );
  INV_X1 U20073 ( .A(n19288), .ZN(n26653) );
  INV_X1 U20074 ( .A(n22729), .ZN(n26654) );
  INV_X1 U20075 ( .A(n20611), .ZN(n26655) );
  INV_X1 U20076 ( .A(n24815), .ZN(n26656) );
  CLKBUF_X1 U20077 ( .A(n26961), .Z(n26657) );
  INV_X1 U20078 ( .A(n24440), .ZN(n26961) );
  INV_X1 U20079 ( .A(n20618), .ZN(n26658) );
  INV_X1 U20080 ( .A(n24819), .ZN(n26659) );
  CLKBUF_X1 U20081 ( .A(n26963), .Z(n26660) );
  INV_X1 U20082 ( .A(n24439), .ZN(n26963) );
  INV_X1 U20083 ( .A(n24818), .ZN(n26661) );
  INV_X1 U20084 ( .A(n20615), .ZN(n26662) );
  CLKBUF_X1 U20085 ( .A(n26964), .Z(n26663) );
  INV_X1 U20086 ( .A(n24440), .ZN(n26964) );
  INV_X1 U20087 ( .A(n22732), .ZN(n26664) );
  INV_X1 U20088 ( .A(n22732), .ZN(n26665) );
  INV_X1 U20089 ( .A(n4819), .ZN(n26666) );
  INV_X1 U20090 ( .A(n22737), .ZN(n26667) );
  INV_X1 U20091 ( .A(n22737), .ZN(n26668) );
  INV_X1 U20092 ( .A(n47050), .ZN(n26669) );
  INV_X1 U20093 ( .A(n22742), .ZN(n26670) );
  INV_X1 U20094 ( .A(n22742), .ZN(n26671) );
  INV_X1 U20095 ( .A(n22747), .ZN(n26672) );
  INV_X1 U20096 ( .A(n22751), .ZN(n26673) );
  INV_X1 U20097 ( .A(n24106), .ZN(n26674) );
  BUF_X1 U20098 ( .A(n25648), .Z(n26675) );
  INV_X1 U20099 ( .A(n22754), .ZN(n26676) );
  INV_X1 U20100 ( .A(n22754), .ZN(n26677) );
  INV_X1 U20101 ( .A(n24142), .ZN(n26678) );
  INV_X1 U20102 ( .A(n24142), .ZN(n26679) );
  INV_X1 U20103 ( .A(n24143), .ZN(n26680) );
  INV_X1 U20104 ( .A(n24143), .ZN(n26681) );
  INV_X1 U20105 ( .A(n24144), .ZN(n26682) );
  INV_X1 U20106 ( .A(n24144), .ZN(n26683) );
  INV_X1 U20107 ( .A(n24145), .ZN(n26684) );
  INV_X1 U20108 ( .A(n24145), .ZN(n26685) );
  INV_X1 U20109 ( .A(n22764), .ZN(n26686) );
  INV_X1 U20110 ( .A(n22764), .ZN(n26687) );
  BUF_X1 U20111 ( .A(n19226), .Z(n26688) );
  BUF_X1 U20112 ( .A(n17082), .Z(n26689) );
  BUF_X1 U20113 ( .A(n19229), .Z(n26690) );
  BUF_X1 U20114 ( .A(n25634), .Z(n26691) );
  INV_X1 U20115 ( .A(n24146), .ZN(n26692) );
  INV_X1 U20116 ( .A(n24146), .ZN(n26693) );
  INV_X1 U20117 ( .A(n24147), .ZN(n26694) );
  INV_X1 U20118 ( .A(n24147), .ZN(n26695) );
  INV_X1 U20119 ( .A(n22771), .ZN(n26696) );
  INV_X1 U20120 ( .A(n22771), .ZN(n26697) );
  INV_X1 U20121 ( .A(n24148), .ZN(n26698) );
  INV_X1 U20122 ( .A(n24148), .ZN(n26699) );
  INV_X1 U20123 ( .A(n24149), .ZN(n26700) );
  INV_X1 U20124 ( .A(n24149), .ZN(n26701) );
  INV_X1 U20125 ( .A(n27789), .ZN(n26702) );
  INV_X1 U20126 ( .A(n22779), .ZN(n26704) );
  INV_X1 U20127 ( .A(n27726), .ZN(n26705) );
  INV_X1 U20128 ( .A(n22781), .ZN(n26707) );
  INV_X1 U20129 ( .A(n4714), .ZN(n26708) );
  INV_X1 U20130 ( .A(n22783), .ZN(n26710) );
  INV_X1 U20131 ( .A(n22785), .ZN(n26711) );
  INV_X1 U20132 ( .A(n4713), .ZN(n26712) );
  INV_X1 U20133 ( .A(n22789), .ZN(n26714) );
  INV_X1 U20134 ( .A(n24170), .ZN(n26715) );
  INV_X1 U20135 ( .A(n24172), .ZN(n26716) );
  INV_X1 U20136 ( .A(n24172), .ZN(n26717) );
  INV_X1 U20137 ( .A(n24175), .ZN(n26718) );
  INV_X1 U20138 ( .A(n24175), .ZN(n26719) );
  INV_X1 U20139 ( .A(n24180), .ZN(n26721) );
  INV_X1 U20140 ( .A(n24180), .ZN(n26722) );
  INV_X1 U20141 ( .A(n24184), .ZN(n26724) );
  INV_X1 U20142 ( .A(n24184), .ZN(n26726) );
  BUF_X1 U20143 ( .A(n25875), .Z(n26727) );
  BUF_X1 U20144 ( .A(n25873), .Z(n26728) );
  INV_X1 U20145 ( .A(n22798), .ZN(n26729) );
  INV_X1 U20146 ( .A(n22808), .ZN(n26730) );
  INV_X1 U20147 ( .A(n22810), .ZN(n26731) );
  INV_X1 U20148 ( .A(n24202), .ZN(n26732) );
  INV_X1 U20149 ( .A(n24202), .ZN(n26733) );
  INV_X1 U20150 ( .A(n24201), .ZN(n26735) );
  INV_X1 U20151 ( .A(n24918), .ZN(n26736) );
  INV_X1 U20152 ( .A(n20722), .ZN(n26737) );
  INV_X1 U20153 ( .A(n24918), .ZN(n26738) );
  INV_X1 U20154 ( .A(n24208), .ZN(n26739) );
  INV_X1 U20155 ( .A(n24208), .ZN(n267401) );
  INV_X1 U20156 ( .A(n24207), .ZN(n26742) );
  INV_X1 U20157 ( .A(n24920), .ZN(n26743) );
  INV_X1 U20158 ( .A(n24920), .ZN(n26744) );
  INV_X1 U20159 ( .A(n24919), .ZN(n26745) );
  INV_X1 U20160 ( .A(n24212), .ZN(n26746) );
  INV_X1 U20161 ( .A(n24212), .ZN(n26747) );
  INV_X1 U20162 ( .A(n22820), .ZN(n26748) );
  INV_X1 U20163 ( .A(n22820), .ZN(n267501) );
  INV_X1 U20164 ( .A(n22823), .ZN(n26751) );
  INV_X1 U20165 ( .A(n22823), .ZN(n26753) );
  INV_X1 U20166 ( .A(n24915), .ZN(n26754) );
  INV_X1 U20167 ( .A(n24914), .ZN(n26755) );
  INV_X1 U20168 ( .A(n20721), .ZN(n26756) );
  INV_X1 U20169 ( .A(n20721), .ZN(n26757) );
  INV_X1 U20170 ( .A(n24917), .ZN(n26758) );
  INV_X1 U20171 ( .A(n24722), .ZN(n26759) );
  INV_X1 U20172 ( .A(n20719), .ZN(n267601) );
  INV_X1 U20173 ( .A(n24912), .ZN(n26761) );
  INV_X1 U20174 ( .A(n20720), .ZN(n26762) );
  INV_X1 U20175 ( .A(n20720), .ZN(n26763) );
  INV_X1 U20176 ( .A(n24908), .ZN(n26764) );
  INV_X1 U20177 ( .A(n24725), .ZN(n26765) );
  INV_X1 U20178 ( .A(n24910), .ZN(n26766) );
  INV_X1 U20179 ( .A(n24723), .ZN(n26767) );
  INV_X1 U20180 ( .A(n20713), .ZN(n26768) );
  INV_X1 U20181 ( .A(n24906), .ZN(n26769) );
  INV_X1 U20182 ( .A(n24907), .ZN(n267701) );
  INV_X1 U20183 ( .A(n24725), .ZN(n26771) );
  INV_X1 U20184 ( .A(n20711), .ZN(n26772) );
  INV_X1 U20185 ( .A(n24902), .ZN(n26773) );
  INV_X1 U20186 ( .A(n20712), .ZN(n26774) );
  INV_X1 U20187 ( .A(n24904), .ZN(n26775) );
  INV_X1 U20188 ( .A(n20709), .ZN(n26776) );
  INV_X1 U20189 ( .A(n24898), .ZN(n26777) );
  INV_X1 U20190 ( .A(n24900), .ZN(n26778) );
  INV_X1 U20191 ( .A(n24894), .ZN(n26779) );
  INV_X1 U20192 ( .A(n20708), .ZN(n267801) );
  INV_X1 U20193 ( .A(n24896), .ZN(n26781) );
  INV_X1 U20194 ( .A(n27204), .ZN(n26782) );
  INV_X1 U20195 ( .A(n24890), .ZN(n26783) );
  INV_X1 U20196 ( .A(n24890), .ZN(n26784) );
  INV_X1 U20197 ( .A(n24891), .ZN(n26785) );
  INV_X1 U20198 ( .A(n22492), .ZN(n26786) );
  INV_X1 U20199 ( .A(n20707), .ZN(n26787) );
  INV_X1 U20200 ( .A(n20707), .ZN(n26788) );
  INV_X1 U20201 ( .A(n24893), .ZN(n26789) );
  INV_X1 U20202 ( .A(n24886), .ZN(n267901) );
  INV_X1 U20203 ( .A(n24885), .ZN(n26791) );
  INV_X1 U20204 ( .A(n24885), .ZN(n26792) );
  INV_X1 U20205 ( .A(n23672), .ZN(n26793) );
  INV_X1 U20206 ( .A(n20706), .ZN(n26794) );
  INV_X1 U20207 ( .A(n20706), .ZN(n26795) );
  INV_X1 U20208 ( .A(n24888), .ZN(n26796) );
  INV_X1 U20209 ( .A(n3185), .ZN(n26797) );
  INV_X1 U20210 ( .A(n24880), .ZN(n26798) );
  INV_X1 U20211 ( .A(n20705), .ZN(n26799) );
  INV_X1 U20212 ( .A(n24883), .ZN(n268001) );
  INV_X1 U20213 ( .A(n24882), .ZN(n26801) );
  INV_X1 U20214 ( .A(n24882), .ZN(n26802) );
  INV_X1 U20215 ( .A(n38050), .ZN(n26803) );
  INV_X1 U20216 ( .A(n24875), .ZN(n26804) );
  INV_X1 U20217 ( .A(n20701), .ZN(n26805) );
  INV_X1 U20218 ( .A(n277401), .ZN(n26806) );
  INV_X1 U20219 ( .A(n20703), .ZN(n26807) );
  INV_X1 U20220 ( .A(n24877), .ZN(n26808) );
  INV_X1 U20221 ( .A(n24316), .ZN(n26809) );
  INV_X1 U20222 ( .A(n24315), .ZN(n268101) );
  INV_X1 U20223 ( .A(n24316), .ZN(n26811) );
  INV_X1 U20224 ( .A(n24315), .ZN(n26812) );
  INV_X1 U20225 ( .A(n24319), .ZN(n26813) );
  INV_X1 U20226 ( .A(n24318), .ZN(n26814) );
  INV_X1 U20227 ( .A(n24319), .ZN(n26815) );
  INV_X1 U20228 ( .A(n24318), .ZN(n26816) );
  INV_X1 U20229 ( .A(n24322), .ZN(n26817) );
  INV_X1 U20230 ( .A(n24321), .ZN(n26818) );
  INV_X1 U20231 ( .A(n24322), .ZN(n26819) );
  INV_X1 U20232 ( .A(n24321), .ZN(n268201) );
  INV_X1 U20233 ( .A(n24325), .ZN(n26821) );
  INV_X1 U20234 ( .A(n24324), .ZN(n26822) );
  INV_X1 U20235 ( .A(n24325), .ZN(n26823) );
  INV_X1 U20236 ( .A(n24324), .ZN(n26824) );
  INV_X1 U20237 ( .A(n24328), .ZN(n26825) );
  INV_X1 U20238 ( .A(n24327), .ZN(n26826) );
  INV_X1 U20239 ( .A(n24328), .ZN(n26827) );
  INV_X1 U20240 ( .A(n24327), .ZN(n26828) );
  INV_X1 U20241 ( .A(n24331), .ZN(n26829) );
  INV_X1 U20242 ( .A(n24330), .ZN(n268301) );
  INV_X1 U20243 ( .A(n24331), .ZN(n26831) );
  INV_X1 U20244 ( .A(n24330), .ZN(n26832) );
  INV_X1 U20245 ( .A(n24334), .ZN(n26833) );
  INV_X1 U20246 ( .A(n24333), .ZN(n26834) );
  INV_X1 U20247 ( .A(n24334), .ZN(n26835) );
  INV_X1 U20248 ( .A(n24333), .ZN(n26836) );
  INV_X1 U20249 ( .A(n24337), .ZN(n26837) );
  INV_X1 U20250 ( .A(n24336), .ZN(n26838) );
  INV_X1 U20251 ( .A(n24337), .ZN(n26839) );
  INV_X1 U20252 ( .A(n24336), .ZN(n268401) );
  INV_X1 U20253 ( .A(n24727), .ZN(n26841) );
  INV_X1 U20254 ( .A(n20698), .ZN(n26842) );
  INV_X1 U20255 ( .A(n20698), .ZN(n26843) );
  INV_X1 U20256 ( .A(n24870), .ZN(n26844) );
  INV_X1 U20257 ( .A(n24726), .ZN(n26845) );
  INV_X1 U20258 ( .A(n20699), .ZN(n26846) );
  INV_X1 U20259 ( .A(n20699), .ZN(n26847) );
  INV_X1 U20260 ( .A(n24872), .ZN(n26848) );
  INV_X1 U20261 ( .A(n20696), .ZN(n26849) );
  INV_X1 U20262 ( .A(n20696), .ZN(n268501) );
  INV_X1 U20263 ( .A(n24866), .ZN(n26851) );
  INV_X1 U20264 ( .A(n20697), .ZN(n26852) );
  INV_X1 U20265 ( .A(n20697), .ZN(n26853) );
  INV_X1 U20266 ( .A(n24868), .ZN(n26854) );
  INV_X1 U20267 ( .A(n20695), .ZN(n26855) );
  INV_X1 U20268 ( .A(n17104), .ZN(n26856) );
  INV_X1 U20269 ( .A(n20695), .ZN(n26857) );
  INV_X1 U20270 ( .A(n17104), .ZN(n26858) );
  INV_X1 U20271 ( .A(n24371), .ZN(n26859) );
  INV_X1 U20272 ( .A(n24370), .ZN(n268601) );
  INV_X1 U20273 ( .A(n24371), .ZN(n26861) );
  INV_X1 U20274 ( .A(n24373), .ZN(n26862) );
  INV_X1 U20275 ( .A(n24373), .ZN(n26863) );
  INV_X1 U20276 ( .A(n24372), .ZN(n26864) );
  INV_X1 U20277 ( .A(n24372), .ZN(n26865) );
  INV_X1 U20278 ( .A(n24648), .ZN(n26866) );
  INV_X1 U20279 ( .A(n24375), .ZN(n26867) );
  INV_X1 U20280 ( .A(n24377), .ZN(n26868) );
  INV_X1 U20281 ( .A(n24379), .ZN(n26869) );
  INV_X1 U20282 ( .A(n24379), .ZN(n268701) );
  INV_X1 U20283 ( .A(n24378), .ZN(n26871) );
  INV_X1 U20284 ( .A(n24378), .ZN(n26872) );
  INV_X1 U20285 ( .A(n24381), .ZN(n26873) );
  INV_X1 U20286 ( .A(n24380), .ZN(n26874) );
  INV_X1 U20287 ( .A(n24381), .ZN(n26875) );
  INV_X1 U20288 ( .A(n24380), .ZN(n26876) );
  INV_X1 U20289 ( .A(n24383), .ZN(n26877) );
  INV_X1 U20290 ( .A(n24383), .ZN(n26878) );
  INV_X1 U20291 ( .A(n24382), .ZN(n26879) );
  INV_X1 U20292 ( .A(n24382), .ZN(n268801) );
  INV_X1 U20293 ( .A(n24385), .ZN(n26881) );
  INV_X1 U20294 ( .A(n24384), .ZN(n26882) );
  INV_X1 U20295 ( .A(n24385), .ZN(n26883) );
  INV_X1 U20296 ( .A(n24384), .ZN(n26884) );
  INV_X1 U20297 ( .A(n24387), .ZN(n26885) );
  INV_X1 U20298 ( .A(n24387), .ZN(n26886) );
  INV_X1 U20299 ( .A(n24386), .ZN(n26887) );
  INV_X1 U20300 ( .A(n24386), .ZN(n26888) );
  INV_X1 U20301 ( .A(n24389), .ZN(n26889) );
  INV_X1 U20302 ( .A(n24388), .ZN(n268901) );
  INV_X1 U20303 ( .A(n24389), .ZN(n26891) );
  INV_X1 U20304 ( .A(n24388), .ZN(n26892) );
  INV_X1 U20305 ( .A(n24391), .ZN(n26893) );
  INV_X1 U20306 ( .A(n24391), .ZN(n26894) );
  INV_X1 U20307 ( .A(n24390), .ZN(n26895) );
  INV_X1 U20308 ( .A(n24390), .ZN(n26896) );
  INV_X1 U20309 ( .A(n24393), .ZN(n26897) );
  INV_X1 U20310 ( .A(n24392), .ZN(n26898) );
  INV_X1 U20311 ( .A(n24393), .ZN(n26899) );
  INV_X1 U20312 ( .A(n24392), .ZN(n269001) );
  INV_X1 U20313 ( .A(n20810), .ZN(n26901) );
  INV_X1 U20314 ( .A(n19067), .ZN(n26902) );
  INV_X1 U20315 ( .A(n277801), .ZN(n26903) );
  INV_X1 U20316 ( .A(n24863), .ZN(n26904) );
  INV_X1 U20317 ( .A(n278001), .ZN(n26905) );
  INV_X1 U20318 ( .A(n24407), .ZN(n26906) );
  INV_X1 U20319 ( .A(n24408), .ZN(n26907) );
  INV_X1 U20320 ( .A(n24408), .ZN(n26908) );
  INV_X1 U20321 ( .A(n24407), .ZN(n26909) );
  INV_X1 U20322 ( .A(n24410), .ZN(n269101) );
  INV_X1 U20323 ( .A(n24409), .ZN(n26911) );
  INV_X1 U20324 ( .A(n24410), .ZN(n26912) );
  INV_X1 U20325 ( .A(n24409), .ZN(n26913) );
  INV_X1 U20326 ( .A(n24412), .ZN(n26914) );
  INV_X1 U20327 ( .A(n24411), .ZN(n26915) );
  INV_X1 U20328 ( .A(n24412), .ZN(n26916) );
  INV_X1 U20329 ( .A(n24411), .ZN(n26917) );
  INV_X1 U20330 ( .A(n24413), .ZN(n26918) );
  INV_X1 U20331 ( .A(n24414), .ZN(n26919) );
  INV_X1 U20332 ( .A(n24413), .ZN(n269201) );
  INV_X1 U20333 ( .A(n24414), .ZN(n26921) );
  INV_X1 U20334 ( .A(n24416), .ZN(n26922) );
  INV_X1 U20335 ( .A(n24416), .ZN(n26923) );
  INV_X1 U20336 ( .A(n24419), .ZN(n26924) );
  INV_X1 U20337 ( .A(n24418), .ZN(n26925) );
  INV_X1 U20338 ( .A(n24418), .ZN(n26926) );
  INV_X1 U20339 ( .A(n20621), .ZN(n26927) );
  INV_X1 U20340 ( .A(n24818), .ZN(n26928) );
  INV_X1 U20341 ( .A(n20615), .ZN(n26929) );
  INV_X1 U20342 ( .A(n20616), .ZN(n269301) );
  INV_X1 U20343 ( .A(n20617), .ZN(n26931) );
  INV_X1 U20344 ( .A(n20617), .ZN(n26932) );
  INV_X1 U20345 ( .A(n24819), .ZN(n26933) );
  INV_X1 U20346 ( .A(n20612), .ZN(n26934) );
  INV_X1 U20347 ( .A(n20611), .ZN(n26935) );
  INV_X1 U20348 ( .A(n24815), .ZN(n26936) );
  INV_X1 U20349 ( .A(n20809), .ZN(n26937) );
  INV_X1 U20350 ( .A(n20809), .ZN(n26938) );
  INV_X1 U20351 ( .A(n3098), .ZN(n26939) );
  INV_X1 U20352 ( .A(n24813), .ZN(n269401) );
  INV_X1 U20353 ( .A(n24428), .ZN(n26941) );
  INV_X1 U20354 ( .A(n24429), .ZN(n26942) );
  INV_X1 U20355 ( .A(n24429), .ZN(n26943) );
  INV_X1 U20356 ( .A(n26976), .ZN(n26948) );
  INV_X1 U20357 ( .A(n24439), .ZN(n26962) );
  INV_X1 U20358 ( .A(n24702), .ZN(n26966) );
  BUF_X1 U20359 ( .A(add_124_aco_B_3_), .Z(n26967) );
  BUF_X1 U20360 ( .A(n26077), .Z(n26968) );
  NAND4_X1 U20361 ( .A1(N7942), .A2(n278201), .A3(n21519), .A4(n17114), .ZN(
        n4542) );
  INV_X1 U20362 ( .A(n20556), .ZN(n27201) );
  INV_X1 U20363 ( .A(n24485), .ZN(n27199) );
  INV_X1 U20364 ( .A(n20789), .ZN(n27766) );
  BUF_X1 U20365 ( .A(n25872), .Z(n27208) );
  BUF_X1 U20366 ( .A(n25872), .Z(n27207) );
  BUF_X1 U20367 ( .A(n25874), .Z(n27209) );
  BUF_X1 U20368 ( .A(n3987), .Z(n27153) );
  BUF_X1 U20369 ( .A(n3160), .Z(n27263) );
  BUF_X1 U20370 ( .A(n25936), .Z(n27155) );
  BUF_X1 U20371 ( .A(n25936), .Z(n27154) );
  BUF_X1 U20372 ( .A(n25935), .Z(n27265) );
  BUF_X1 U20373 ( .A(n25935), .Z(n27264) );
  BUF_X1 U20374 ( .A(n21368), .Z(n27148) );
  BUF_X1 U20375 ( .A(n21371), .Z(n27270) );
  BUF_X1 U20376 ( .A(n21369), .Z(n27150) );
  BUF_X1 U20377 ( .A(n21368), .Z(n27149) );
  BUF_X1 U20378 ( .A(n21372), .Z(n27272) );
  BUF_X1 U20379 ( .A(n21371), .Z(n27271) );
  INV_X1 U20380 ( .A(n24709), .ZN(n27188) );
  INV_X1 U20381 ( .A(n24703), .ZN(n27244) );
  INV_X1 U20382 ( .A(n24708), .ZN(n27197) );
  INV_X1 U20383 ( .A(n24511), .ZN(n27222) );
  BUF_X1 U20384 ( .A(n20481), .Z(n27027) );
  BUF_X1 U20385 ( .A(n25186), .Z(n27028) );
  BUF_X1 U20386 ( .A(n5305), .Z(n27029) );
  INV_X1 U20387 ( .A(n48840), .ZN(n27085) );
  INV_X1 U20388 ( .A(n48840), .ZN(n27086) );
  INV_X1 U20389 ( .A(n53060), .ZN(n27001) );
  INV_X1 U20390 ( .A(n53060), .ZN(n27002) );
  INV_X1 U20391 ( .A(n5304), .ZN(n27014) );
  INV_X1 U20392 ( .A(n5304), .ZN(n27015) );
  NAND2_X1 U20393 ( .A1(n25087), .A2(n19756), .ZN(n4818) );
  AND2_X1 U20394 ( .A1(n27811), .A2(n26529), .ZN(n3078) );
  AND2_X1 U20395 ( .A1(n27807), .A2(n26081), .ZN(n32600) );
  AND2_X1 U20396 ( .A1(n27817), .A2(n26527), .ZN(n38050) );
  AND2_X1 U20397 ( .A1(n27809), .A2(n26528), .ZN(n3185) );
  AND2_X1 U20398 ( .A1(n871), .A2(n22707), .ZN(n4543) );
  AND2_X1 U20399 ( .A1(n866), .A2(n27140), .ZN(n45180) );
  AND2_X1 U20400 ( .A1(n861), .A2(n21611), .ZN(n4494) );
  AND2_X1 U20401 ( .A1(n856), .A2(n26392), .ZN(n44700) );
  AND2_X1 U20402 ( .A1(n851), .A2(n21783), .ZN(n44450) );
  AND2_X1 U20403 ( .A1(n846), .A2(n21651), .ZN(n4421) );
  AND2_X1 U20404 ( .A1(n841), .A2(n25896), .ZN(n4396) );
  AND2_X1 U20405 ( .A1(n836), .A2(n21286), .ZN(n4371) );
  AND2_X1 U20406 ( .A1(n831), .A2(n27141), .ZN(n43470) );
  AND2_X1 U20407 ( .A1(n826), .A2(n24473), .ZN(n4324) );
  AND2_X1 U20408 ( .A1(n821), .A2(n26386), .ZN(n43020) );
  AND2_X1 U20409 ( .A1(n816), .A2(n21787), .ZN(n4280) );
  AND2_X1 U20410 ( .A1(n811), .A2(n21645), .ZN(n4258) );
  AND2_X1 U20411 ( .A1(n806), .A2(n25900), .ZN(n4236) );
  AND2_X1 U20412 ( .A1(n801), .A2(n21299), .ZN(n42140) );
  AND2_X1 U20413 ( .A1(n796), .A2(n25876), .ZN(n41880) );
  AND2_X1 U20414 ( .A1(n791), .A2(n21615), .ZN(n4164) );
  AND2_X1 U20415 ( .A1(n786), .A2(n25214), .ZN(n41410) );
  AND2_X1 U20416 ( .A1(n781), .A2(n21775), .ZN(n4119) );
  AND2_X1 U20417 ( .A1(n776), .A2(n24449), .ZN(n40970) );
  AND2_X1 U20418 ( .A1(n771), .A2(n24793), .ZN(n4075) );
  AND2_X1 U20419 ( .A1(n766), .A2(n256101), .ZN(n40530) );
  AND2_X1 U20420 ( .A1(n761), .A2(n25866), .ZN(n4031) );
  AND2_X1 U20421 ( .A1(n756), .A2(n21637), .ZN(n4005) );
  AND2_X1 U20422 ( .A1(n751), .A2(n26396), .ZN(n3981) );
  AND2_X1 U20423 ( .A1(n746), .A2(n21779), .ZN(n3958) );
  AND2_X1 U20424 ( .A1(n741), .A2(n20599), .ZN(n39360) );
  AND2_X1 U20425 ( .A1(n736), .A2(n21430), .ZN(n3914) );
  AND2_X1 U20426 ( .A1(n731), .A2(n21302), .ZN(n3892) );
  AND2_X1 U20427 ( .A1(n726), .A2(n20550), .ZN(n3870) );
  AND2_X1 U20428 ( .A1(n721), .A2(n21641), .ZN(n38480) );
  AND2_X1 U20429 ( .A1(n716), .A2(n21807), .ZN(n3823) );
  AND2_X1 U20430 ( .A1(n711), .A2(n24297), .ZN(n37990) );
  AND2_X1 U20431 ( .A1(n706), .A2(n20597), .ZN(n3776) );
  AND2_X1 U20432 ( .A1(n701), .A2(n24467), .ZN(n3754) );
  AND2_X1 U20433 ( .A1(n696), .A2(n17120), .ZN(n3732) );
  AND2_X1 U20434 ( .A1(n691), .A2(n24490), .ZN(n37100) );
  AND2_X1 U20435 ( .A1(n686), .A2(n24451), .ZN(n3688) );
  AND2_X1 U20436 ( .A1(n681), .A2(n21811), .ZN(n3666) );
  AND2_X1 U20437 ( .A1(n676), .A2(n26381), .ZN(n3642) );
  AND2_X1 U20438 ( .A1(n671), .A2(n21633), .ZN(n3618) );
  AND2_X1 U20439 ( .A1(n666), .A2(n25884), .ZN(n35950) );
  AND2_X1 U20440 ( .A1(n661), .A2(n24470), .ZN(n3573) );
  AND2_X1 U20441 ( .A1(n656), .A2(n24488), .ZN(n35510) );
  AND2_X1 U20442 ( .A1(n651), .A2(n20589), .ZN(n3529) );
  AND2_X1 U20443 ( .A1(n646), .A2(n21791), .ZN(n35070) );
  AND2_X1 U20444 ( .A1(n641), .A2(n25201), .ZN(n3485) );
  AND2_X1 U20445 ( .A1(n636), .A2(n21607), .ZN(n34600) );
  AND2_X1 U20446 ( .A1(n631), .A2(n25888), .ZN(n3436) );
  AND2_X1 U20447 ( .A1(n626), .A2(n22799), .ZN(n3413) );
  AND2_X1 U20448 ( .A1(n621), .A2(n25858), .ZN(n3391) );
  AND2_X1 U20449 ( .A1(n616), .A2(n20595), .ZN(n33690) );
  AND2_X1 U20450 ( .A1(n611), .A2(n21795), .ZN(n3347) );
  AND2_X1 U20451 ( .A1(n606), .A2(n25211), .ZN(n3325) );
  AND2_X1 U20452 ( .A1(n601), .A2(n24476), .ZN(n33030) );
  AND2_X1 U20453 ( .A1(n596), .A2(n27288), .ZN(n3278) );
  AND2_X1 U20454 ( .A1(n591), .A2(n21290), .ZN(n32540) );
  AND2_X1 U20455 ( .A1(n586), .A2(n25862), .ZN(n3229) );
  AND2_X1 U20456 ( .A1(n581), .A2(n21625), .ZN(n32040) );
  AND2_X1 U20457 ( .A1(n576), .A2(n24279), .ZN(n3179) );
  AND2_X1 U20458 ( .A1(n571), .A2(n26389), .ZN(n3154) );
  AND2_X1 U20459 ( .A1(n566), .A2(n21620), .ZN(n31290) );
  AND2_X1 U20460 ( .A1(n561), .A2(n27289), .ZN(n3104) );
  AND2_X1 U20461 ( .A1(n556), .A2(n22704), .ZN(n3072) );
  AND2_X1 U20462 ( .A1(n27816), .A2(n21519), .ZN(n3987) );
  AND2_X1 U20463 ( .A1(n27812), .A2(n26089), .ZN(n3160) );
  BUF_X1 U20464 ( .A(n4715), .Z(n26995) );
  AND2_X1 U20465 ( .A1(n27815), .A2(n21507), .ZN(n4170) );
  AND2_X1 U20466 ( .A1(n27813), .A2(n26082), .ZN(n3135) );
  BUF_X1 U20467 ( .A(n4716), .Z(n26996) );
  INV_X1 U20468 ( .A(n19215), .ZN(n27192) );
  INV_X1 U20469 ( .A(n21296), .ZN(n27191) );
  INV_X1 U20470 ( .A(n25263), .ZN(n27190) );
  INV_X1 U20471 ( .A(n21293), .ZN(n27189) );
  INV_X1 U20472 ( .A(n19219), .ZN(n27213) );
  INV_X1 U20473 ( .A(n21308), .ZN(n27212) );
  INV_X1 U20474 ( .A(n25272), .ZN(n27211) );
  INV_X1 U20475 ( .A(n21305), .ZN(n27210) );
  INV_X1 U20476 ( .A(n19221), .ZN(n27195) );
  INV_X1 U20477 ( .A(n21314), .ZN(n27194) );
  INV_X1 U20478 ( .A(n21311), .ZN(n27193) );
  INV_X1 U20479 ( .A(n19223), .ZN(n27216) );
  INV_X1 U20480 ( .A(n21320), .ZN(n27215) );
  INV_X1 U20481 ( .A(n21317), .ZN(n27214) );
  INV_X1 U20482 ( .A(n24700), .ZN(n27219) );
  INV_X1 U20483 ( .A(n20511), .ZN(n27177) );
  INV_X1 U20484 ( .A(n24731), .ZN(n27178) );
  INV_X1 U20485 ( .A(n20507), .ZN(n27232) );
  INV_X1 U20486 ( .A(n24730), .ZN(n27233) );
  INV_X1 U20487 ( .A(n25101), .ZN(n27186) );
  INV_X1 U20488 ( .A(n25102), .ZN(n27185) );
  INV_X1 U20489 ( .A(n19026), .ZN(n27184) );
  INV_X1 U20490 ( .A(n25102), .ZN(n27183) );
  INV_X1 U20491 ( .A(n19022), .ZN(n27182) );
  INV_X1 U20492 ( .A(n25096), .ZN(n27181) );
  INV_X1 U20493 ( .A(n25095), .ZN(n27180) );
  INV_X1 U20494 ( .A(n25096), .ZN(n27179) );
  INV_X1 U20495 ( .A(n25097), .ZN(n27241) );
  INV_X1 U20496 ( .A(n25098), .ZN(n27240) );
  INV_X1 U20497 ( .A(n19023), .ZN(n27239) );
  INV_X1 U20498 ( .A(n25098), .ZN(n27238) );
  INV_X1 U20499 ( .A(n19020), .ZN(n27237) );
  INV_X1 U20500 ( .A(n25091), .ZN(n27236) );
  INV_X1 U20501 ( .A(n24618), .ZN(n27242) );
  INV_X1 U20502 ( .A(n25090), .ZN(n27235) );
  INV_X1 U20503 ( .A(n25091), .ZN(n27234) );
  BUF_X1 U20504 ( .A(n17990), .Z(n27047) );
  INV_X1 U20505 ( .A(n24614), .ZN(n27161) );
  INV_X1 U20506 ( .A(n24629), .ZN(n27249) );
  INV_X1 U20507 ( .A(n24609), .ZN(n27165) );
  INV_X1 U20508 ( .A(n24611), .ZN(n27164) );
  INV_X1 U20509 ( .A(n24612), .ZN(n27162) );
  INV_X1 U20510 ( .A(n24624), .ZN(n27253) );
  INV_X1 U20511 ( .A(n24626), .ZN(n27252) );
  INV_X1 U20512 ( .A(n24627), .ZN(n27250) );
  NAND2_X1 U20513 ( .A1(n26986), .A2(n26555), .ZN(n4989) );
  AND2_X1 U20514 ( .A1(n22421), .A2(n22954), .ZN(n48840) );
  AND2_X1 U20515 ( .A1(n24706), .A2(n26374), .ZN(n53060) );
  AND2_X1 U20516 ( .A1(n24705), .A2(n25754), .ZN(n5304) );
  INV_X1 U20517 ( .A(n24606), .ZN(n27170) );
  INV_X1 U20518 ( .A(n24606), .ZN(n27168) );
  INV_X1 U20519 ( .A(n24609), .ZN(n27167) );
  INV_X1 U20520 ( .A(n24621), .ZN(n27258) );
  INV_X1 U20521 ( .A(n24621), .ZN(n27256) );
  INV_X1 U20522 ( .A(n24624), .ZN(n27255) );
  AND2_X1 U20523 ( .A1(n24706), .A2(n26147), .ZN(n5305) );
  INV_X1 U20524 ( .A(n24701), .ZN(n27073) );
  INV_X1 U20525 ( .A(n4889), .ZN(n27048) );
  INV_X1 U20526 ( .A(n24702), .ZN(n27074) );
  INV_X1 U20527 ( .A(n20493), .ZN(n27099) );
  INV_X1 U20528 ( .A(n24701), .ZN(n27075) );
  INV_X1 U20529 ( .A(n20488), .ZN(n27062) );
  INV_X1 U20530 ( .A(n4889), .ZN(n27049) );
  INV_X1 U20531 ( .A(n5206), .ZN(n27030) );
  INV_X1 U20532 ( .A(n5206), .ZN(n27031) );
  INV_X1 U20533 ( .A(n44660), .ZN(n27817) );
  INV_X1 U20534 ( .A(n43920), .ZN(n27807) );
  INV_X1 U20535 ( .A(n3481), .ZN(n27813) );
  INV_X1 U20536 ( .A(n3097), .ZN(n27811) );
  INV_X1 U20537 ( .A(n4026), .ZN(n27808) );
  NAND2_X1 U20538 ( .A1(n20895), .A2(n21508), .ZN(n4819) );
  INV_X1 U20539 ( .A(n20498), .ZN(n27796) );
  INV_X1 U20540 ( .A(n20496), .ZN(n27804) );
  AND2_X1 U20541 ( .A1(n26083), .A2(n17266), .ZN(n45490) );
  NOR2_X1 U20542 ( .A1(n27767), .A2(n23732), .ZN(n4979) );
  INV_X1 U20543 ( .A(n3988), .ZN(n27797) );
  INV_X1 U20544 ( .A(n3161), .ZN(n27803) );
  BUF_X1 U20545 ( .A(n21860), .Z(n27172) );
  BUF_X1 U20546 ( .A(n26319), .Z(n27174) );
  BUF_X1 U20547 ( .A(n21859), .Z(n27173) );
  BUF_X1 U20548 ( .A(n21863), .Z(n27226) );
  BUF_X1 U20549 ( .A(n21862), .Z(n27225) );
  BUF_X1 U20550 ( .A(n26320), .Z(n27228) );
  BUF_X1 U20551 ( .A(n21861), .Z(n27227) );
  INV_X1 U20552 ( .A(n24693), .ZN(n27795) );
  INV_X1 U20553 ( .A(n24695), .ZN(n27805) );
  BUF_X1 U20554 ( .A(n21864), .Z(n27229) );
  BUF_X1 U20555 ( .A(n21337), .Z(n27157) );
  BUF_X1 U20556 ( .A(n19229), .Z(n27156) );
  BUF_X1 U20557 ( .A(n21326), .Z(n27245) );
  BUF_X1 U20558 ( .A(n19226), .Z(n27246) );
  BUF_X1 U20559 ( .A(n21338), .Z(n27158) );
  NOR2_X1 U20560 ( .A1(n22734), .A2(n26938), .ZN(n4715) );
  NOR2_X1 U20561 ( .A1(n22739), .A2(n24426), .ZN(n4716) );
  AND2_X1 U20562 ( .A1(n25631), .A2(n21632), .ZN(n5205) );
  AND2_X1 U20563 ( .A1(n22425), .A2(n26084), .ZN(n27098) );
  AND2_X1 U20564 ( .A1(n22421), .A2(n26085), .ZN(n4885) );
  AND2_X1 U20565 ( .A1(n26501), .A2(n21875), .ZN(n27061) );
  AND2_X1 U20566 ( .A1(n22424), .A2(n21876), .ZN(n4890) );
  BUF_X1 U20567 ( .A(n17268), .Z(n26988) );
  BUF_X1 U20568 ( .A(n4987), .Z(n27044) );
  BUF_X1 U20569 ( .A(n4982), .Z(n27045) );
  BUF_X1 U20570 ( .A(n4983), .Z(n27046) );
  BUF_X1 U20571 ( .A(n24693), .Z(n27125) );
  BUF_X1 U20572 ( .A(n24695), .Z(n27273) );
  BUF_X1 U20573 ( .A(n43460), .Z(n27126) );
  BUF_X1 U20574 ( .A(n3103), .Z(n27274) );
  BUF_X1 U20575 ( .A(n20900), .Z(n27127) );
  BUF_X1 U20576 ( .A(n20905), .Z(n27275) );
  NAND2_X1 U20577 ( .A1(n21872), .A2(n23685), .ZN(n4990) );
  BUF_X1 U20578 ( .A(n25661), .Z(n27152) );
  BUF_X1 U20579 ( .A(n21402), .Z(n27151) );
  BUF_X1 U20580 ( .A(n21397), .Z(n27261) );
  BUF_X1 U20581 ( .A(n21398), .Z(n27262) );
  BUF_X1 U20582 ( .A(n25945), .Z(n27145) );
  BUF_X1 U20583 ( .A(n25953), .Z(n27266) );
  BUF_X1 U20584 ( .A(n25948), .Z(n27146) );
  BUF_X1 U20585 ( .A(n25956), .Z(n27268) );
  BUF_X1 U20586 ( .A(n25953), .Z(n27267) );
  NAND2_X1 U20587 ( .A1(n25949), .A2(n265501), .ZN(n4985) );
  NAND2_X1 U20588 ( .A1(n23679), .A2(n25312), .ZN(n4986) );
  BUF_X1 U20589 ( .A(n25948), .Z(n27147) );
  BUF_X1 U20590 ( .A(n25956), .Z(n27269) );
  INV_X1 U20591 ( .A(n37980), .ZN(n27160) );
  INV_X1 U20592 ( .A(n37980), .ZN(n27159) );
  INV_X1 U20593 ( .A(n20902), .ZN(n27176) );
  INV_X1 U20594 ( .A(n20903), .ZN(n27175) );
  INV_X1 U20595 ( .A(n20907), .ZN(n27231) );
  INV_X1 U20596 ( .A(n20908), .ZN(n27230) );
  INV_X1 U20597 ( .A(n31780), .ZN(n27248) );
  INV_X1 U20598 ( .A(n31780), .ZN(n27247) );
  AND2_X1 U20599 ( .A1(n22424), .A2(n25937), .ZN(n4889) );
  AND2_X1 U20600 ( .A1(n20896), .A2(n26326), .ZN(n47890) );
  AND2_X1 U20601 ( .A1(n25087), .A2(n25941), .ZN(n47880) );
  AND2_X1 U20602 ( .A1(n21330), .A2(n26373), .ZN(n5206) );
  BUF_X1 U20603 ( .A(n26968), .Z(n26989) );
  BUF_X1 U20604 ( .A(n26968), .Z(n26990) );
  NAND3_X1 U20605 ( .A1(n25508), .A2(n25518), .A3(n24690), .ZN(n44660) );
  NAND3_X1 U20606 ( .A1(n24720), .A2(n17121), .A3(n4028), .ZN(n43920) );
  NAND3_X1 U20607 ( .A1(n24721), .A2(n17121), .A3(n24689), .ZN(n3481) );
  BUF_X1 U20608 ( .A(n26997), .Z(n26998) );
  NAND2_X1 U20609 ( .A1(n24690), .A2(n24691), .ZN(n3097) );
  BUF_X1 U20610 ( .A(n20888), .Z(n26999) );
  NAND2_X1 U20611 ( .A1(n17997), .A2(n24691), .ZN(n4026) );
  INV_X1 U20612 ( .A(n4491), .ZN(n27816) );
  INV_X1 U20613 ( .A(n44420), .ZN(n27818) );
  INV_X1 U20614 ( .A(n4539), .ZN(n27814) );
  INV_X1 U20615 ( .A(n4417), .ZN(n27819) );
  INV_X1 U20616 ( .A(n45150), .ZN(n27815) );
  INV_X1 U20617 ( .A(n3663), .ZN(n27812) );
  INV_X1 U20618 ( .A(n32990), .ZN(n278101) );
  INV_X1 U20619 ( .A(n38440), .ZN(n27809) );
  AOI211_X1 U20620 ( .C1(n22448), .C2(N7942), .A(n24073), .B(n17266), .ZN(
        n4567) );
  NOR3_X1 U20621 ( .A1(n22727), .A2(n19266), .A3(n27811), .ZN(n3099) );
  AND2_X1 U20622 ( .A1(n25746), .A2(n26677), .ZN(n4713) );
  AND2_X1 U20623 ( .A1(n25758), .A2(n20746), .ZN(n4714) );
  NOR2_X1 U20624 ( .A1(alu_start), .A2(n25001), .ZN(n3098) );
  AOI211_X1 U20625 ( .C1(n26505), .C2(r929_LT_LE), .A(n27807), .B(n22728), 
        .ZN(n43930) );
  INV_X1 U20626 ( .A(n19754), .ZN(n27792) );
  INV_X1 U20627 ( .A(n45660), .ZN(n278201) );
  NOR2_X1 U20628 ( .A1(n25927), .A2(n44670), .ZN(n38060) );
  AOI211_X1 U20629 ( .C1(n22432), .C2(N5213), .A(n27817), .B(n25002), .ZN(
        n44670) );
  NOR2_X1 U20630 ( .A1(n25289), .A2(n38450), .ZN(n3186) );
  AOI211_X1 U20631 ( .C1(n22434), .C2(N2903), .A(n27809), .B(n24071), .ZN(
        n38450) );
  NOR2_X1 U20632 ( .A1(n20609), .A2(n44430), .ZN(n36250) );
  AOI211_X1 U20633 ( .C1(n21866), .C2(N4509), .A(n27818), .B(n26653), .ZN(
        n44430) );
  NOR2_X1 U20634 ( .A1(n22530), .A2(n4027), .ZN(n32110) );
  AOI211_X1 U20635 ( .C1(n26514), .C2(N2985), .A(n27808), .B(n24073), .ZN(
        n4027) );
  NOR2_X1 U20636 ( .A1(n25316), .A2(n4418), .ZN(n3443) );
  AOI211_X1 U20637 ( .C1(n17073), .C2(r948_LT_LE), .A(n27819), .B(n22728), 
        .ZN(n4418) );
  NOR2_X1 U20638 ( .A1(n25282), .A2(n42100), .ZN(n3236) );
  AOI211_X1 U20639 ( .C1(n26322), .C2(r924_LT_LE), .A(n20798), .B(n17265), 
        .ZN(n42100) );
  NOR2_X1 U20640 ( .A1(n21279), .A2(n4492), .ZN(n3988) );
  AOI211_X1 U20641 ( .C1(n22447), .C2(N5888), .A(n27816), .B(n24074), .ZN(
        n4492) );
  NOR2_X1 U20642 ( .A1(n21323), .A2(n3664), .ZN(n3161) );
  AOI211_X1 U20643 ( .C1(n21867), .C2(N2811), .A(n27812), .B(n25002), .ZN(
        n3664) );
  INV_X1 U20644 ( .A(n24714), .ZN(n27791) );
  NOR2_X1 U20645 ( .A1(n22744), .A2(n21491), .ZN(n4987) );
  AOI211_X1 U20646 ( .C1(n26506), .C2(N7267), .A(n27814), .B(n24074), .ZN(
        n4540) );
  AOI211_X1 U20647 ( .C1(n26505), .C2(N2637), .A(n278101), .B(n20798), .ZN(
        n33000) );
  INV_X1 U20648 ( .A(n42090), .ZN(n27806) );
  AND3_X1 U20649 ( .A1(n18431), .A2(n5200), .A3(n21331), .ZN(n27043) );
  NOR2_X1 U20650 ( .A1(n22727), .A2(n26941), .ZN(n30950) );
  BUF_X1 U20651 ( .A(n25377), .Z(n27112) );
  BUF_X1 U20652 ( .A(n25377), .Z(n27111) );
  AOI211_X1 U20653 ( .C1(n22448), .C2(N2729), .A(n27813), .B(n26652), .ZN(
        n3482) );
  AOI211_X1 U20654 ( .C1(n26322), .C2(N6563), .A(n27815), .B(n26653), .ZN(
        n45160) );
  NOR2_X1 U20655 ( .A1(n24712), .A2(n21504), .ZN(n4982) );
  NOR2_X1 U20656 ( .A1(n24715), .A2(n21465), .ZN(n4983) );
  AND4_X1 U20657 ( .A1(N5888), .A2(n22468), .A3(n19266), .A4(n4491), .ZN(
        n39800) );
  INV_X1 U20658 ( .A(n20752), .ZN(n27782) );
  AND4_X1 U20659 ( .A1(N2729), .A2(n260901), .A3(n21868), .A4(n3481), .ZN(
        n31280) );
  AND4_X1 U20660 ( .A1(N6563), .A2(n21517), .A3(n26506), .A4(n45150), .ZN(
        n4163) );
  NAND3_X1 U20661 ( .A1(n27794), .A2(n25663), .A3(n24686), .ZN(n26987) );
  AND4_X1 U20662 ( .A1(N5213), .A2(n22472), .A3(n17073), .A4(n44660), .ZN(
        n37980) );
  AND4_X1 U20663 ( .A1(N2903), .A2(n26089), .A3(n21866), .A4(n38440), .ZN(
        n31780) );
  AND4_X1 U20664 ( .A1(N2637), .A2(n265301), .A3(n26515), .A4(n32990), .ZN(
        n3103) );
  AND4_X1 U20665 ( .A1(N7267), .A2(n21506), .A3(n22447), .A4(n4539), .ZN(
        n43460) );
  INV_X1 U20666 ( .A(n53950), .ZN(n27741) );
  OAI22_X1 U20667 ( .A1(n24684), .A2(n22951), .B1(n24675), .B2(n24678), .ZN(
        n4419) );
  INV_X1 U20668 ( .A(n17102), .ZN(n27726) );
  BUF_X1 U20669 ( .A(n26675), .Z(n26991) );
  INV_X1 U20670 ( .A(n24711), .ZN(n27789) );
  OAI22_X1 U20671 ( .A1(n22950), .A2(n24677), .B1(n24676), .B2(n24683), .ZN(
        n3483) );
  BUF_X1 U20672 ( .A(n25649), .Z(n26992) );
  OAI22_X1 U20673 ( .A1(n24683), .A2(n42110), .B1(n24677), .B2(n42120), .ZN(
        n42090) );
  OAI22_X1 U20674 ( .A1(n24678), .A2(n42110), .B1(n24684), .B2(n42120), .ZN(
        n45660) );
  OAI21_X1 U20675 ( .B1(n17085), .B2(n18514), .A(n17996), .ZN(n44680) );
  NAND3_X1 U20676 ( .A1(n24676), .A2(n19178), .A3(n24681), .ZN(n42120) );
  BUF_X1 U20677 ( .A(n25645), .Z(n26993) );
  NAND3_X1 U20678 ( .A1(n25509), .A2(n25518), .A3(n24687), .ZN(n4491) );
  BUF_X1 U20679 ( .A(n19237), .Z(n26994) );
  NAND2_X1 U20680 ( .A1(n17085), .A2(n27302), .ZN(n4569) );
  NAND3_X1 U20681 ( .A1(n25512), .A2(n19174), .A3(n24687), .ZN(n44420) );
  NAND3_X1 U20682 ( .A1(n25512), .A2(n25509), .A3(n17997), .ZN(n4539) );
  NAND3_X1 U20683 ( .A1(n25511), .A2(n25508), .A3(n24689), .ZN(n4417) );
  NAND3_X1 U20684 ( .A1(n19175), .A2(n19174), .A3(n24681), .ZN(n45150) );
  NAND3_X1 U20685 ( .A1(n24720), .A2(n19178), .A3(n24688), .ZN(n3663) );
  NAND3_X1 U20686 ( .A1(n22950), .A2(n25510), .A3(n24682), .ZN(n42110) );
  NAND2_X1 U20687 ( .A1(n5299), .A2(n25957), .ZN(n26997) );
  NAND2_X1 U20688 ( .A1(n24688), .A2(n24692), .ZN(n32990) );
  AND2_X1 U20689 ( .A1(n24717), .A2(n22953), .ZN(n4028) );
  INV_X1 U20690 ( .A(n19756), .ZN(n26977) );
  NAND2_X1 U20691 ( .A1(n24682), .A2(n24692), .ZN(n38440) );
  INV_X1 U20692 ( .A(n20885), .ZN(n27304) );
  INV_X1 U20693 ( .A(n27295), .ZN(n27306) );
  INV_X1 U20694 ( .A(n27294), .ZN(n27305) );
  NAND3_X1 U20695 ( .A1(n880), .A2(n885), .A3(n17083), .ZN(n47050) );
  NAND3_X1 U20696 ( .A1(n884), .A2(n24686), .A3(n878), .ZN(n51360) );
  NAND3_X1 U20697 ( .A1(n882), .A2(n25665), .A3(n19109), .ZN(n47060) );
  NAND2_X1 U20698 ( .A1(n5293), .A2(n5294), .ZN(mul_outcome[126]) );
  AOI221_X1 U20699 ( .B1(n24397), .B2(matrix_mul_2D_6__5__0_), .C1(n24313), 
        .C2(matrix_mul_2D_6__7__0_), .A(n5298), .ZN(n5293) );
  NAND2_X1 U20700 ( .A1(n5289), .A2(n5290), .ZN(mul_outcome[127]) );
  AOI221_X1 U20701 ( .B1(n25027), .B2(matrix_mul_2D_6__5__1_), .C1(n17116), 
        .C2(matrix_mul_2D_6__7__1_), .A(n5292), .ZN(n5289) );
  NAND2_X1 U20702 ( .A1(n5285), .A2(n5286), .ZN(mul_outcome[128]) );
  AOI221_X1 U20703 ( .B1(n24425), .B2(matrix_mul_2D_6__5__2_), .C1(n22427), 
        .C2(matrix_mul_2D_6__7__2_), .A(n5288), .ZN(n5285) );
  NAND2_X1 U20704 ( .A1(n5281), .A2(n5282), .ZN(mul_outcome[129]) );
  AOI221_X1 U20705 ( .B1(n24427), .B2(matrix_mul_2D_6__5__3_), .C1(n24310), 
        .C2(matrix_mul_2D_6__7__3_), .A(n5284), .ZN(n5281) );
  NAND2_X1 U20706 ( .A1(n5273), .A2(n5274), .ZN(mul_outcome[130]) );
  AOI221_X1 U20707 ( .B1(n25029), .B2(matrix_mul_2D_6__5__4_), .C1(n26498), 
        .C2(matrix_mul_2D_6__7__4_), .A(n5276), .ZN(n5273) );
  NAND2_X1 U20708 ( .A1(n52690), .A2(n52700), .ZN(mul_outcome[131]) );
  AOI221_X1 U20709 ( .B1(n24395), .B2(matrix_mul_2D_6__5__5_), .C1(n23378), 
        .C2(matrix_mul_2D_6__7__5_), .A(n5272), .ZN(n52690) );
  NAND2_X1 U20710 ( .A1(n52650), .A2(n52660), .ZN(mul_outcome[132]) );
  AOI221_X1 U20711 ( .B1(n24817), .B2(matrix_mul_2D_6__5__6_), .C1(n22419), 
        .C2(matrix_mul_2D_6__7__6_), .A(n52680), .ZN(n52650) );
  NAND2_X1 U20712 ( .A1(n52610), .A2(n52620), .ZN(mul_outcome[133]) );
  AOI221_X1 U20713 ( .B1(n21971), .B2(matrix_mul_2D_6__5__7_), .C1(n26240), 
        .C2(matrix_mul_2D_6__7__7_), .A(n52640), .ZN(n52610) );
  NAND2_X1 U20714 ( .A1(n52570), .A2(n52580), .ZN(mul_outcome[134]) );
  AOI221_X1 U20715 ( .B1(n20614), .B2(matrix_mul_2D_6__5__8_), .C1(n19311), 
        .C2(matrix_mul_2D_6__7__8_), .A(n52600), .ZN(n52570) );
  NAND2_X1 U20716 ( .A1(n52530), .A2(n52540), .ZN(mul_outcome[135]) );
  AOI221_X1 U20717 ( .B1(n24399), .B2(matrix_mul_2D_6__5__9_), .C1(n26503), 
        .C2(matrix_mul_2D_6__7__9_), .A(n52560), .ZN(n52530) );
  NAND2_X1 U20718 ( .A1(n5249), .A2(n52500), .ZN(mul_outcome[136]) );
  AOI221_X1 U20719 ( .B1(n25033), .B2(matrix_mul_2D_6__5__10_), .C1(n26244), 
        .C2(matrix_mul_2D_6__7__10_), .A(n52520), .ZN(n5249) );
  NAND2_X1 U20720 ( .A1(n5245), .A2(n5246), .ZN(mul_outcome[137]) );
  AOI221_X1 U20721 ( .B1(n21976), .B2(matrix_mul_2D_6__5__11_), .C1(n26504), 
        .C2(matrix_mul_2D_6__7__11_), .A(n5248), .ZN(n5245) );
  NAND2_X1 U20722 ( .A1(n5241), .A2(n5242), .ZN(mul_outcome[138]) );
  AOI221_X1 U20723 ( .B1(n25029), .B2(matrix_mul_2D_6__5__12_), .C1(n26243), 
        .C2(matrix_mul_2D_6__7__12_), .A(n5244), .ZN(n5241) );
  NAND2_X1 U20724 ( .A1(n5237), .A2(n5238), .ZN(mul_outcome[139]) );
  AOI221_X1 U20725 ( .B1(n26937), .B2(matrix_mul_2D_6__5__13_), .C1(n26497), 
        .C2(matrix_mul_2D_6__7__13_), .A(n5240), .ZN(n5237) );
  NAND2_X1 U20726 ( .A1(n52290), .A2(n52300), .ZN(mul_outcome[140]) );
  AOI221_X1 U20727 ( .B1(n20811), .B2(matrix_mul_2D_6__5__14_), .C1(n22430), 
        .C2(matrix_mul_2D_6__7__14_), .A(n52320), .ZN(n52290) );
  NAND2_X1 U20728 ( .A1(n5197), .A2(n5198), .ZN(mul_outcome[147]) );
  AOI221_X1 U20729 ( .B1(n22431), .B2(matrix_mul_2D_7__6__0_), .C1(n24942), 
        .C2(matrix_mul_2D_7__7__0_), .A(n5202), .ZN(n5197) );
  NAND2_X1 U20730 ( .A1(n5193), .A2(n5194), .ZN(mul_outcome[148]) );
  AOI221_X1 U20731 ( .B1(n22428), .B2(matrix_mul_2D_7__6__1_), .C1(n25330), 
        .C2(matrix_mul_2D_7__7__1_), .A(n5196), .ZN(n5193) );
  NAND2_X1 U20732 ( .A1(n5189), .A2(n5190), .ZN(mul_outcome[149]) );
  AOI221_X1 U20733 ( .B1(n26502), .B2(matrix_mul_2D_7__6__2_), .C1(n24159), 
        .C2(matrix_mul_2D_7__7__2_), .A(n5192), .ZN(n5189) );
  NAND2_X1 U20734 ( .A1(n51810), .A2(n51820), .ZN(mul_outcome[150]) );
  AOI221_X1 U20735 ( .B1(n22420), .B2(matrix_mul_2D_7__6__3_), .C1(n24942), 
        .C2(matrix_mul_2D_7__7__3_), .A(n51840), .ZN(n51810) );
  NAND2_X1 U20736 ( .A1(n51770), .A2(n51780), .ZN(mul_outcome[151]) );
  AOI221_X1 U20737 ( .B1(n22431), .B2(matrix_mul_2D_7__6__4_), .C1(n24157), 
        .C2(matrix_mul_2D_7__7__4_), .A(n51800), .ZN(n51770) );
  NAND2_X1 U20738 ( .A1(n51730), .A2(n51740), .ZN(mul_outcome[152]) );
  AOI221_X1 U20739 ( .B1(n26496), .B2(matrix_mul_2D_7__6__5_), .C1(n25331), 
        .C2(matrix_mul_2D_7__7__5_), .A(n51760), .ZN(n51730) );
  NAND2_X1 U20740 ( .A1(n51690), .A2(n51700), .ZN(mul_outcome[153]) );
  AOI221_X1 U20741 ( .B1(n26808), .B2(matrix_mul_2D_7__6__6_), .C1(n25331), 
        .C2(matrix_mul_2D_7__7__6_), .A(n51720), .ZN(n51690) );
  NAND2_X1 U20742 ( .A1(n5165), .A2(n5166), .ZN(mul_outcome[154]) );
  AOI221_X1 U20743 ( .B1(n24312), .B2(matrix_mul_2D_7__6__7_), .C1(n19299), 
        .C2(matrix_mul_2D_7__7__7_), .A(n51680), .ZN(n5165) );
  NAND2_X1 U20744 ( .A1(n5161), .A2(n5162), .ZN(mul_outcome[155]) );
  AOI221_X1 U20745 ( .B1(n24309), .B2(matrix_mul_2D_7__6__8_), .C1(n19086), 
        .C2(matrix_mul_2D_7__7__8_), .A(n5164), .ZN(n5161) );
  NAND2_X1 U20746 ( .A1(n5157), .A2(n5158), .ZN(mul_outcome[156]) );
  AOI221_X1 U20747 ( .B1(n26244), .B2(matrix_mul_2D_7__6__9_), .C1(n24941), 
        .C2(matrix_mul_2D_7__7__9_), .A(n5160), .ZN(n5157) );
  NAND2_X1 U20748 ( .A1(n5153), .A2(n5154), .ZN(mul_outcome[157]) );
  AOI221_X1 U20749 ( .B1(n23377), .B2(matrix_mul_2D_7__6__10_), .C1(n24938), 
        .C2(matrix_mul_2D_7__7__10_), .A(n5156), .ZN(n5153) );
  NAND2_X1 U20750 ( .A1(n51490), .A2(n51500), .ZN(mul_outcome[158]) );
  AOI221_X1 U20751 ( .B1(n26498), .B2(matrix_mul_2D_7__6__11_), .C1(n24939), 
        .C2(matrix_mul_2D_7__7__11_), .A(n5152), .ZN(n51490) );
  NAND2_X1 U20752 ( .A1(n51450), .A2(n51460), .ZN(mul_outcome[159]) );
  AOI221_X1 U20753 ( .B1(n26807), .B2(matrix_mul_2D_7__6__12_), .C1(n26707), 
        .C2(matrix_mul_2D_7__7__12_), .A(n51480), .ZN(n51450) );
  NAND2_X1 U20754 ( .A1(n51370), .A2(n51380), .ZN(mul_outcome[160]) );
  AOI221_X1 U20755 ( .B1(n26504), .B2(matrix_mul_2D_7__6__13_), .C1(n24160), 
        .C2(matrix_mul_2D_7__7__13_), .A(n51400), .ZN(n51370) );
  NAND2_X1 U20756 ( .A1(n5130), .A2(n5131), .ZN(mul_outcome[161]) );
  AOI221_X1 U20757 ( .B1(n24313), .B2(matrix_mul_2D_7__6__14_), .C1(n24160), 
        .C2(matrix_mul_2D_7__7__14_), .A(n5134), .ZN(n5130) );
  NAND3_X1 U20758 ( .A1(n49750), .A2(n49760), .A3(n4977), .ZN(mul_outcome[42])
         );
  AOI22_X1 U20759 ( .A1(n27059), .A2(matrix_mul_2D_2__2__0_), .B1(n25635), 
        .B2(matrix_mul_2D_2__3__0_), .ZN(n49750) );
  NAND3_X1 U20760 ( .A1(n49710), .A2(n49720), .A3(n49730), .ZN(mul_outcome[43]) );
  AOI22_X1 U20761 ( .A1(n27050), .A2(matrix_mul_2D_2__2__1_), .B1(n25636), 
        .B2(matrix_mul_2D_2__3__1_), .ZN(n49710) );
  NAND3_X1 U20762 ( .A1(n49670), .A2(n49680), .A3(n49690), .ZN(mul_outcome[44]) );
  AOI22_X1 U20763 ( .A1(n27051), .A2(matrix_mul_2D_2__2__2_), .B1(n19228), 
        .B2(matrix_mul_2D_2__3__2_), .ZN(n49670) );
  NAND3_X1 U20764 ( .A1(n49630), .A2(n49640), .A3(n49650), .ZN(mul_outcome[45]) );
  AOI22_X1 U20765 ( .A1(n27052), .A2(matrix_mul_2D_2__2__3_), .B1(n25635), 
        .B2(matrix_mul_2D_2__3__3_), .ZN(n49630) );
  NAND3_X1 U20766 ( .A1(n4959), .A2(n4960), .A3(n49610), .ZN(mul_outcome[46])
         );
  AOI22_X1 U20767 ( .A1(n27053), .A2(matrix_mul_2D_2__2__4_), .B1(n25636), 
        .B2(matrix_mul_2D_2__3__4_), .ZN(n4959) );
  NAND3_X1 U20768 ( .A1(n4955), .A2(n4956), .A3(n4957), .ZN(mul_outcome[47])
         );
  AOI22_X1 U20769 ( .A1(n27054), .A2(matrix_mul_2D_2__2__5_), .B1(n25632), 
        .B2(matrix_mul_2D_2__3__5_), .ZN(n4955) );
  NAND3_X1 U20770 ( .A1(n4951), .A2(n4952), .A3(n4953), .ZN(mul_outcome[48])
         );
  AOI22_X1 U20771 ( .A1(n27055), .A2(matrix_mul_2D_2__2__6_), .B1(n21340), 
        .B2(matrix_mul_2D_2__3__6_), .ZN(n4951) );
  NAND3_X1 U20772 ( .A1(n4947), .A2(n4948), .A3(n4949), .ZN(mul_outcome[49])
         );
  AOI22_X1 U20773 ( .A1(n27056), .A2(matrix_mul_2D_2__2__7_), .B1(n21344), 
        .B2(matrix_mul_2D_2__3__7_), .ZN(n4947) );
  NAND3_X1 U20774 ( .A1(n4939), .A2(n4940), .A3(n4941), .ZN(mul_outcome[50])
         );
  AOI22_X1 U20775 ( .A1(n27057), .A2(matrix_mul_2D_2__2__8_), .B1(n25632), 
        .B2(matrix_mul_2D_2__3__8_), .ZN(n4939) );
  NAND3_X1 U20776 ( .A1(n4935), .A2(n4936), .A3(n4937), .ZN(mul_outcome[51])
         );
  AOI22_X1 U20777 ( .A1(n27055), .A2(matrix_mul_2D_2__2__9_), .B1(n21341), 
        .B2(matrix_mul_2D_2__3__9_), .ZN(n4935) );
  NAND3_X1 U20778 ( .A1(n4931), .A2(n4932), .A3(n4933), .ZN(mul_outcome[52])
         );
  AOI22_X1 U20779 ( .A1(n27056), .A2(matrix_mul_2D_2__2__10_), .B1(n21345), 
        .B2(matrix_mul_2D_2__3__10_), .ZN(n4931) );
  NAND3_X1 U20780 ( .A1(n4927), .A2(n4928), .A3(n4929), .ZN(mul_outcome[53])
         );
  AOI22_X1 U20781 ( .A1(n27057), .A2(matrix_mul_2D_2__2__11_), .B1(n21333), 
        .B2(matrix_mul_2D_2__3__11_), .ZN(n4927) );
  NAND3_X1 U20782 ( .A1(n4923), .A2(n4924), .A3(n4925), .ZN(mul_outcome[54])
         );
  AOI22_X1 U20783 ( .A1(n27058), .A2(matrix_mul_2D_2__2__12_), .B1(n19230), 
        .B2(matrix_mul_2D_2__3__12_), .ZN(n4923) );
  NAND3_X1 U20784 ( .A1(n49190), .A2(n49200), .A3(n49210), .ZN(mul_outcome[55]) );
  AOI22_X1 U20785 ( .A1(n27059), .A2(matrix_mul_2D_2__2__13_), .B1(n21345), 
        .B2(matrix_mul_2D_2__3__13_), .ZN(n49190) );
  NAND3_X1 U20786 ( .A1(n49150), .A2(n49160), .A3(n49170), .ZN(mul_outcome[56]) );
  AOI22_X1 U20787 ( .A1(n27060), .A2(matrix_mul_2D_2__2__14_), .B1(n21334), 
        .B2(matrix_mul_2D_2__3__14_), .ZN(n49150) );
  NAND3_X1 U20788 ( .A1(n4779), .A2(n4780), .A3(n4781), .ZN(mul_outcome[84])
         );
  AOI221_X1 U20789 ( .B1(n21062), .B2(matrix_mul_2D_4__6__0_), .C1(n24817), 
        .C2(matrix_mul_2D_4__7__0_), .A(n4782), .ZN(n4781) );
  NAND3_X1 U20790 ( .A1(n4775), .A2(n4776), .A3(n4777), .ZN(mul_outcome[85])
         );
  AOI221_X1 U20791 ( .B1(n21000), .B2(matrix_mul_2D_4__6__1_), .C1(n25027), 
        .C2(matrix_mul_2D_4__7__1_), .A(n4778), .ZN(n4777) );
  NAND3_X1 U20792 ( .A1(n4771), .A2(n4772), .A3(n4773), .ZN(mul_outcome[86])
         );
  AOI221_X1 U20793 ( .B1(n19312), .B2(matrix_mul_2D_4__6__2_), .C1(n24425), 
        .C2(matrix_mul_2D_4__7__2_), .A(n4774), .ZN(n4773) );
  NAND3_X1 U20794 ( .A1(n4767), .A2(n4768), .A3(n4769), .ZN(mul_outcome[87])
         );
  AOI221_X1 U20795 ( .B1(n26622), .B2(matrix_mul_2D_4__6__3_), .C1(n24427), 
        .C2(matrix_mul_2D_4__7__3_), .A(n4770), .ZN(n4769) );
  NAND3_X1 U20796 ( .A1(n4763), .A2(n4764), .A3(n4765), .ZN(mul_outcome[88])
         );
  AOI221_X1 U20797 ( .B1(n23973), .B2(matrix_mul_2D_4__6__4_), .C1(n24398), 
        .C2(matrix_mul_2D_4__7__4_), .A(n4766), .ZN(n4765) );
  NAND3_X1 U20798 ( .A1(n4759), .A2(n4760), .A3(n4761), .ZN(mul_outcome[89])
         );
  AOI221_X1 U20799 ( .B1(n23981), .B2(matrix_mul_2D_4__6__5_), .C1(n25033), 
        .C2(matrix_mul_2D_4__7__5_), .A(n4762), .ZN(n4761) );
  NAND3_X1 U20800 ( .A1(n4751), .A2(n4752), .A3(n4753), .ZN(mul_outcome[90])
         );
  AOI221_X1 U20801 ( .B1(n26620), .B2(matrix_mul_2D_4__6__6_), .C1(n24402), 
        .C2(matrix_mul_2D_4__7__6_), .A(n4754), .ZN(n4753) );
  NAND3_X1 U20802 ( .A1(n47470), .A2(n47480), .A3(n4749), .ZN(mul_outcome[91])
         );
  AOI221_X1 U20803 ( .B1(n23970), .B2(matrix_mul_2D_4__6__7_), .C1(n21975), 
        .C2(matrix_mul_2D_4__7__7_), .A(n4750), .ZN(n4749) );
  NAND3_X1 U20804 ( .A1(n47430), .A2(n47440), .A3(n47450), .ZN(mul_outcome[92]) );
  AOI221_X1 U20805 ( .B1(n26927), .B2(matrix_mul_2D_4__6__8_), .C1(n24424), 
        .C2(matrix_mul_2D_4__7__8_), .A(n47460), .ZN(n47450) );
  NAND3_X1 U20806 ( .A1(n47390), .A2(n47400), .A3(n47410), .ZN(mul_outcome[93]) );
  AOI221_X1 U20807 ( .B1(n23658), .B2(matrix_mul_2D_4__6__9_), .C1(n20814), 
        .C2(matrix_mul_2D_4__7__9_), .A(n47420), .ZN(n47410) );
  NAND3_X1 U20808 ( .A1(n47350), .A2(n47360), .A3(n47370), .ZN(mul_outcome[94]) );
  AOI221_X1 U20809 ( .B1(n23978), .B2(matrix_mul_2D_4__6__10_), .C1(n20810), 
        .C2(matrix_mul_2D_4__7__10_), .A(n47380), .ZN(n47370) );
  NAND3_X1 U20810 ( .A1(n47310), .A2(n47320), .A3(n47330), .ZN(mul_outcome[95]) );
  AOI221_X1 U20811 ( .B1(n22676), .B2(matrix_mul_2D_4__6__11_), .C1(n26938), 
        .C2(matrix_mul_2D_4__7__11_), .A(n47340), .ZN(n47330) );
  NAND3_X1 U20812 ( .A1(n4727), .A2(n47280), .A3(n47290), .ZN(mul_outcome[96])
         );
  AOI221_X1 U20813 ( .B1(n19273), .B2(matrix_mul_2D_4__6__12_), .C1(n23493), 
        .C2(matrix_mul_2D_4__7__12_), .A(n47300), .ZN(n47290) );
  NAND3_X1 U20814 ( .A1(n4723), .A2(n4724), .A3(n4725), .ZN(mul_outcome[97])
         );
  AOI221_X1 U20815 ( .B1(n19274), .B2(matrix_mul_2D_4__6__13_), .C1(n20613), 
        .C2(matrix_mul_2D_4__7__13_), .A(n4726), .ZN(n4725) );
  NAND3_X1 U20816 ( .A1(n4717), .A2(n4718), .A3(n4719), .ZN(mul_outcome[98])
         );
  AOI221_X1 U20817 ( .B1(n25024), .B2(matrix_mul_2D_4__6__14_), .C1(n21970), 
        .C2(matrix_mul_2D_4__7__14_), .A(n4720), .ZN(n4719) );
  NAND3_X1 U20818 ( .A1(n48760), .A2(n48770), .A3(n48780), .ZN(mul_outcome[63]) );
  AOI22_X1 U20819 ( .A1(n21185), .A2(matrix_mul_2D_3__2__0_), .B1(n23726), 
        .B2(matrix_mul_2D_3__6__0_), .ZN(n48760) );
  NAND3_X1 U20820 ( .A1(n48720), .A2(n48730), .A3(n48740), .ZN(mul_outcome[64]) );
  AOI22_X1 U20821 ( .A1(n25759), .A2(matrix_mul_2D_3__2__1_), .B1(n24856), 
        .B2(matrix_mul_2D_3__6__1_), .ZN(n48720) );
  NAND3_X1 U20822 ( .A1(n4868), .A2(n48690), .A3(n48700), .ZN(mul_outcome[65])
         );
  AOI22_X1 U20823 ( .A1(n25756), .A2(matrix_mul_2D_3__2__2_), .B1(n20861), 
        .B2(matrix_mul_2D_3__6__2_), .ZN(n4868) );
  NAND3_X1 U20824 ( .A1(n4864), .A2(n4865), .A3(n4866), .ZN(mul_outcome[66])
         );
  AOI22_X1 U20825 ( .A1(n25757), .A2(matrix_mul_2D_3__2__3_), .B1(n26589), 
        .B2(matrix_mul_2D_3__6__3_), .ZN(n4864) );
  NAND3_X1 U20826 ( .A1(n4860), .A2(n4861), .A3(n4862), .ZN(mul_outcome[67])
         );
  AOI22_X1 U20827 ( .A1(n21186), .A2(matrix_mul_2D_3__2__4_), .B1(n20687), 
        .B2(matrix_mul_2D_3__6__4_), .ZN(n4860) );
  NAND3_X1 U20828 ( .A1(n4856), .A2(n4857), .A3(n4858), .ZN(mul_outcome[68])
         );
  AOI22_X1 U20829 ( .A1(n25761), .A2(matrix_mul_2D_3__2__5_), .B1(n21146), 
        .B2(matrix_mul_2D_3__6__5_), .ZN(n4856) );
  NAND3_X1 U20830 ( .A1(n4852), .A2(n4853), .A3(n4854), .ZN(mul_outcome[69])
         );
  AOI22_X1 U20831 ( .A1(n25758), .A2(matrix_mul_2D_3__2__6_), .B1(n23733), 
        .B2(matrix_mul_2D_3__6__6_), .ZN(n4852) );
  NAND3_X1 U20832 ( .A1(n4844), .A2(n4845), .A3(n4846), .ZN(mul_outcome[70])
         );
  AOI22_X1 U20833 ( .A1(n25757), .A2(matrix_mul_2D_3__2__7_), .B1(n22535), 
        .B2(matrix_mul_2D_3__6__7_), .ZN(n4844) );
  NAND3_X1 U20834 ( .A1(n48400), .A2(n4841), .A3(n4842), .ZN(mul_outcome[71])
         );
  AOI22_X1 U20835 ( .A1(n25539), .A2(matrix_mul_2D_3__2__8_), .B1(n22538), 
        .B2(matrix_mul_2D_3__6__8_), .ZN(n48400) );
  NAND3_X1 U20836 ( .A1(n48360), .A2(n48370), .A3(n48380), .ZN(mul_outcome[72]) );
  AOI22_X1 U20837 ( .A1(n19185), .A2(matrix_mul_2D_3__2__9_), .B1(n20692), 
        .B2(matrix_mul_2D_3__6__9_), .ZN(n48360) );
  NAND3_X1 U20838 ( .A1(n48320), .A2(n48330), .A3(n48340), .ZN(mul_outcome[73]) );
  AOI22_X1 U20839 ( .A1(n25760), .A2(matrix_mul_2D_3__2__10_), .B1(n20693), 
        .B2(matrix_mul_2D_3__6__10_), .ZN(n48320) );
  NAND3_X1 U20840 ( .A1(n48280), .A2(n48290), .A3(n48300), .ZN(mul_outcome[74]) );
  AOI22_X1 U20841 ( .A1(n25755), .A2(matrix_mul_2D_3__2__11_), .B1(n22533), 
        .B2(matrix_mul_2D_3__6__11_), .ZN(n48280) );
  NAND3_X1 U20842 ( .A1(n48240), .A2(n48250), .A3(n48260), .ZN(mul_outcome[75]) );
  AOI22_X1 U20843 ( .A1(n25754), .A2(matrix_mul_2D_3__2__12_), .B1(n23729), 
        .B2(matrix_mul_2D_3__6__12_), .ZN(n48240) );
  NAND3_X1 U20844 ( .A1(n48200), .A2(n48210), .A3(n48220), .ZN(mul_outcome[76]) );
  AOI22_X1 U20845 ( .A1(n25539), .A2(matrix_mul_2D_3__2__13_), .B1(n24859), 
        .B2(matrix_mul_2D_3__6__13_), .ZN(n48200) );
  NAND3_X1 U20846 ( .A1(n4814), .A2(n4815), .A3(n4816), .ZN(mul_outcome[77])
         );
  AOI22_X1 U20847 ( .A1(n25761), .A2(matrix_mul_2D_3__2__14_), .B1(n26588), 
        .B2(matrix_mul_2D_3__6__14_), .ZN(n4814) );
  NAND2_X1 U20848 ( .A1(n5075), .A2(n50760), .ZN(mul_outcome[21]) );
  AOI221_X1 U20849 ( .B1(n26341), .B2(matrix_mul_2D_1__6__0_), .C1(n26762), 
        .C2(matrix_mul_2D_1__7__0_), .A(n50800), .ZN(n5075) );
  NAND2_X1 U20850 ( .A1(n5071), .A2(n5072), .ZN(mul_outcome[22]) );
  AOI221_X1 U20851 ( .B1(n26339), .B2(matrix_mul_2D_1__6__1_), .C1(n21833), 
        .C2(matrix_mul_2D_1__7__1_), .A(n5074), .ZN(n5071) );
  NAND2_X1 U20852 ( .A1(n5067), .A2(n5068), .ZN(mul_outcome[23]) );
  AOI221_X1 U20853 ( .B1(n26106), .B2(matrix_mul_2D_1__6__2_), .C1(n21434), 
        .C2(matrix_mul_2D_1__7__2_), .A(n5070), .ZN(n5067) );
  NAND2_X1 U20854 ( .A1(n5063), .A2(n5064), .ZN(mul_outcome[24]) );
  AOI221_X1 U20855 ( .B1(n21548), .B2(matrix_mul_2D_1__6__3_), .C1(n24259), 
        .C2(matrix_mul_2D_1__7__3_), .A(n5066), .ZN(n5063) );
  NAND2_X1 U20856 ( .A1(n5059), .A2(n5060), .ZN(mul_outcome[25]) );
  AOI221_X1 U20857 ( .B1(n26340), .B2(matrix_mul_2D_1__6__4_), .C1(n21831), 
        .C2(matrix_mul_2D_1__7__4_), .A(n5062), .ZN(n5059) );
  NAND2_X1 U20858 ( .A1(n50550), .A2(n50560), .ZN(mul_outcome[26]) );
  AOI221_X1 U20859 ( .B1(n21893), .B2(matrix_mul_2D_1__6__5_), .C1(n19247), 
        .C2(matrix_mul_2D_1__7__5_), .A(n50580), .ZN(n50550) );
  NAND2_X1 U20860 ( .A1(n50510), .A2(n50520), .ZN(mul_outcome[27]) );
  AOI221_X1 U20861 ( .B1(n26106), .B2(matrix_mul_2D_1__6__6_), .C1(n24262), 
        .C2(matrix_mul_2D_1__7__6_), .A(n50540), .ZN(n50510) );
  NAND2_X1 U20862 ( .A1(n50470), .A2(n50480), .ZN(mul_outcome[28]) );
  AOI221_X1 U20863 ( .B1(n21549), .B2(matrix_mul_2D_1__6__7_), .C1(n25916), 
        .C2(matrix_mul_2D_1__7__7_), .A(n50500), .ZN(n50470) );
  NAND2_X1 U20864 ( .A1(n50430), .A2(n50440), .ZN(mul_outcome[29]) );
  AOI221_X1 U20865 ( .B1(n21892), .B2(matrix_mul_2D_1__6__8_), .C1(n21489), 
        .C2(matrix_mul_2D_1__7__8_), .A(n50460), .ZN(n50430) );
  NAND2_X1 U20866 ( .A1(n5035), .A2(n5036), .ZN(mul_outcome[30]) );
  AOI221_X1 U20867 ( .B1(n21895), .B2(matrix_mul_2D_1__6__9_), .C1(n21462), 
        .C2(matrix_mul_2D_1__7__9_), .A(n5038), .ZN(n5035) );
  NAND2_X1 U20868 ( .A1(n5031), .A2(n5032), .ZN(mul_outcome[31]) );
  AOI221_X1 U20869 ( .B1(n21547), .B2(matrix_mul_2D_1__6__10_), .C1(n21504), 
        .C2(matrix_mul_2D_1__7__10_), .A(n5034), .ZN(n5031) );
  NAND2_X1 U20870 ( .A1(n5027), .A2(n5028), .ZN(mul_outcome[32]) );
  AOI221_X1 U20871 ( .B1(n26105), .B2(matrix_mul_2D_1__6__11_), .C1(n21491), 
        .C2(matrix_mul_2D_1__7__11_), .A(n5030), .ZN(n5027) );
  NAND2_X1 U20872 ( .A1(n5023), .A2(n5024), .ZN(mul_outcome[33]) );
  AOI221_X1 U20873 ( .B1(n21896), .B2(matrix_mul_2D_1__6__12_), .C1(n260601), 
        .C2(matrix_mul_2D_1__7__12_), .A(n5026), .ZN(n5023) );
  NAND2_X1 U20874 ( .A1(n5019), .A2(n5020), .ZN(mul_outcome[34]) );
  AOI221_X1 U20875 ( .B1(n26341), .B2(matrix_mul_2D_1__6__13_), .C1(n21499), 
        .C2(matrix_mul_2D_1__7__13_), .A(n5022), .ZN(n5019) );
  NAND2_X1 U20876 ( .A1(n5015), .A2(n5016), .ZN(mul_outcome[35]) );
  AOI221_X1 U20877 ( .B1(n21550), .B2(matrix_mul_2D_1__6__14_), .C1(n26074), 
        .C2(matrix_mul_2D_1__7__14_), .A(n5018), .ZN(n5015) );
  NAND3_X1 U20878 ( .A1(n54180), .A2(n54190), .A3(n54200), .ZN(mul_outcome[0])
         );
  AOI22_X1 U20879 ( .A1(n26979), .A2(matrix_mul_2D_0__6__0_), .B1(n24156), 
        .B2(matrix_mul_2D_0__1__0_), .ZN(n54180) );
  NAND3_X1 U20880 ( .A1(n50850), .A2(n50860), .A3(n50870), .ZN(mul_outcome[1])
         );
  AOI22_X1 U20881 ( .A1(n26983), .A2(matrix_mul_2D_0__6__1_), .B1(n24156), 
        .B2(matrix_mul_2D_0__1__1_), .ZN(n50850) );
  NAND3_X1 U20882 ( .A1(n5039), .A2(n5040), .A3(n5041), .ZN(mul_outcome[2]) );
  AOI22_X1 U20883 ( .A1(n26978), .A2(matrix_mul_2D_0__6__2_), .B1(n19085), 
        .B2(matrix_mul_2D_0__1__2_), .ZN(n5039) );
  NAND3_X1 U20884 ( .A1(n49950), .A2(n49960), .A3(n49970), .ZN(mul_outcome[3])
         );
  AOI22_X1 U20885 ( .A1(n22957), .A2(matrix_mul_2D_0__6__3_), .B1(n24155), 
        .B2(matrix_mul_2D_0__1__3_), .ZN(n49950) );
  NAND3_X1 U20886 ( .A1(n4943), .A2(n4944), .A3(n4945), .ZN(mul_outcome[4]) );
  AOI22_X1 U20887 ( .A1(n26985), .A2(matrix_mul_2D_0__6__4_), .B1(n24153), 
        .B2(matrix_mul_2D_0__1__4_), .ZN(n4943) );
  NAND3_X1 U20888 ( .A1(n4899), .A2(n4900), .A3(n4901), .ZN(mul_outcome[5]) );
  AOI22_X1 U20889 ( .A1(n22954), .A2(matrix_mul_2D_0__6__5_), .B1(n26704), 
        .B2(matrix_mul_2D_0__1__5_), .ZN(n4899) );
  NAND3_X1 U20890 ( .A1(n4848), .A2(n4849), .A3(n4850), .ZN(mul_outcome[6]) );
  AOI22_X1 U20891 ( .A1(n22958), .A2(matrix_mul_2D_0__6__6_), .B1(n24153), 
        .B2(matrix_mul_2D_0__1__6_), .ZN(n4848) );
  NAND3_X1 U20892 ( .A1(n48020), .A2(n4803), .A3(n4804), .ZN(mul_outcome[7])
         );
  AOI22_X1 U20893 ( .A1(n26985), .A2(matrix_mul_2D_0__6__7_), .B1(n24150), 
        .B2(matrix_mul_2D_0__1__7_), .ZN(n48020) );
  NAND3_X1 U20894 ( .A1(n4755), .A2(n4756), .A3(n4757), .ZN(mul_outcome[8]) );
  AOI22_X1 U20895 ( .A1(n22957), .A2(matrix_mul_2D_0__6__8_), .B1(n25328), 
        .B2(matrix_mul_2D_0__1__8_), .ZN(n4755) );
  NAND3_X1 U20896 ( .A1(n47000), .A2(n47010), .A3(n47020), .ZN(mul_outcome[9])
         );
  AOI22_X1 U20897 ( .A1(n26986), .A2(matrix_mul_2D_0__6__9_), .B1(n24152), 
        .B2(matrix_mul_2D_0__1__9_), .ZN(n47000) );
  NAND3_X1 U20898 ( .A1(n5371), .A2(n5372), .A3(n5373), .ZN(mul_outcome[10])
         );
  AOI22_X1 U20899 ( .A1(n26980), .A2(matrix_mul_2D_0__6__10_), .B1(n24944), 
        .B2(matrix_mul_2D_0__1__10_), .ZN(n5371) );
  NAND3_X1 U20900 ( .A1(n5327), .A2(n5328), .A3(n5329), .ZN(mul_outcome[11])
         );
  AOI22_X1 U20901 ( .A1(n26981), .A2(matrix_mul_2D_0__6__11_), .B1(n24945), 
        .B2(matrix_mul_2D_0__1__11_), .ZN(n5327) );
  NAND3_X1 U20902 ( .A1(n5277), .A2(n5278), .A3(n5279), .ZN(mul_outcome[12])
         );
  AOI22_X1 U20903 ( .A1(n26982), .A2(matrix_mul_2D_0__6__12_), .B1(n25329), 
        .B2(matrix_mul_2D_0__1__12_), .ZN(n5277) );
  NAND3_X1 U20904 ( .A1(n5233), .A2(n5234), .A3(n5235), .ZN(mul_outcome[13])
         );
  AOI22_X1 U20905 ( .A1(n26983), .A2(matrix_mul_2D_0__6__13_), .B1(n25329), 
        .B2(matrix_mul_2D_0__1__13_), .ZN(n5233) );
  NAND3_X1 U20906 ( .A1(n51850), .A2(n51860), .A3(n51870), .ZN(mul_outcome[14]) );
  AOI22_X1 U20907 ( .A1(n26984), .A2(matrix_mul_2D_0__6__14_), .B1(n19298), 
        .B2(matrix_mul_2D_0__1__14_), .ZN(n51850) );
  NAND3_X1 U20908 ( .A1(n53910), .A2(n53920), .A3(n53930), .ZN(
        mul_outcome[105]) );
  AOI221_X1 U20909 ( .B1(n24396), .B2(matrix_mul_2D_5__6__0_), .C1(n25910), 
        .C2(matrix_mul_2D_5__7__0_), .A(n53940), .ZN(n53930) );
  NAND3_X1 U20910 ( .A1(n53870), .A2(n53880), .A3(n53890), .ZN(
        mul_outcome[106]) );
  AOI221_X1 U20911 ( .B1(n26404), .B2(matrix_mul_2D_5__6__1_), .C1(n21502), 
        .C2(matrix_mul_2D_5__7__1_), .A(n53900), .ZN(n53890) );
  NAND3_X1 U20912 ( .A1(n5383), .A2(n5384), .A3(n53850), .ZN(mul_outcome[107])
         );
  AOI221_X1 U20913 ( .B1(n26403), .B2(matrix_mul_2D_5__6__2_), .C1(n19249), 
        .C2(matrix_mul_2D_5__7__2_), .A(n53860), .ZN(n53850) );
  NAND3_X1 U20914 ( .A1(n5379), .A2(n5380), .A3(n5381), .ZN(mul_outcome[108])
         );
  AOI221_X1 U20915 ( .B1(n24426), .B2(matrix_mul_2D_5__6__3_), .C1(n21495), 
        .C2(matrix_mul_2D_5__7__3_), .A(n5382), .ZN(n5381) );
  NAND3_X1 U20916 ( .A1(n5375), .A2(n5376), .A3(n5377), .ZN(mul_outcome[109])
         );
  AOI221_X1 U20917 ( .B1(n26401), .B2(matrix_mul_2D_5__6__4_), .C1(n26068), 
        .C2(matrix_mul_2D_5__7__4_), .A(n5378), .ZN(n5377) );
  NAND3_X1 U20918 ( .A1(n5367), .A2(n5368), .A3(n5369), .ZN(mul_outcome[110])
         );
  AOI221_X1 U20919 ( .B1(n24401), .B2(matrix_mul_2D_5__6__5_), .C1(n21436), 
        .C2(matrix_mul_2D_5__7__5_), .A(n5370), .ZN(n5369) );
  NAND3_X1 U20920 ( .A1(n5363), .A2(n5364), .A3(n5365), .ZN(mul_outcome[111])
         );
  AOI221_X1 U20921 ( .B1(n20815), .B2(matrix_mul_2D_5__6__6_), .C1(n26076), 
        .C2(matrix_mul_2D_5__7__6_), .A(n5366), .ZN(n5365) );
  NAND3_X1 U20922 ( .A1(n53590), .A2(n5360), .A3(n5361), .ZN(mul_outcome[112])
         );
  AOI221_X1 U20923 ( .B1(n26400), .B2(matrix_mul_2D_5__6__7_), .C1(n26067), 
        .C2(matrix_mul_2D_5__7__7_), .A(n5362), .ZN(n5361) );
  NAND3_X1 U20924 ( .A1(n53550), .A2(n53560), .A3(n53570), .ZN(
        mul_outcome[113]) );
  AOI221_X1 U20925 ( .B1(n24400), .B2(matrix_mul_2D_5__6__8_), .C1(n26758), 
        .C2(matrix_mul_2D_5__7__8_), .A(n53580), .ZN(n53570) );
  NAND3_X1 U20926 ( .A1(n53510), .A2(n53520), .A3(n53530), .ZN(
        mul_outcome[114]) );
  AOI221_X1 U20927 ( .B1(n21972), .B2(matrix_mul_2D_5__6__9_), .C1(n17077), 
        .C2(matrix_mul_2D_5__7__9_), .A(n53540), .ZN(n53530) );
  NAND3_X1 U20928 ( .A1(n53470), .A2(n53480), .A3(n53490), .ZN(
        mul_outcome[115]) );
  AOI221_X1 U20929 ( .B1(n25026), .B2(matrix_mul_2D_5__6__10_), .C1(n25908), 
        .C2(matrix_mul_2D_5__7__10_), .A(n53500), .ZN(n53490) );
  NAND3_X1 U20930 ( .A1(n53430), .A2(n53440), .A3(n53450), .ZN(
        mul_outcome[116]) );
  AOI221_X1 U20931 ( .B1(n19272), .B2(matrix_mul_2D_5__6__11_), .C1(n22830), 
        .C2(matrix_mul_2D_5__7__11_), .A(n53460), .ZN(n53450) );
  NAND3_X1 U20932 ( .A1(n53390), .A2(n53400), .A3(n53410), .ZN(
        mul_outcome[117]) );
  AOI221_X1 U20933 ( .B1(n21967), .B2(matrix_mul_2D_5__6__12_), .C1(n26066), 
        .C2(matrix_mul_2D_5__7__12_), .A(n53420), .ZN(n53410) );
  NAND3_X1 U20934 ( .A1(n5335), .A2(n5336), .A3(n5337), .ZN(mul_outcome[118])
         );
  AOI221_X1 U20935 ( .B1(n23492), .B2(matrix_mul_2D_5__6__13_), .C1(n26756), 
        .C2(matrix_mul_2D_5__7__13_), .A(n5338), .ZN(n5337) );
  NAND3_X1 U20936 ( .A1(n5331), .A2(n5332), .A3(n5333), .ZN(mul_outcome[119])
         );
  AOI221_X1 U20937 ( .B1(n26395), .B2(matrix_mul_2D_5__6__14_), .C1(n26075), 
        .C2(matrix_mul_2D_5__7__14_), .A(n5334), .ZN(n5333) );
  NOR3_X1 U20938 ( .A1(n462), .A2(n545), .A3(n536), .ZN(add_124_aco_B_3_) );
  NAND3_X1 U20939 ( .A1(n883), .A2(n20891), .A3(n878), .ZN(n54230) );
  NAND4_X1 U20940 ( .A1(n457), .A2(n880), .A3(n27741), .A4(n21438), .ZN(n5200)
         );
  INV_X1 U20941 ( .A(n883), .ZN(n27794) );
  NAND3_X1 U20942 ( .A1(n24685), .A2(n17080), .A3(n879), .ZN(n5133) );
  NAND3_X1 U20943 ( .A1(n24685), .A2(n25662), .A3(n882), .ZN(n4721) );
  INV_X1 U20944 ( .A(n877), .ZN(n277901) );
  NAND3_X1 U20945 ( .A1(n17086), .A2(n17080), .A3(n879), .ZN(n50780) );
  NAND2_X1 U20946 ( .A1(srstn), .A2(n23961), .ZN(n4571) );
  NAND3_X1 U20947 ( .A1(n47980), .A2(n47990), .A3(n48000), .ZN(mul_outcome[80]) );
  AOI22_X1 U20948 ( .A1(n19185), .A2(n17721), .B1(n24858), .B2(n17673), .ZN(
        n47980) );
  AOI22_X1 U20949 ( .A1(n27102), .A2(n17745), .B1(n19184), .B2(n17733), .ZN(
        n47990) );
  AOI221_X1 U20950 ( .B1(n26762), .B2(n17685), .C1(n23971), .C2(n17661), .A(
        n27763), .ZN(n48000) );
  NAND3_X1 U20951 ( .A1(n4810), .A2(n4811), .A3(n4812), .ZN(mul_outcome[78])
         );
  AOI22_X1 U20952 ( .A1(n25760), .A2(n17725), .B1(n25065), .B2(n17677), .ZN(
        n4810) );
  AOI22_X1 U20953 ( .A1(n27100), .A2(n17749), .B1(n25536), .B2(n17737), .ZN(
        n4811) );
  AOI221_X1 U20954 ( .B1(n26306), .B2(n17689), .C1(n23982), .C2(n17665), .A(
        n27765), .ZN(n4812) );
  AOI221_X1 U20955 ( .B1(n26305), .B2(matrix_mul_2D_3__5__0_), .C1(n23979), 
        .C2(matrix_mul_2D_3__7__0_), .A(n48790), .ZN(n48780) );
  OAI22_X1 U20956 ( .A1(n2306), .A2(n24090), .B1(n2321), .B2(n24094), .ZN(
        n48790) );
  AOI221_X1 U20957 ( .B1(n22838), .B2(matrix_mul_2D_3__5__1_), .C1(n19102), 
        .C2(matrix_mul_2D_3__7__1_), .A(n48750), .ZN(n48740) );
  OAI22_X1 U20958 ( .A1(n2305), .A2(n24091), .B1(n2320), .B2(n24095), .ZN(
        n48750) );
  AOI221_X1 U20959 ( .B1(n25917), .B2(matrix_mul_2D_3__5__2_), .C1(n22879), 
        .C2(matrix_mul_2D_3__7__2_), .A(n48710), .ZN(n48700) );
  OAI22_X1 U20960 ( .A1(n2304), .A2(n24991), .B1(n2319), .B2(n24994), .ZN(
        n48710) );
  AOI221_X1 U20961 ( .B1(n24258), .B2(matrix_mul_2D_3__5__3_), .C1(n23974), 
        .C2(matrix_mul_2D_3__7__3_), .A(n4867), .ZN(n4866) );
  OAI22_X1 U20962 ( .A1(n2303), .A2(n20790), .B1(n2318), .B2(n20791), .ZN(
        n4867) );
  AOI221_X1 U20963 ( .B1(n26055), .B2(matrix_mul_2D_3__5__4_), .C1(n22678), 
        .C2(matrix_mul_2D_3__7__4_), .A(n4863), .ZN(n4862) );
  OAI22_X1 U20964 ( .A1(n2302), .A2(n26664), .B1(n2317), .B2(n26667), .ZN(
        n4863) );
  AOI221_X1 U20965 ( .B1(n26755), .B2(matrix_mul_2D_3__5__5_), .C1(n23982), 
        .C2(matrix_mul_2D_3__7__5_), .A(n4859), .ZN(n4858) );
  OAI22_X1 U20966 ( .A1(n2301), .A2(n26665), .B1(n2316), .B2(n24092), .ZN(
        n4859) );
  AOI221_X1 U20967 ( .B1(n24261), .B2(matrix_mul_2D_3__5__6_), .C1(n23971), 
        .C2(matrix_mul_2D_3__7__6_), .A(n4855), .ZN(n4854) );
  OAI22_X1 U20968 ( .A1(n2300), .A2(n26665), .B1(n2315), .B2(n19291), .ZN(
        n4855) );
  AOI221_X1 U20969 ( .B1(n26058), .B2(matrix_mul_2D_3__5__7_), .C1(n25366), 
        .C2(matrix_mul_2D_3__7__7_), .A(n4847), .ZN(n4846) );
  OAI22_X1 U20970 ( .A1(n2299), .A2(n22734), .B1(n2314), .B2(n22739), .ZN(
        n4847) );
  AOI221_X1 U20971 ( .B1(n26072), .B2(matrix_mul_2D_3__5__8_), .C1(n23967), 
        .C2(matrix_mul_2D_3__7__8_), .A(n4843), .ZN(n4842) );
  OAI22_X1 U20972 ( .A1(n2298), .A2(n22735), .B1(n2313), .B2(n22740), .ZN(
        n4843) );
  AOI221_X1 U20973 ( .B1(n21465), .B2(matrix_mul_2D_3__5__9_), .C1(n23975), 
        .C2(matrix_mul_2D_3__7__9_), .A(n48390), .ZN(n48380) );
  OAI22_X1 U20974 ( .A1(n2297), .A2(n19290), .B1(n2312), .B2(n26668), .ZN(
        n48390) );
  AOI221_X1 U20975 ( .B1(n26763), .B2(matrix_mul_2D_3__5__10_), .C1(n25239), 
        .C2(matrix_mul_2D_3__7__10_), .A(n48350), .ZN(n48340) );
  OAI22_X1 U20976 ( .A1(n2296), .A2(n24088), .B1(n2311), .B2(n26668), .ZN(
        n48350) );
  AOI221_X1 U20977 ( .B1(n18496), .B2(matrix_mul_2D_3__5__11_), .C1(n26624), 
        .C2(matrix_mul_2D_3__7__11_), .A(n48310), .ZN(n48300) );
  OAI22_X1 U20978 ( .A1(n2295), .A2(n24991), .B1(n2310), .B2(n24994), .ZN(
        n48310) );
  AOI221_X1 U20979 ( .B1(n26001), .B2(matrix_mul_2D_3__5__12_), .C1(n25025), 
        .C2(matrix_mul_2D_3__7__12_), .A(n48270), .ZN(n48260) );
  OAI22_X1 U20980 ( .A1(n2294), .A2(n24090), .B1(n2309), .B2(n24094), .ZN(
        n48270) );
  AOI221_X1 U20981 ( .B1(n19248), .B2(matrix_mul_2D_3__5__13_), .C1(n17103), 
        .C2(matrix_mul_2D_3__7__13_), .A(n48230), .ZN(n48220) );
  OAI22_X1 U20982 ( .A1(n2293), .A2(n20789), .B1(n2308), .B2(n20791), .ZN(
        n48230) );
  AOI221_X1 U20983 ( .B1(n26078), .B2(matrix_mul_2D_3__5__14_), .C1(n19064), 
        .C2(matrix_mul_2D_3__7__14_), .A(n4817), .ZN(n4816) );
  OAI22_X1 U20984 ( .A1(n2292), .A2(n24091), .B1(n2307), .B2(n24095), .ZN(
        n4817) );
  NAND2_X1 U20985 ( .A1(n5105), .A2(n5106), .ZN(mul_outcome[167]) );
  AOI221_X1 U20986 ( .B1(n24310), .B2(n17283), .C1(n24939), .C2(n17271), .A(
        n27727), .ZN(n5105) );
  AOI221_X1 U20987 ( .B1(n19238), .B2(n17355), .C1(n260801), .C2(n17343), .A(
        n27768), .ZN(n5106) );
  INV_X1 U20988 ( .A(n5109), .ZN(n27727) );
  NAND2_X1 U20989 ( .A1(n5118), .A2(n5119), .ZN(mul_outcome[164]) );
  AOI221_X1 U20990 ( .B1(n22427), .B2(n17289), .C1(n24941), .C2(n17277), .A(
        n277301), .ZN(n5118) );
  AOI221_X1 U20991 ( .B1(n21381), .B2(n17361), .C1(n26056), .C2(n17349), .A(
        n27771), .ZN(n5119) );
  INV_X1 U20992 ( .A(n5121), .ZN(n277301) );
  AOI221_X1 U20993 ( .B1(n25656), .B2(matrix_mul_2D_7__0__0_), .C1(n21490), 
        .C2(matrix_mul_2D_7__1__0_), .A(n5199), .ZN(n5198) );
  OAI22_X1 U20994 ( .A1(n28160), .A2(n24661), .B1(n2801), .B2(n25345), .ZN(
        n5199) );
  AOI221_X1 U20995 ( .B1(n256501), .B2(matrix_mul_2D_7__0__1_), .C1(n21463), 
        .C2(matrix_mul_2D_7__1__1_), .A(n5195), .ZN(n5194) );
  OAI22_X1 U20996 ( .A1(n28150), .A2(n26516), .B1(n2800), .B2(n20748), .ZN(
        n5195) );
  AOI221_X1 U20997 ( .B1(n25652), .B2(matrix_mul_2D_7__0__2_), .C1(n260001), 
        .C2(matrix_mul_2D_7__1__2_), .A(n5191), .ZN(n5190) );
  OAI22_X1 U20998 ( .A1(n2814), .A2(n22451), .B1(n2799), .B2(n20742), .ZN(
        n5191) );
  AOI221_X1 U20999 ( .B1(n25656), .B2(matrix_mul_2D_7__0__3_), .C1(n21834), 
        .C2(matrix_mul_2D_7__1__3_), .A(n51830), .ZN(n51820) );
  OAI22_X1 U21000 ( .A1(n2813), .A2(n24654), .B1(n2798), .B2(n20740), .ZN(
        n51830) );
  AOI221_X1 U21001 ( .B1(n256501), .B2(matrix_mul_2D_7__0__4_), .C1(n21505), 
        .C2(matrix_mul_2D_7__1__4_), .A(n51790), .ZN(n51780) );
  OAI22_X1 U21002 ( .A1(n2812), .A2(n26518), .B1(n2797), .B2(n19091), .ZN(
        n51790) );
  AOI221_X1 U21003 ( .B1(n25652), .B2(matrix_mul_2D_7__0__5_), .C1(n21505), 
        .C2(matrix_mul_2D_7__1__5_), .A(n51750), .ZN(n51740) );
  OAI22_X1 U21004 ( .A1(n28110), .A2(n22949), .B1(n2796), .B2(n25346), .ZN(
        n51750) );
  AOI221_X1 U21005 ( .B1(n21390), .B2(matrix_mul_2D_7__0__6_), .C1(n17119), 
        .C2(matrix_mul_2D_7__1__6_), .A(n51710), .ZN(n51700) );
  OAI22_X1 U21006 ( .A1(n2810), .A2(n22466), .B1(n2795), .B2(n19021), .ZN(
        n51710) );
  AOI221_X1 U21007 ( .B1(n21377), .B2(matrix_mul_2D_7__0__7_), .C1(n21492), 
        .C2(matrix_mul_2D_7__1__7_), .A(n5167), .ZN(n5166) );
  OAI22_X1 U21008 ( .A1(n2809), .A2(n22463), .B1(n2794), .B2(n21150), .ZN(
        n5167) );
  AOI221_X1 U21009 ( .B1(n21382), .B2(matrix_mul_2D_7__0__8_), .C1(n26779), 
        .C2(matrix_mul_2D_7__1__8_), .A(n5163), .ZN(n5162) );
  OAI22_X1 U21010 ( .A1(n2808), .A2(n22463), .B1(n2793), .B2(n26678), .ZN(
        n5163) );
  AOI221_X1 U21011 ( .B1(n25655), .B2(matrix_mul_2D_7__0__9_), .C1(n21434), 
        .C2(matrix_mul_2D_7__1__9_), .A(n5159), .ZN(n5158) );
  OAI22_X1 U21012 ( .A1(n2807), .A2(n24667), .B1(n2792), .B2(n20744), .ZN(
        n5159) );
  AOI221_X1 U21013 ( .B1(n21378), .B2(matrix_mul_2D_7__0__10_), .C1(n25907), 
        .C2(matrix_mul_2D_7__1__10_), .A(n5155), .ZN(n5154) );
  OAI22_X1 U21014 ( .A1(n2806), .A2(n23451), .B1(n2791), .B2(n26682), .ZN(
        n5155) );
  AOI221_X1 U21015 ( .B1(n19238), .B2(matrix_mul_2D_7__0__11_), .C1(n25907), 
        .C2(matrix_mul_2D_7__1__11_), .A(n5151), .ZN(n51500) );
  OAI22_X1 U21016 ( .A1(n2805), .A2(n24665), .B1(n2790), .B2(n25521), .ZN(
        n5151) );
  AOI221_X1 U21017 ( .B1(n21389), .B2(matrix_mul_2D_7__0__12_), .C1(n21500), 
        .C2(matrix_mul_2D_7__1__12_), .A(n51470), .ZN(n51460) );
  OAI22_X1 U21018 ( .A1(n2804), .A2(n22454), .B1(n2789), .B2(n22762), .ZN(
        n51470) );
  AOI221_X1 U21019 ( .B1(n21378), .B2(matrix_mul_2D_7__0__13_), .C1(n17119), 
        .C2(matrix_mul_2D_7__1__13_), .A(n51390), .ZN(n51380) );
  OAI22_X1 U21020 ( .A1(n2803), .A2(n24662), .B1(n2788), .B2(n25094), .ZN(
        n51390) );
  AOI221_X1 U21021 ( .B1(n21381), .B2(matrix_mul_2D_7__0__14_), .C1(n26754), 
        .C2(matrix_mul_2D_7__1__14_), .A(n5132), .ZN(n5131) );
  OAI22_X1 U21022 ( .A1(n2802), .A2(n24668), .B1(n2787), .B2(n19179), .ZN(
        n5132) );
  NAND3_X1 U21023 ( .A1(n50890), .A2(n50900), .A3(n50910), .ZN(mul_outcome[19]) );
  AOI22_X1 U21024 ( .A1(n26982), .A2(n17909), .B1(n26704), .B2(n17969), .ZN(
        n50890) );
  AOI22_X1 U21025 ( .A1(n265101), .A2(n17981), .B1(n26711), .B2(n17957), .ZN(
        n50900) );
  AOI221_X1 U21026 ( .B1(n25938), .B2(n17933), .C1(n17945), .C2(n19078), .A(
        n27784), .ZN(n50910) );
  NAND3_X1 U21027 ( .A1(n50810), .A2(n50820), .A3(n50830), .ZN(mul_outcome[20]) );
  AOI22_X1 U21028 ( .A1(n26984), .A2(n17907), .B1(n24945), .B2(n17967), .ZN(
        n50810) );
  AOI22_X1 U21029 ( .A1(n26512), .A2(n17979), .B1(n22787), .B2(n17955), .ZN(
        n50820) );
  AOI221_X1 U21030 ( .B1(n25944), .B2(n17931), .C1(n17943), .C2(n25313), .A(
        n27783), .ZN(n50830) );
  NAND3_X1 U21031 ( .A1(n5097), .A2(n5098), .A3(n5099), .ZN(mul_outcome[17])
         );
  AOI22_X1 U21032 ( .A1(n26980), .A2(n17913), .B1(n24152), .B2(n17973), .ZN(
        n5097) );
  AOI22_X1 U21033 ( .A1(n22441), .A2(n17985), .B1(n24931), .B2(n17961), .ZN(
        n5098) );
  AOI221_X1 U21034 ( .B1(n259501), .B2(n17937), .C1(n17949), .C2(n26716), .A(
        n27786), .ZN(n5099) );
  NAND3_X1 U21035 ( .A1(n51410), .A2(n51420), .A3(n51430), .ZN(mul_outcome[15]) );
  AOI22_X1 U21036 ( .A1(n26978), .A2(n17917), .B1(n19085), .B2(n17977), .ZN(
        n51410) );
  AOI22_X1 U21037 ( .A1(n22444), .A2(n17989), .B1(n19081), .B2(n17965), .ZN(
        n51420) );
  AOI221_X1 U21038 ( .B1(n25943), .B2(n17941), .C1(n17953), .C2(n26716), .A(
        n27788), .ZN(n51430) );
  NAND3_X1 U21039 ( .A1(n48810), .A2(n48820), .A3(n48830), .ZN(mul_outcome[62]) );
  AOI22_X1 U21040 ( .A1(n27054), .A2(n17811), .B1(n19228), .B2(n17799), .ZN(
        n48810) );
  AOI22_X1 U21041 ( .A1(n27068), .A2(n17835), .B1(n27080), .B2(n17823), .ZN(
        n48820) );
  AOI221_X1 U21042 ( .B1(n27092), .B2(n17787), .C1(n19232), .C2(n17775), .A(
        n27743), .ZN(n48830) );
  AOI221_X1 U21043 ( .B1(n27087), .B2(matrix_mul_2D_2__4__0_), .C1(n21359), 
        .C2(matrix_mul_2D_2__5__0_), .A(n4978), .ZN(n4977) );
  OAI22_X1 U21044 ( .A1(n2240), .A2(n21140), .B1(n2225), .B2(n26551), .ZN(
        n4978) );
  AOI221_X1 U21045 ( .B1(n27088), .B2(matrix_mul_2D_2__4__1_), .C1(n21348), 
        .C2(matrix_mul_2D_2__5__1_), .A(n49740), .ZN(n49730) );
  OAI22_X1 U21046 ( .A1(n2239), .A2(n21150), .B1(n2224), .B2(n22510), .ZN(
        n49740) );
  AOI221_X1 U21047 ( .B1(n27089), .B2(matrix_mul_2D_2__4__2_), .C1(n25638), 
        .C2(matrix_mul_2D_2__5__2_), .A(n49700), .ZN(n49690) );
  OAI22_X1 U21048 ( .A1(n2238), .A2(n22759), .B1(n2223), .B2(n26532), .ZN(
        n49700) );
  AOI221_X1 U21049 ( .B1(n27090), .B2(matrix_mul_2D_2__4__3_), .C1(n25641), 
        .C2(matrix_mul_2D_2__5__3_), .A(n49660), .ZN(n49650) );
  OAI22_X1 U21050 ( .A1(n2237), .A2(n25516), .B1(n2222), .B2(n26521), .ZN(
        n49660) );
  AOI221_X1 U21051 ( .B1(n27091), .B2(matrix_mul_2D_2__4__4_), .C1(n25637), 
        .C2(matrix_mul_2D_2__5__4_), .A(n49620), .ZN(n49610) );
  OAI22_X1 U21052 ( .A1(n2236), .A2(n24970), .B1(n2221), .B2(n26553), .ZN(
        n49620) );
  AOI221_X1 U21053 ( .B1(n27092), .B2(matrix_mul_2D_2__4__5_), .C1(n19232), 
        .C2(matrix_mul_2D_2__5__5_), .A(n4958), .ZN(n4957) );
  OAI22_X1 U21054 ( .A1(n2235), .A2(n24965), .B1(n2220), .B2(n22475), .ZN(
        n4958) );
  AOI221_X1 U21055 ( .B1(n27097), .B2(matrix_mul_2D_2__4__6_), .C1(n21358), 
        .C2(matrix_mul_2D_2__5__6_), .A(n4954), .ZN(n4953) );
  OAI22_X1 U21056 ( .A1(n2234), .A2(n24961), .B1(n2219), .B2(n22507), .ZN(
        n4954) );
  AOI221_X1 U21057 ( .B1(n27093), .B2(matrix_mul_2D_2__4__7_), .C1(n21347), 
        .C2(matrix_mul_2D_2__5__7_), .A(n4950), .ZN(n4949) );
  OAI22_X1 U21058 ( .A1(n2233), .A2(n24963), .B1(n2218), .B2(n23685), .ZN(
        n4950) );
  AOI221_X1 U21059 ( .B1(n27094), .B2(matrix_mul_2D_2__4__8_), .C1(n25638), 
        .C2(matrix_mul_2D_2__5__8_), .A(n4942), .ZN(n4941) );
  OAI22_X1 U21060 ( .A1(n2232), .A2(n21148), .B1(n2217), .B2(n26534), .ZN(
        n4942) );
  AOI221_X1 U21061 ( .B1(n27096), .B2(matrix_mul_2D_2__4__9_), .C1(n25641), 
        .C2(matrix_mul_2D_2__5__9_), .A(n4938), .ZN(n4937) );
  OAI22_X1 U21062 ( .A1(n2231), .A2(n24959), .B1(n2216), .B2(n26523), .ZN(
        n4938) );
  AOI221_X1 U21063 ( .B1(n27093), .B2(matrix_mul_2D_2__4__10_), .C1(n25637), 
        .C2(matrix_mul_2D_2__5__10_), .A(n4934), .ZN(n4933) );
  OAI22_X1 U21064 ( .A1(n2230), .A2(n25522), .B1(n2215), .B2(n22478), .ZN(
        n4934) );
  AOI221_X1 U21065 ( .B1(n27094), .B2(matrix_mul_2D_2__4__11_), .C1(n21350), 
        .C2(matrix_mul_2D_2__5__11_), .A(n4930), .ZN(n4929) );
  OAI22_X1 U21066 ( .A1(n2229), .A2(n25521), .B1(n2214), .B2(n22460), .ZN(
        n4930) );
  AOI221_X1 U21067 ( .B1(n25642), .B2(matrix_mul_2D_6__0__0_), .C1(n27032), 
        .C2(matrix_mul_2D_6__1__0_), .A(n5295), .ZN(n5294) );
  OAI22_X1 U21068 ( .A1(n268400), .A2(n25346), .B1(n2669), .B2(n22506), .ZN(
        n5295) );
  AOI221_X1 U21069 ( .B1(n25643), .B2(matrix_mul_2D_6__0__1_), .C1(n27033), 
        .C2(matrix_mul_2D_6__1__1_), .A(n5291), .ZN(n5290) );
  OAI22_X1 U21070 ( .A1(n268300), .A2(n20745), .B1(n2668), .B2(n26535), .ZN(
        n5291) );
  AOI221_X1 U21071 ( .B1(n19233), .B2(matrix_mul_2D_6__0__2_), .C1(n27034), 
        .C2(matrix_mul_2D_6__1__2_), .A(n5287), .ZN(n5286) );
  OAI22_X1 U21072 ( .A1(n268200), .A2(n25344), .B1(n2667), .B2(n22456), .ZN(
        n5287) );
  AOI221_X1 U21073 ( .B1(n25642), .B2(matrix_mul_2D_6__0__3_), .C1(n27035), 
        .C2(matrix_mul_2D_6__1__3_), .A(n5283), .ZN(n5282) );
  OAI22_X1 U21074 ( .A1(n268100), .A2(n26679), .B1(n2666), .B2(n22507), .ZN(
        n5283) );
  AOI221_X1 U21075 ( .B1(n25643), .B2(matrix_mul_2D_6__0__4_), .C1(n27036), 
        .C2(matrix_mul_2D_6__1__4_), .A(n5275), .ZN(n5274) );
  OAI22_X1 U21076 ( .A1(n268000), .A2(n20749), .B1(n2665), .B2(n26533), .ZN(
        n5275) );
  AOI221_X1 U21077 ( .B1(n256401), .B2(matrix_mul_2D_6__0__5_), .C1(n27037), 
        .C2(matrix_mul_2D_6__1__5_), .A(n5271), .ZN(n52700) );
  OAI22_X1 U21078 ( .A1(n267900), .A2(n22763), .B1(n2664), .B2(n22503), .ZN(
        n5271) );
  AOI221_X1 U21079 ( .B1(n21361), .B2(matrix_mul_2D_6__0__6_), .C1(n27042), 
        .C2(matrix_mul_2D_6__1__6_), .A(n52670), .ZN(n52660) );
  OAI22_X1 U21080 ( .A1(n267800), .A2(n20741), .B1(n2663), .B2(n23686), .ZN(
        n52670) );
  AOI221_X1 U21081 ( .B1(n21365), .B2(matrix_mul_2D_6__0__7_), .C1(n27038), 
        .C2(matrix_mul_2D_6__1__7_), .A(n52630), .ZN(n52620) );
  OAI22_X1 U21082 ( .A1(n267700), .A2(n19177), .B1(n2662), .B2(n22474), .ZN(
        n52630) );
  AOI221_X1 U21083 ( .B1(n256401), .B2(matrix_mul_2D_6__0__8_), .C1(n27039), 
        .C2(matrix_mul_2D_6__1__8_), .A(n52590), .ZN(n52580) );
  OAI22_X1 U21084 ( .A1(n267600), .A2(n20743), .B1(n2661), .B2(n26524), .ZN(
        n52590) );
  AOI221_X1 U21085 ( .B1(n21362), .B2(matrix_mul_2D_6__0__9_), .C1(n27041), 
        .C2(matrix_mul_2D_6__1__9_), .A(n52550), .ZN(n52540) );
  OAI22_X1 U21086 ( .A1(n267500), .A2(n19092), .B1(n2660), .B2(n22477), .ZN(
        n52550) );
  AOI221_X1 U21087 ( .B1(n21366), .B2(matrix_mul_2D_6__0__10_), .C1(n27038), 
        .C2(matrix_mul_2D_6__1__10_), .A(n52510), .ZN(n52500) );
  OAI22_X1 U21088 ( .A1(n267400), .A2(n19021), .B1(n2659), .B2(n22459), .ZN(
        n52510) );
  AOI221_X1 U21089 ( .B1(n21354), .B2(matrix_mul_2D_6__0__11_), .C1(n27039), 
        .C2(matrix_mul_2D_6__1__11_), .A(n5247), .ZN(n5246) );
  OAI22_X1 U21090 ( .A1(n2673), .A2(n26681), .B1(n2658), .B2(n26522), .ZN(
        n5247) );
  NAND3_X1 U21091 ( .A1(n5323), .A2(n5324), .A3(n5325), .ZN(mul_outcome[120])
         );
  AOI221_X1 U21092 ( .B1(n24398), .B2(n17485), .C1(n21496), .C2(n17473), .A(
        n27779), .ZN(n5325) );
  AOI22_X1 U21093 ( .A1(n27016), .A2(n17557), .B1(n22896), .B2(n17545), .ZN(
        n5324) );
  AOI22_X1 U21094 ( .A1(n27013), .A2(n17533), .B1(n25904), .B2(n17521), .ZN(
        n5323) );
  AOI22_X1 U21095 ( .A1(n27012), .A2(matrix_mul_2D_5__2__0_), .B1(n26002), 
        .B2(matrix_mul_2D_5__3__0_), .ZN(n53910) );
  AOI22_X1 U21096 ( .A1(n27003), .A2(matrix_mul_2D_5__2__1_), .B1(n21433), 
        .B2(matrix_mul_2D_5__3__1_), .ZN(n53870) );
  AOI22_X1 U21097 ( .A1(n27004), .A2(matrix_mul_2D_5__2__2_), .B1(n22826), 
        .B2(matrix_mul_2D_5__3__2_), .ZN(n5383) );
  AOI22_X1 U21098 ( .A1(n27005), .A2(matrix_mul_2D_5__2__3_), .B1(n26079), 
        .B2(matrix_mul_2D_5__3__3_), .ZN(n5379) );
  AOI22_X1 U21099 ( .A1(n27006), .A2(matrix_mul_2D_5__2__4_), .B1(n26073), 
        .B2(matrix_mul_2D_5__3__4_), .ZN(n5375) );
  AOI22_X1 U21100 ( .A1(n27007), .A2(matrix_mul_2D_5__2__5_), .B1(n26306), 
        .B2(matrix_mul_2D_5__3__5_), .ZN(n5367) );
  AOI22_X1 U21101 ( .A1(n27008), .A2(matrix_mul_2D_5__2__6_), .B1(n22871), 
        .B2(matrix_mul_2D_5__3__6_), .ZN(n5363) );
  AOI22_X1 U21102 ( .A1(n27009), .A2(matrix_mul_2D_5__2__7_), .B1(n26056), 
        .B2(matrix_mul_2D_5__3__7_), .ZN(n53590) );
  AOI22_X1 U21103 ( .A1(n27010), .A2(matrix_mul_2D_5__2__8_), .B1(n26059), 
        .B2(matrix_mul_2D_5__3__8_), .ZN(n53550) );
  AOI22_X1 U21104 ( .A1(n27008), .A2(matrix_mul_2D_5__2__9_), .B1(n260801), 
        .B2(matrix_mul_2D_5__3__9_), .ZN(n53510) );
  AOI22_X1 U21105 ( .A1(n27009), .A2(matrix_mul_2D_5__2__10_), .B1(n25918), 
        .B2(matrix_mul_2D_5__3__10_), .ZN(n53470) );
  AOI22_X1 U21106 ( .A1(n27010), .A2(matrix_mul_2D_5__2__11_), .B1(n17078), 
        .B2(matrix_mul_2D_5__3__11_), .ZN(n53430) );
  OAI22_X1 U21107 ( .A1(n23934), .A2(n11862), .B1(n22004), .B2(n1779), .ZN(
        n6896) );
  OAI22_X1 U21108 ( .A1(n23886), .A2(n11876), .B1(n22040), .B2(n1777), .ZN(
        n68940) );
  OAI22_X1 U21109 ( .A1(n25230), .A2(n11890), .B1(n22076), .B2(n1775), .ZN(
        n68920) );
  OAI22_X1 U21110 ( .A1(n22607), .A2(n11904), .B1(n22112), .B2(n1773), .ZN(
        n68900) );
  OAI22_X1 U21111 ( .A1(n22582), .A2(n11918), .B1(n22344), .B2(n1771), .ZN(
        n68880) );
  OAI22_X1 U21112 ( .A1(n23926), .A2(n11932), .B1(n22368), .B2(n1769), .ZN(
        n68860) );
  OAI22_X1 U21113 ( .A1(n23878), .A2(n11946), .B1(n22392), .B2(n1767), .ZN(
        n68840) );
  OAI22_X1 U21114 ( .A1(n24974), .A2(n11960), .B1(n22416), .B2(n1765), .ZN(
        n68820) );
  OAI22_X1 U21115 ( .A1(n23922), .A2(n11974), .B1(n22152), .B2(n1763), .ZN(
        n68800) );
  OAI22_X1 U21116 ( .A1(n23874), .A2(n11988), .B1(n22197), .B2(n1761), .ZN(
        n68780) );
  OAI22_X1 U21117 ( .A1(n24978), .A2(n12002), .B1(n22243), .B2(n1759), .ZN(
        n68760) );
  OAI22_X1 U21118 ( .A1(n22580), .A2(n12016), .B1(n22278), .B2(n1757), .ZN(
        n68740) );
  OAI22_X1 U21119 ( .A1(n23909), .A2(n12030), .B1(n22158), .B2(n1755), .ZN(
        n6872) );
  OAI22_X1 U21120 ( .A1(n23861), .A2(n12044), .B1(n22204), .B2(n1753), .ZN(
        n6870) );
  OAI22_X1 U21121 ( .A1(n24971), .A2(n12058), .B1(n22236), .B2(n1751), .ZN(
        n6868) );
  OAI22_X1 U21122 ( .A1(n22564), .A2(n12072), .B1(n22268), .B2(n1749), .ZN(
        n6866) );
  OAI22_X1 U21123 ( .A1(n23897), .A2(n12086), .B1(n22008), .B2(n1747), .ZN(
        n6864) );
  OAI22_X1 U21124 ( .A1(n23849), .A2(n12100), .B1(n22044), .B2(n1745), .ZN(
        n6862) );
  OAI22_X1 U21125 ( .A1(n20770), .A2(n12114), .B1(n22080), .B2(n1743), .ZN(
        n6860) );
  OAI22_X1 U21126 ( .A1(n22551), .A2(n12128), .B1(n22116), .B2(n1741), .ZN(
        n6858) );
  OAI22_X1 U21127 ( .A1(n23927), .A2(n12142), .B1(n21990), .B2(n1739), .ZN(
        n68560) );
  OAI22_X1 U21128 ( .A1(n23879), .A2(n12156), .B1(n22026), .B2(n1737), .ZN(
        n68540) );
  OAI22_X1 U21129 ( .A1(n24976), .A2(n12170), .B1(n22062), .B2(n1735), .ZN(
        n68520) );
  OAI22_X1 U21130 ( .A1(n22602), .A2(n12184), .B1(n22098), .B2(n1733), .ZN(
        n68500) );
  OAI22_X1 U21131 ( .A1(n22566), .A2(n12198), .B1(n22338), .B2(n1731), .ZN(
        n68480) );
  OAI22_X1 U21132 ( .A1(n23914), .A2(n12212), .B1(n22362), .B2(n1729), .ZN(
        n68460) );
  OAI22_X1 U21133 ( .A1(n23866), .A2(n12226), .B1(n22386), .B2(n1727), .ZN(
        n68440) );
  OAI22_X1 U21134 ( .A1(n20766), .A2(n12240), .B1(n22410), .B2(n1725), .ZN(
        n68420) );
  OAI22_X1 U21135 ( .A1(n23915), .A2(n12254), .B1(n22134), .B2(n1723), .ZN(
        n6840) );
  OAI22_X1 U21136 ( .A1(n23867), .A2(n12268), .B1(n22179), .B2(n1721), .ZN(
        n6838) );
  OAI22_X1 U21137 ( .A1(n25349), .A2(n12282), .B1(n22229), .B2(n1719), .ZN(
        n6836) );
  OAI22_X1 U21138 ( .A1(n22590), .A2(n12296), .B1(n22265), .B2(n1717), .ZN(
        n6834) );
  OAI22_X1 U21139 ( .A1(n22546), .A2(n1779), .B1(n21720), .B2(n1715), .ZN(
        n6832) );
  OAI22_X1 U21140 ( .A1(n23902), .A2(n1777), .B1(n21736), .B2(n1713), .ZN(
        n6830) );
  OAI22_X1 U21141 ( .A1(n23854), .A2(n1775), .B1(n21752), .B2(n1711), .ZN(
        n6828) );
  OAI22_X1 U21142 ( .A1(n23964), .A2(n1773), .B1(n21768), .B2(n1709), .ZN(
        n6826) );
  OAI22_X1 U21143 ( .A1(n23904), .A2(n1771), .B1(n21659), .B2(n1707), .ZN(
        n6824) );
  OAI22_X1 U21144 ( .A1(n23856), .A2(n1769), .B1(n21667), .B2(n1705), .ZN(
        n6822) );
  OAI22_X1 U21145 ( .A1(n25361), .A2(n1767), .B1(n21675), .B2(n1703), .ZN(
        n6820) );
  OAI22_X1 U21146 ( .A1(n22574), .A2(n1765), .B1(n21683), .B2(n1701), .ZN(
        n6818) );
  OAI22_X1 U21147 ( .A1(n22594), .A2(n1763), .B1(n21724), .B2(n1699), .ZN(
        n6816) );
  OAI22_X1 U21148 ( .A1(n23890), .A2(n1761), .B1(n21740), .B2(n1697), .ZN(
        n6814) );
  OAI22_X1 U21149 ( .A1(n23842), .A2(n1759), .B1(n21756), .B2(n1695), .ZN(
        n6812) );
  OAI22_X1 U21150 ( .A1(n19098), .A2(n1757), .B1(n21772), .B2(n1693), .ZN(
        n6810) );
  OAI22_X1 U21151 ( .A1(n23891), .A2(n1755), .B1(n21691), .B2(n1691), .ZN(
        n6808) );
  OAI22_X1 U21152 ( .A1(n23843), .A2(n1753), .B1(n21699), .B2(n1689), .ZN(
        n6806) );
  OAI22_X1 U21153 ( .A1(n19097), .A2(n1751), .B1(n21707), .B2(n1687), .ZN(
        n6804) );
  OAI22_X1 U21154 ( .A1(n22546), .A2(n1749), .B1(n23583), .B2(n1685), .ZN(
        n68020) );
  OAI22_X1 U21155 ( .A1(n20686), .A2(n1747), .B1(n22149), .B2(n1683), .ZN(
        n68000) );
  OAI22_X1 U21156 ( .A1(n20654), .A2(n1745), .B1(n22194), .B2(n1681), .ZN(
        n67980) );
  OAI22_X1 U21157 ( .A1(n19063), .A2(n1743), .B1(n22241), .B2(n1679), .ZN(
        n67960) );
  OAI22_X1 U21158 ( .A1(n22599), .A2(n1741), .B1(n22275), .B2(n1677), .ZN(
        n67940) );
  OAI22_X1 U21159 ( .A1(n24849), .A2(n1739), .B1(n22001), .B2(n1675), .ZN(
        n67920) );
  OAI22_X1 U21160 ( .A1(n24833), .A2(n1737), .B1(n22037), .B2(n1673), .ZN(
        n67900) );
  OAI22_X1 U21161 ( .A1(n25364), .A2(n1735), .B1(n22073), .B2(n1671), .ZN(
        n67880) );
  OAI22_X1 U21162 ( .A1(n22586), .A2(n1733), .B1(n22109), .B2(n1669), .ZN(
        n67860) );
  OAI22_X1 U21163 ( .A1(n24844), .A2(n1731), .B1(n264101), .B2(n1667), .ZN(
        n67840) );
  OAI22_X1 U21164 ( .A1(n24827), .A2(n1729), .B1(n26416), .B2(n1665), .ZN(
        n67820) );
  OAI22_X1 U21165 ( .A1(n24120), .A2(n1727), .B1(n26422), .B2(n1663), .ZN(
        n6780) );
  OAI22_X1 U21166 ( .A1(n22571), .A2(n1725), .B1(n26428), .B2(n1661), .ZN(
        n6778) );
  OAI22_X1 U21167 ( .A1(n22578), .A2(n1723), .B1(n22341), .B2(n1659), .ZN(
        n6776) );
  OAI22_X1 U21168 ( .A1(n20679), .A2(n1721), .B1(n22365), .B2(n1657), .ZN(
        n6774) );
  OAI22_X1 U21169 ( .A1(n20647), .A2(n1719), .B1(n22389), .B2(n1655), .ZN(
        n6772) );
  OAI22_X1 U21170 ( .A1(n24132), .A2(n1717), .B1(n22413), .B2(n1653), .ZN(
        n6770) );
  OAI22_X1 U21171 ( .A1(n25044), .A2(n1715), .B1(n26436), .B2(n1651), .ZN(
        n6768) );
  OAI22_X1 U21172 ( .A1(n25061), .A2(n1713), .B1(n26445), .B2(n1649), .ZN(
        n6766) );
  OAI22_X1 U21173 ( .A1(n24138), .A2(n1711), .B1(n264501), .B2(n1647), .ZN(
        n67640) );
  OAI22_X1 U21174 ( .A1(n22559), .A2(n1709), .B1(n68), .B2(n1645), .ZN(n67620)
         );
  OAI22_X1 U21175 ( .A1(n22562), .A2(n1707), .B1(n22335), .B2(n1643), .ZN(
        n67600) );
  OAI22_X1 U21176 ( .A1(n20822), .A2(n1705), .B1(n22359), .B2(n1641), .ZN(
        n67580) );
  OAI22_X1 U21177 ( .A1(n20846), .A2(n1703), .B1(n22383), .B2(n1639), .ZN(
        n67560) );
  OAI22_X1 U21178 ( .A1(n24107), .A2(n1701), .B1(n22407), .B2(n1637), .ZN(
        n67540) );
  OAI22_X1 U21179 ( .A1(n24855), .A2(n1699), .B1(n26407), .B2(n1635), .ZN(
        n67520) );
  OAI22_X1 U21180 ( .A1(n24839), .A2(n1697), .B1(n26413), .B2(n1633), .ZN(
        n67500) );
  OAI22_X1 U21181 ( .A1(n24114), .A2(n1695), .B1(n26419), .B2(n1631), .ZN(
        n6748) );
  OAI22_X1 U21182 ( .A1(n22595), .A2(n1693), .B1(n26425), .B2(n1629), .ZN(
        n6746) );
  OAI22_X1 U21183 ( .A1(n22558), .A2(n1691), .B1(n26213), .B2(n1627), .ZN(
        n6744) );
  OAI22_X1 U21184 ( .A1(n20830), .A2(n1689), .B1(n26221), .B2(n1625), .ZN(
        n6742) );
  OAI22_X1 U21185 ( .A1(n20854), .A2(n1687), .B1(n26229), .B2(n1623), .ZN(
        n6740) );
  OAI22_X1 U21186 ( .A1(n24126), .A2(n1685), .B1(n26237), .B2(n1621), .ZN(
        n6738) );
  OAI22_X1 U21187 ( .A1(n20677), .A2(n1683), .B1(n26431), .B2(n1619), .ZN(
        n6736) );
  OAI22_X1 U21188 ( .A1(n20645), .A2(n1681), .B1(n26441), .B2(n1617), .ZN(
        n6734) );
  OAI22_X1 U21189 ( .A1(n19095), .A2(n1679), .B1(n26449), .B2(n1615), .ZN(
        n6732) );
  OAI22_X1 U21190 ( .A1(n22583), .A2(n1677), .B1(n24362), .B2(n1613), .ZN(
        n6730) );
  OAI22_X1 U21191 ( .A1(n24847), .A2(n1675), .B1(n26183), .B2(n1611), .ZN(
        n6728) );
  OAI22_X1 U21192 ( .A1(n24830), .A2(n1673), .B1(n26187), .B2(n1609), .ZN(
        n6726) );
  OAI22_X1 U21193 ( .A1(n25350), .A2(n1671), .B1(n26191), .B2(n1607), .ZN(
        n6724) );
  OAI22_X1 U21194 ( .A1(n22567), .A2(n1669), .B1(n24368), .B2(n1605), .ZN(
        n6722) );
  OAI22_X1 U21195 ( .A1(n24843), .A2(n1667), .B1(n26167), .B2(n1603), .ZN(
        n67200) );
  OAI22_X1 U21196 ( .A1(n24826), .A2(n1665), .B1(n26171), .B2(n1601), .ZN(
        n67180) );
  OAI22_X1 U21197 ( .A1(n19100), .A2(n1663), .B1(n26175), .B2(n1599), .ZN(
        n67160) );
  OAI22_X1 U21198 ( .A1(n23760), .A2(n1661), .B1(n26179), .B2(n1597), .ZN(
        n67140) );
  OAI22_X1 U21199 ( .A1(n23932), .A2(n1659), .B1(n26409), .B2(n1595), .ZN(
        n67120) );
  OAI22_X1 U21200 ( .A1(n23884), .A2(n1657), .B1(n26415), .B2(n1593), .ZN(
        n67100) );
  OAI22_X1 U21201 ( .A1(n25357), .A2(n1655), .B1(n26421), .B2(n1591), .ZN(
        n67080) );
  OAI22_X1 U21202 ( .A1(n23838), .A2(n1653), .B1(n26427), .B2(n1589), .ZN(
        n67060) );
  OAI22_X1 U21203 ( .A1(n23837), .A2(n1651), .B1(n26215), .B2(n1587), .ZN(
        n67040) );
  OAI22_X1 U21204 ( .A1(n20661), .A2(n1649), .B1(n26223), .B2(n1585), .ZN(
        n67020) );
  OAI22_X1 U21205 ( .A1(n20628), .A2(n1647), .B1(n26231), .B2(n1583), .ZN(
        n67000) );
  OAI22_X1 U21206 ( .A1(n25241), .A2(n1645), .B1(n26239), .B2(n1581), .ZN(
        n6698) );
  OAI22_X1 U21207 ( .A1(n23920), .A2(n1643), .B1(n26435), .B2(n1579), .ZN(
        n6696) );
  OAI22_X1 U21208 ( .A1(n23872), .A2(n1641), .B1(n26867), .B2(n1577), .ZN(
        n6694) );
  OAI22_X1 U21209 ( .A1(n24134), .A2(n1639), .B1(n26451), .B2(n1575), .ZN(
        n6692) );
  OAI22_X1 U21210 ( .A1(n22578), .A2(n1637), .B1(n26455), .B2(n1573), .ZN(
        n6690) );
  OAI22_X1 U21211 ( .A1(n23813), .A2(n1635), .B1(n26483), .B2(n1571), .ZN(
        n6688) );
  OAI22_X1 U21212 ( .A1(n20813), .A2(n1633), .B1(n26487), .B2(n1569), .ZN(
        n6686) );
  OAI22_X1 U21213 ( .A1(n20837), .A2(n1631), .B1(n26491), .B2(n1567), .ZN(
        n6684) );
  OAI22_X1 U21214 ( .A1(n25360), .A2(n1629), .B1(n26495), .B2(n1565), .ZN(
        n66820) );
  OAI22_X1 U21215 ( .A1(n23908), .A2(n1627), .B1(n22012), .B2(n1563), .ZN(
        n66800) );
  OAI22_X1 U21216 ( .A1(n23860), .A2(n1625), .B1(n22048), .B2(n1561), .ZN(
        n66780) );
  OAI22_X1 U21217 ( .A1(n24110), .A2(n1623), .B1(n22084), .B2(n1559), .ZN(
        n66760) );
  OAI22_X1 U21218 ( .A1(n22562), .A2(n1621), .B1(n22120), .B2(n1557), .ZN(
        n66740) );
  OAI22_X1 U21219 ( .A1(n23789), .A2(n1619), .B1(n26482), .B2(n1555), .ZN(
        n66720) );
  OAI22_X1 U21220 ( .A1(n25038), .A2(n1617), .B1(n26486), .B2(n1553), .ZN(
        n66700) );
  OAI22_X1 U21221 ( .A1(n25054), .A2(n1615), .B1(n264901), .B2(n1551), .ZN(
        n66680) );
  OAI22_X1 U21222 ( .A1(n23961), .A2(n1613), .B1(n26494), .B2(n1549), .ZN(
        n6666) );
  OAI22_X1 U21223 ( .A1(n23896), .A2(n1611), .B1(n22163), .B2(n1547), .ZN(
        n6664) );
  OAI22_X1 U21224 ( .A1(n23848), .A2(n1609), .B1(n22210), .B2(n1545), .ZN(
        n6662) );
  OAI22_X1 U21225 ( .A1(n24122), .A2(n1607), .B1(n22240), .B2(n1543), .ZN(
        n6660) );
  OAI22_X1 U21226 ( .A1(n23754), .A2(n1605), .B1(n22274), .B2(n1541), .ZN(
        n6658) );
  OAI22_X1 U21227 ( .A1(n23926), .A2(n1603), .B1(n22140), .B2(n1539), .ZN(
        n6656) );
  OAI22_X1 U21228 ( .A1(n23878), .A2(n1601), .B1(n22186), .B2(n1537), .ZN(
        n6654) );
  OAI22_X1 U21229 ( .A1(n24140), .A2(n1599), .B1(n22234), .B2(n1535), .ZN(
        n6652) );
  OAI22_X1 U21230 ( .A1(n23832), .A2(n1597), .B1(n24366), .B2(n1533), .ZN(
        n6650) );
  OAI22_X1 U21231 ( .A1(n23914), .A2(n1595), .B1(n21994), .B2(n1531), .ZN(
        n6648) );
  OAI22_X1 U21232 ( .A1(n23866), .A2(n1593), .B1(n22030), .B2(n1529), .ZN(
        n6646) );
  OAI22_X1 U21233 ( .A1(n24116), .A2(n1591), .B1(n22066), .B2(n1527), .ZN(
        n6644) );
  OAI22_X1 U21234 ( .A1(n23814), .A2(n1589), .B1(n22102), .B2(n1525), .ZN(
        n6642) );
  OAI22_X1 U21235 ( .A1(n23902), .A2(n1587), .B1(n26166), .B2(n1523), .ZN(
        n6640) );
  OAI22_X1 U21236 ( .A1(n23854), .A2(n1585), .B1(n26170), .B2(n1521), .ZN(
        n6638) );
  OAI22_X1 U21237 ( .A1(n24127), .A2(n1583), .B1(n26174), .B2(n1519), .ZN(
        n6636) );
  OAI22_X1 U21238 ( .A1(n23790), .A2(n1581), .B1(n26178), .B2(n1517), .ZN(
        n6634) );
  OAI22_X1 U21239 ( .A1(n23759), .A2(n1579), .B1(n26212), .B2(n1515), .ZN(
        n6632) );
  OAI22_X1 U21240 ( .A1(n25040), .A2(n1577), .B1(n26220), .B2(n1513), .ZN(
        n6630) );
  OAI22_X1 U21241 ( .A1(n25056), .A2(n1575), .B1(n26228), .B2(n1511), .ZN(
        n6628) );
  OAI22_X1 U21242 ( .A1(n22675), .A2(n1573), .B1(n26236), .B2(n1509), .ZN(
        n6626) );
  OAI22_X1 U21243 ( .A1(n23890), .A2(n1571), .B1(n26182), .B2(n1507), .ZN(
        n6624) );
  OAI22_X1 U21244 ( .A1(n23842), .A2(n1569), .B1(n26186), .B2(n1505), .ZN(
        n6622) );
  OAI22_X1 U21245 ( .A1(n25236), .A2(n1567), .B1(n26190), .B2(n1503), .ZN(
        n66200) );
  OAI22_X1 U21246 ( .A1(n23748), .A2(n1565), .B1(n24363), .B2(n1501), .ZN(
        n66180) );
  OAI22_X1 U21247 ( .A1(n23831), .A2(n1563), .B1(n26214), .B2(n1499), .ZN(
        n66160) );
  OAI22_X1 U21248 ( .A1(n25046), .A2(n1561), .B1(n26222), .B2(n1497), .ZN(
        n66140) );
  OAI22_X1 U21249 ( .A1(n25063), .A2(n1559), .B1(n26230), .B2(n1495), .ZN(
        n66120) );
  OAI22_X1 U21250 ( .A1(n19061), .A2(n1557), .B1(n26238), .B2(n1493), .ZN(
        n66100) );
  OAI22_X1 U21251 ( .A1(n24853), .A2(n1555), .B1(n22006), .B2(n1491), .ZN(
        n66080) );
  OAI22_X1 U21252 ( .A1(n24837), .A2(n1553), .B1(n22042), .B2(n1489), .ZN(
        n66060) );
  OAI22_X1 U21253 ( .A1(n19056), .A2(n1551), .B1(n22078), .B2(n1487), .ZN(
        n66040) );
  OAI22_X1 U21254 ( .A1(n23826), .A2(n1549), .B1(n22114), .B2(n1485), .ZN(
        n66020) );
  OAI22_X1 U21255 ( .A1(n23807), .A2(n1547), .B1(n22346), .B2(n1483), .ZN(
        n66000) );
  OAI22_X1 U21256 ( .A1(n22672), .A2(n1545), .B1(n22370), .B2(n1481), .ZN(
        n6598) );
  OAI22_X1 U21257 ( .A1(n22640), .A2(n1543), .B1(n22394), .B2(n1479), .ZN(
        n6596) );
  OAI22_X1 U21258 ( .A1(n19062), .A2(n1541), .B1(n22418), .B2(n1477), .ZN(
        n6594) );
  OAI22_X1 U21259 ( .A1(n20671), .A2(n1539), .B1(n22156), .B2(n1475), .ZN(
        n6592) );
  OAI22_X1 U21260 ( .A1(n20638), .A2(n1537), .B1(n22201), .B2(n1473), .ZN(
        n6590) );
  OAI22_X1 U21261 ( .A1(n25359), .A2(n1535), .B1(n22246), .B2(n1471), .ZN(
        n6588) );
  OAI22_X1 U21262 ( .A1(n23808), .A2(n1533), .B1(n22282), .B2(n1469), .ZN(
        n6586) );
  OAI22_X1 U21263 ( .A1(n20824), .A2(n1531), .B1(n22161), .B2(n1467), .ZN(
        n6584) );
  OAI22_X1 U21264 ( .A1(n20848), .A2(n1529), .B1(n22207), .B2(n1465), .ZN(
        n65820) );
  OAI22_X1 U21265 ( .A1(n20760), .A2(n1527), .B1(n22237), .B2(n1463), .ZN(
        n65800) );
  OAI22_X1 U21266 ( .A1(n23784), .A2(n1525), .B1(n22270), .B2(n1461), .ZN(
        n65780) );
  OAI22_X1 U21267 ( .A1(n25049), .A2(n1523), .B1(n22010), .B2(n1459), .ZN(
        n65760) );
  OAI22_X1 U21268 ( .A1(n25066), .A2(n1521), .B1(n22046), .B2(n1457), .ZN(
        n65740) );
  OAI22_X1 U21269 ( .A1(n25229), .A2(n1519), .B1(n22082), .B2(n1455), .ZN(
        n65720) );
  OAI22_X1 U21270 ( .A1(n23766), .A2(n1517), .B1(n22118), .B2(n1453), .ZN(
        n65700) );
  OAI22_X1 U21271 ( .A1(n20682), .A2(n1515), .B1(n21992), .B2(n1451), .ZN(
        n65680) );
  OAI22_X1 U21272 ( .A1(n20650), .A2(n1513), .B1(n22028), .B2(n1449), .ZN(
        n6566) );
  OAI22_X1 U21273 ( .A1(n20768), .A2(n1511), .B1(n22064), .B2(n1447), .ZN(
        n6564) );
  OAI22_X1 U21274 ( .A1(n23820), .A2(n1509), .B1(n22100), .B2(n1445), .ZN(
        n6562) );
  OAI22_X1 U21275 ( .A1(n23783), .A2(n1507), .B1(n22340), .B2(n1443), .ZN(
        n6560) );
  OAI22_X1 U21276 ( .A1(n22664), .A2(n1505), .B1(n22364), .B2(n1441), .ZN(
        n6558) );
  OAI22_X1 U21277 ( .A1(n22632), .A2(n1503), .B1(n22388), .B2(n1439), .ZN(
        n6556) );
  OAI22_X1 U21278 ( .A1(n26674), .A2(n1501), .B1(n22412), .B2(n1437), .ZN(
        n6554) );
  OAI22_X1 U21279 ( .A1(n20674), .A2(n1499), .B1(n22137), .B2(n1435), .ZN(
        n6552) );
  OAI22_X1 U21280 ( .A1(n20642), .A2(n1497), .B1(n22182), .B2(n1433), .ZN(
        n6550) );
  OAI22_X1 U21281 ( .A1(n24975), .A2(n1495), .B1(n22231), .B2(n1431), .ZN(
        n6548) );
  OAI22_X1 U21282 ( .A1(n23802), .A2(n1493), .B1(n24366), .B2(n1429), .ZN(
        n6546) );
  OAI22_X1 U21283 ( .A1(n23753), .A2(n1491), .B1(n21721), .B2(n1427), .ZN(
        n6544) );
  OAI22_X1 U21284 ( .A1(n22656), .A2(n1489), .B1(n21737), .B2(n1425), .ZN(
        n6542) );
  OAI22_X1 U21285 ( .A1(n22624), .A2(n1487), .B1(n21753), .B2(n1423), .ZN(
        n6540) );
  OAI22_X1 U21286 ( .A1(n23965), .A2(n1485), .B1(n21769), .B2(n1421), .ZN(
        n65380) );
  OAI22_X1 U21287 ( .A1(n20666), .A2(n1483), .B1(n21662), .B2(n1419), .ZN(
        n65360) );
  OAI22_X1 U21288 ( .A1(n20633), .A2(n1481), .B1(n21670), .B2(n1417), .ZN(
        n65340) );
  OAI22_X1 U21289 ( .A1(n24983), .A2(n1479), .B1(n21678), .B2(n1415), .ZN(
        n65320) );
  OAI22_X1 U21290 ( .A1(n23778), .A2(n1477), .B1(n21686), .B2(n1413), .ZN(
        n65300) );
  OAI22_X1 U21291 ( .A1(n23825), .A2(n1475), .B1(n21726), .B2(n1411), .ZN(
        n65280) );
  OAI22_X1 U21292 ( .A1(n22648), .A2(n1473), .B1(n21742), .B2(n1409), .ZN(
        n65260) );
  OAI22_X1 U21293 ( .A1(n22616), .A2(n1471), .B1(n21758), .B2(n1407), .ZN(
        n65240) );
  OAI22_X1 U21294 ( .A1(n23963), .A2(n1469), .B1(n21774), .B2(n1405), .ZN(
        n65220) );
  OAI22_X1 U21295 ( .A1(n20658), .A2(n1467), .B1(n21694), .B2(n1403), .ZN(
        n65200) );
  OAI22_X1 U21296 ( .A1(n20625), .A2(n1465), .B1(n21702), .B2(n1401), .ZN(
        n65180) );
  OAI22_X1 U21297 ( .A1(n24979), .A2(n1463), .B1(n21710), .B2(n1399), .ZN(
        n6516) );
  OAI22_X1 U21298 ( .A1(n23758), .A2(n1461), .B1(n24365), .B2(n1397), .ZN(
        n6514) );
  OAI22_X1 U21299 ( .A1(n22672), .A2(n1459), .B1(n22153), .B2(n27883), .ZN(
        n6512) );
  INV_X1 U21300 ( .A(sram_rdata_w1[1]), .ZN(n27883) );
  OAI22_X1 U21301 ( .A1(n22640), .A2(n1457), .B1(n22198), .B2(n27881), .ZN(
        n6510) );
  INV_X1 U21302 ( .A(sram_rdata_w1[3]), .ZN(n27881) );
  OAI22_X1 U21303 ( .A1(n25237), .A2(n1455), .B1(n22243), .B2(n27879), .ZN(
        n6508) );
  INV_X1 U21304 ( .A(sram_rdata_w1[5]), .ZN(n27879) );
  OAI22_X1 U21305 ( .A1(n23751), .A2(n1453), .B1(n22278), .B2(n27877), .ZN(
        n6506) );
  INV_X1 U21306 ( .A(sram_rdata_w1[7]), .ZN(n27877) );
  OAI22_X1 U21307 ( .A1(n22664), .A2(n1451), .B1(n22003), .B2(n27875), .ZN(
        n6504) );
  INV_X1 U21308 ( .A(sram_rdata_w1[9]), .ZN(n27875) );
  OAI22_X1 U21309 ( .A1(n22632), .A2(n1449), .B1(n22039), .B2(n27873), .ZN(
        n6502) );
  INV_X1 U21310 ( .A(sram_rdata_w1[11]), .ZN(n27873) );
  OAI22_X1 U21311 ( .A1(n25226), .A2(n1447), .B1(n22075), .B2(n27871), .ZN(
        n65000) );
  INV_X1 U21312 ( .A(sram_rdata_w1[13]), .ZN(n27871) );
  OAI22_X1 U21313 ( .A1(n23835), .A2(n1445), .B1(n22111), .B2(n27869), .ZN(
        n64980) );
  INV_X1 U21314 ( .A(sram_rdata_w1[15]), .ZN(n27869) );
  OAI22_X1 U21315 ( .A1(n22656), .A2(n1443), .B1(n22007), .B2(n27867), .ZN(
        n64960) );
  INV_X1 U21316 ( .A(sram_rdata_w1[17]), .ZN(n27867) );
  OAI22_X1 U21317 ( .A1(n22624), .A2(n1441), .B1(n22043), .B2(n27865), .ZN(
        n64940) );
  INV_X1 U21318 ( .A(sram_rdata_w1[19]), .ZN(n27865) );
  OAI22_X1 U21319 ( .A1(n25227), .A2(n1439), .B1(n22079), .B2(n27863), .ZN(
        n64920) );
  INV_X1 U21320 ( .A(sram_rdata_w1[21]), .ZN(n27863) );
  OAI22_X1 U21321 ( .A1(n23795), .A2(n1437), .B1(n22115), .B2(n27861), .ZN(
        n64900) );
  INV_X1 U21322 ( .A(sram_rdata_w1[23]), .ZN(n27861) );
  OAI22_X1 U21323 ( .A1(n23801), .A2(n1435), .B1(n22343), .B2(n27859), .ZN(
        n64880) );
  INV_X1 U21324 ( .A(sram_rdata_w1[25]), .ZN(n27859) );
  OAI22_X1 U21325 ( .A1(n22669), .A2(n1433), .B1(n22367), .B2(n27857), .ZN(
        n64860) );
  INV_X1 U21326 ( .A(sram_rdata_w1[27]), .ZN(n27857) );
  OAI22_X1 U21327 ( .A1(n22637), .A2(n1431), .B1(n22391), .B2(n27855), .ZN(
        n6484) );
  INV_X1 U21328 ( .A(sram_rdata_w1[29]), .ZN(n27855) );
  OAI22_X1 U21329 ( .A1(n25356), .A2(n1429), .B1(n22415), .B2(n27853), .ZN(
        n6482) );
  INV_X1 U21330 ( .A(sram_rdata_w1[31]), .ZN(n27853) );
  OAI22_X1 U21331 ( .A1(n22648), .A2(n1427), .B1(n22157), .B2(n27851), .ZN(
        n6480) );
  INV_X1 U21332 ( .A(sram_rdata_w0[1]), .ZN(n27851) );
  OAI22_X1 U21333 ( .A1(n22616), .A2(n1425), .B1(n22203), .B2(n27849), .ZN(
        n6478) );
  INV_X1 U21334 ( .A(sram_rdata_w0[3]), .ZN(n27849) );
  OAI22_X1 U21335 ( .A1(n25240), .A2(n1423), .B1(n22235), .B2(n27847), .ZN(
        n6476) );
  INV_X1 U21336 ( .A(sram_rdata_w0[5]), .ZN(n27847) );
  OAI22_X1 U21337 ( .A1(n23771), .A2(n1421), .B1(n22267), .B2(n27845), .ZN(
        n6474) );
  INV_X1 U21338 ( .A(sram_rdata_w0[7]), .ZN(n27845) );
  OAI22_X1 U21339 ( .A1(n23777), .A2(n1419), .B1(n22337), .B2(n27843), .ZN(
        n6472) );
  INV_X1 U21340 ( .A(sram_rdata_w0[9]), .ZN(n27843) );
  OAI22_X1 U21341 ( .A1(n22660), .A2(n1417), .B1(n22361), .B2(n27841), .ZN(
        n6470) );
  INV_X1 U21342 ( .A(sram_rdata_w0[11]), .ZN(n27841) );
  OAI22_X1 U21343 ( .A1(n22628), .A2(n1415), .B1(n22385), .B2(n27839), .ZN(
        n6468) );
  INV_X1 U21344 ( .A(sram_rdata_w0[13]), .ZN(n27839) );
  OAI22_X1 U21345 ( .A1(n24974), .A2(n1413), .B1(n22409), .B2(n27837), .ZN(
        n6466) );
  INV_X1 U21346 ( .A(sram_rdata_w0[15]), .ZN(n27837) );
  OAI22_X1 U21347 ( .A1(n22668), .A2(n1411), .B1(n21989), .B2(n27835), .ZN(
        n6464) );
  INV_X1 U21348 ( .A(sram_rdata_w0[17]), .ZN(n27835) );
  OAI22_X1 U21349 ( .A1(n22636), .A2(n1409), .B1(n22025), .B2(n27833), .ZN(
        n6462) );
  INV_X1 U21350 ( .A(sram_rdata_w0[19]), .ZN(n27833) );
  OAI22_X1 U21351 ( .A1(n19100), .A2(n1407), .B1(n22061), .B2(n27831), .ZN(
        n6460) );
  INV_X1 U21352 ( .A(sram_rdata_w0[21]), .ZN(n27831) );
  OAI22_X1 U21353 ( .A1(n23745), .A2(n1405), .B1(n22097), .B2(n27829), .ZN(
        n6458) );
  INV_X1 U21354 ( .A(sram_rdata_w0[23]), .ZN(n27829) );
  OAI22_X1 U21355 ( .A1(n23747), .A2(n1403), .B1(n21719), .B2(n27827), .ZN(
        n6456) );
  INV_X1 U21356 ( .A(sram_rdata_w0[25]), .ZN(n27827) );
  OAI22_X1 U21357 ( .A1(n22652), .A2(n1401), .B1(n21735), .B2(n27825), .ZN(
        n6454) );
  INV_X1 U21358 ( .A(sram_rdata_w0[27]), .ZN(n27825) );
  OAI22_X1 U21359 ( .A1(n22620), .A2(n1399), .B1(n21751), .B2(n27823), .ZN(
        n6452) );
  INV_X1 U21360 ( .A(sram_rdata_w0[29]), .ZN(n27823) );
  OAI22_X1 U21361 ( .A1(n20770), .A2(n1397), .B1(n21767), .B2(n27821), .ZN(
        n6450) );
  INV_X1 U21362 ( .A(sram_rdata_w0[31]), .ZN(n27821) );
  OAI22_X1 U21363 ( .A1(n22660), .A2(n14247), .B1(n22144), .B2(n1388), .ZN(
        n74090) );
  OAI22_X1 U21364 ( .A1(n22628), .A2(n14261), .B1(n22190), .B2(n1386), .ZN(
        n74070) );
  OAI22_X1 U21365 ( .A1(n20762), .A2(n14275), .B1(n22225), .B2(n1384), .ZN(
        n74050) );
  OAI22_X1 U21366 ( .A1(n23830), .A2(n14289), .B1(n22260), .B2(n1382), .ZN(
        n74030) );
  OAI22_X1 U21367 ( .A1(n23819), .A2(n1388), .B1(n22332), .B2(n1380), .ZN(
        n74010) );
  OAI22_X1 U21368 ( .A1(n22644), .A2(n1386), .B1(n22356), .B2(n1378), .ZN(
        n73990) );
  OAI22_X1 U21369 ( .A1(n22612), .A2(n1384), .B1(n22380), .B2(n1376), .ZN(
        n73970) );
  OAI22_X1 U21370 ( .A1(n20758), .A2(n1382), .B1(n22404), .B2(n1374), .ZN(
        n73950) );
  OAI22_X1 U21371 ( .A1(n22652), .A2(n1380), .B1(n21997), .B2(n1372), .ZN(
        n73930) );
  OAI22_X1 U21372 ( .A1(n22620), .A2(n1378), .B1(n22033), .B2(n1370), .ZN(
        n7391) );
  OAI22_X1 U21373 ( .A1(n20751), .A2(n1376), .B1(n22069), .B2(n1368), .ZN(
        n7389) );
  OAI22_X1 U21374 ( .A1(n23812), .A2(n1374), .B1(n22105), .B2(n1366), .ZN(
        n7387) );
  OAI22_X1 U21375 ( .A1(n23796), .A2(n1372), .B1(n22325), .B2(n1364), .ZN(
        n7385) );
  OAI22_X1 U21376 ( .A1(n20681), .A2(n1370), .B1(n22349), .B2(n1362), .ZN(
        n7383) );
  OAI22_X1 U21377 ( .A1(n20649), .A2(n1368), .B1(n22373), .B2(n1360), .ZN(
        n7381) );
  OAI22_X1 U21378 ( .A1(n19065), .A2(n1366), .B1(n22397), .B2(n1358), .ZN(
        n7379) );
  OAI22_X1 U21379 ( .A1(n22645), .A2(n1364), .B1(n22121), .B2(n1356), .ZN(
        n7377) );
  OAI22_X1 U21380 ( .A1(n22613), .A2(n1362), .B1(n22164), .B2(n1354), .ZN(
        n73750) );
  OAI22_X1 U21381 ( .A1(n24980), .A2(n1360), .B1(n22217), .B2(n1352), .ZN(
        n73730) );
  OAI22_X1 U21382 ( .A1(n23788), .A2(n1358), .B1(n22253), .B2(n1350), .ZN(
        n73710) );
  OAI22_X1 U21383 ( .A1(n25031), .A2(n1356), .B1(n22127), .B2(n1348), .ZN(
        n73690) );
  OAI22_X1 U21384 ( .A1(n25048), .A2(n1354), .B1(n22171), .B2(n1346), .ZN(
        n73670) );
  OAI22_X1 U21385 ( .A1(n19060), .A2(n1352), .B1(n22211), .B2(n1344), .ZN(
        n73650) );
  OAI22_X1 U21386 ( .A1(n23824), .A2(n1350), .B1(n22247), .B2(n1342), .ZN(
        n73630) );
  OAI22_X1 U21387 ( .A1(n25038), .A2(n1348), .B1(n21977), .B2(n27948), .ZN(
        n73610) );
  INV_X1 U21388 ( .A(sram_rdata_d1[0]), .ZN(n27948) );
  OAI22_X1 U21389 ( .A1(n25054), .A2(n1346), .B1(n22013), .B2(n27946), .ZN(
        n7359) );
  INV_X1 U21390 ( .A(sram_rdata_d1[2]), .ZN(n27946) );
  OAI22_X1 U21391 ( .A1(n25354), .A2(n1344), .B1(n22049), .B2(n27944), .ZN(
        n7357) );
  INV_X1 U21392 ( .A(sram_rdata_d1[4]), .ZN(n27944) );
  OAI22_X1 U21393 ( .A1(n23805), .A2(n1342), .B1(n22085), .B2(n27942), .ZN(
        n7355) );
  INV_X1 U21394 ( .A(sram_rdata_d1[6]), .ZN(n27942) );
  OAI22_X1 U21395 ( .A1(n25042), .A2(n14567), .B1(n21984), .B2(n1332), .ZN(
        n7345) );
  OAI22_X1 U21396 ( .A1(n25058), .A2(n14581), .B1(n22020), .B2(n1330), .ZN(
        n7343) );
  OAI22_X1 U21397 ( .A1(n25230), .A2(n14595), .B1(n22056), .B2(n1328), .ZN(
        n7341) );
  OAI22_X1 U21398 ( .A1(n23782), .A2(n14609), .B1(n22092), .B2(n1326), .ZN(
        n7339) );
  OAI22_X1 U21399 ( .A1(n23772), .A2(n1332), .B1(n21712), .B2(n1324), .ZN(
        n7337) );
  OAI22_X1 U21400 ( .A1(n20673), .A2(n1330), .B1(n21728), .B2(n1322), .ZN(
        n7335) );
  OAI22_X1 U21401 ( .A1(n20641), .A2(n1328), .B1(n21744), .B2(n1320), .ZN(
        n7333) );
  OAI22_X1 U21402 ( .A1(n25361), .A2(n1326), .B1(n21760), .B2(n1318), .ZN(
        n7331) );
  OAI22_X1 U21403 ( .A1(n24843), .A2(n1324), .B1(n21680), .B2(n1316), .ZN(
        n7329) );
  OAI22_X1 U21404 ( .A1(n24826), .A2(n1322), .B1(n21688), .B2(n1314), .ZN(
        n7327) );
  OAI22_X1 U21405 ( .A1(n25358), .A2(n1320), .B1(n21696), .B2(n1312), .ZN(
        n7325) );
  OAI22_X1 U21406 ( .A1(n23764), .A2(n1318), .B1(n21704), .B2(n1310), .ZN(
        n73230) );
  OAI22_X1 U21407 ( .A1(n23765), .A2(n1316), .B1(n21716), .B2(n1308), .ZN(
        n73210) );
  OAI22_X1 U21408 ( .A1(n20663), .A2(n1314), .B1(n21732), .B2(n1306), .ZN(
        n73190) );
  OAI22_X1 U21409 ( .A1(n20630), .A2(n1312), .B1(n21748), .B2(n1304), .ZN(
        n73170) );
  OAI22_X1 U21410 ( .A1(n23962), .A2(n1310), .B1(n21764), .B2(n1302), .ZN(
        n73150) );
  OAI22_X1 U21411 ( .A1(n20680), .A2(n1308), .B1(n22266), .B2(n1300), .ZN(
        n73130) );
  OAI22_X1 U21412 ( .A1(n20648), .A2(n1306), .B1(n21656), .B2(n1298), .ZN(
        n73110) );
  OAI22_X1 U21413 ( .A1(n24131), .A2(n1304), .B1(n21664), .B2(n1296), .ZN(
        n73090) );
  OAI22_X1 U21414 ( .A1(n23818), .A2(n1302), .B1(n21672), .B2(n1294), .ZN(
        n73070) );
  OAI22_X1 U21415 ( .A1(n23836), .A2(n1300), .B1(n22329), .B2(n1292), .ZN(
        n73050) );
  OAI22_X1 U21416 ( .A1(n20655), .A2(n1298), .B1(n22353), .B2(n1290), .ZN(
        n7303) );
  OAI22_X1 U21417 ( .A1(n20622), .A2(n1296), .B1(n22377), .B2(n1288), .ZN(
        n7301) );
  OAI22_X1 U21418 ( .A1(n24119), .A2(n1294), .B1(n22401), .B2(n1286), .ZN(
        n7299) );
  OAI22_X1 U21419 ( .A1(n20672), .A2(n1292), .B1(n22143), .B2(n27940), .ZN(
        n7297) );
  INV_X1 U21420 ( .A(sram_rdata_d1[8]), .ZN(n27940) );
  OAI22_X1 U21421 ( .A1(n20639), .A2(n1290), .B1(n22189), .B2(n27938), .ZN(
        n7295) );
  INV_X1 U21422 ( .A(sram_rdata_d1[10]), .ZN(n27938) );
  OAI22_X1 U21423 ( .A1(n24108), .A2(n1288), .B1(n22224), .B2(n27936), .ZN(
        n7293) );
  INV_X1 U21424 ( .A(sram_rdata_d1[12]), .ZN(n27936) );
  OAI22_X1 U21425 ( .A1(n23800), .A2(n1286), .B1(n22259), .B2(n27934), .ZN(
        n7291) );
  INV_X1 U21426 ( .A(sram_rdata_d1[14]), .ZN(n27934) );
  OAI22_X1 U21427 ( .A1(n24844), .A2(n14887), .B1(n26429), .B2(n1276), .ZN(
        n72810) );
  OAI22_X1 U21428 ( .A1(n24827), .A2(n14901), .B1(n26437), .B2(n1274), .ZN(
        n72790) );
  OAI22_X1 U21429 ( .A1(n24125), .A2(n14915), .B1(n26447), .B2(n1272), .ZN(
        n72770) );
  OAI22_X1 U21430 ( .A1(n23776), .A2(n14929), .B1(n26453), .B2(n1270), .ZN(
        n72750) );
  OAI22_X1 U21431 ( .A1(n20656), .A2(n1276), .B1(n21995), .B2(n1268), .ZN(
        n72730) );
  OAI22_X1 U21432 ( .A1(n20623), .A2(n1274), .B1(n22031), .B2(n1266), .ZN(
        n72710) );
  OAI22_X1 U21433 ( .A1(n24137), .A2(n1272), .B1(n22067), .B2(n1264), .ZN(
        n7269) );
  OAI22_X1 U21434 ( .A1(n22556), .A2(n1270), .B1(n22103), .B2(n1262), .ZN(
        n72670) );
  OAI22_X1 U21435 ( .A1(n22671), .A2(n1268), .B1(n26405), .B2(n1260), .ZN(
        n7265) );
  OAI22_X1 U21436 ( .A1(n22639), .A2(n1266), .B1(n26411), .B2(n1258), .ZN(
        n7263) );
  OAI22_X1 U21437 ( .A1(n24113), .A2(n1264), .B1(n26417), .B2(n1256), .ZN(
        n7261) );
  OAI22_X1 U21438 ( .A1(n22608), .A2(n1262), .B1(n26423), .B2(n1254), .ZN(
        n7259) );
  OAI22_X1 U21439 ( .A1(n23811), .A2(n1260), .B1(n22323), .B2(n1252), .ZN(
        n7257) );
  OAI22_X1 U21440 ( .A1(n25035), .A2(n1258), .B1(n22347), .B2(n1250), .ZN(
        n7255) );
  OAI22_X1 U21441 ( .A1(n25051), .A2(n1256), .B1(n22371), .B2(n1248), .ZN(
        n7253) );
  OAI22_X1 U21442 ( .A1(n19096), .A2(n1254), .B1(n22395), .B2(n1246), .ZN(
        n7251) );
  OAI22_X1 U21443 ( .A1(n22663), .A2(n1252), .B1(n264301), .B2(n1244), .ZN(
        n7249) );
  OAI22_X1 U21444 ( .A1(n22631), .A2(n1250), .B1(n70), .B2(n1242), .ZN(n7247)
         );
  OAI22_X1 U21445 ( .A1(n25356), .A2(n1248), .B1(n26446), .B2(n1240), .ZN(
        n7245) );
  OAI22_X1 U21446 ( .A1(n23794), .A2(n1246), .B1(n26452), .B2(n1238), .ZN(
        n7243) );
  OAI22_X1 U21447 ( .A1(n23787), .A2(n1244), .B1(n26209), .B2(n1236), .ZN(
        n72410) );
  OAI22_X1 U21448 ( .A1(n25036), .A2(n1242), .B1(n26217), .B2(n1234), .ZN(
        n72390) );
  OAI22_X1 U21449 ( .A1(n25052), .A2(n1240), .B1(n26225), .B2(n1232), .ZN(
        n72370) );
  OAI22_X1 U21450 ( .A1(n19101), .A2(n1238), .B1(n26233), .B2(n1230), .ZN(
        n72350) );
  OAI22_X1 U21451 ( .A1(n22654), .A2(n1236), .B1(n26406), .B2(n27932), .ZN(
        n72330) );
  INV_X1 U21452 ( .A(sram_rdata_d1[16]), .ZN(n27932) );
  OAI22_X1 U21453 ( .A1(n22622), .A2(n1234), .B1(n26412), .B2(n27930), .ZN(
        n72310) );
  INV_X1 U21454 ( .A(sram_rdata_d1[18]), .ZN(n27930) );
  OAI22_X1 U21455 ( .A1(n19065), .A2(n1232), .B1(n26418), .B2(n27928), .ZN(
        n72290) );
  INV_X1 U21456 ( .A(sram_rdata_d1[20]), .ZN(n27928) );
  OAI22_X1 U21457 ( .A1(n23770), .A2(n1230), .B1(n26424), .B2(n27926), .ZN(
        n72270) );
  INV_X1 U21458 ( .A(sram_rdata_d1[22]), .ZN(n27926) );
  OAI22_X1 U21459 ( .A1(n23757), .A2(n15207), .B1(n26211), .B2(n1220), .ZN(
        n7217) );
  OAI22_X1 U21460 ( .A1(n25043), .A2(n15221), .B1(n26219), .B2(n1218), .ZN(
        n7215) );
  OAI22_X1 U21461 ( .A1(n25059), .A2(n15235), .B1(n26227), .B2(n1216), .ZN(
        n7213) );
  OAI22_X1 U21462 ( .A1(n22674), .A2(n15249), .B1(n26235), .B2(n1214), .ZN(
        n7211) );
  OAI22_X1 U21463 ( .A1(n22647), .A2(n1220), .B1(n26177), .B2(n1212), .ZN(
        n7209) );
  OAI22_X1 U21464 ( .A1(n22615), .A2(n1218), .B1(n26181), .B2(n1210), .ZN(
        n7207) );
  OAI22_X1 U21465 ( .A1(n25224), .A2(n1216), .B1(n26185), .B2(n1208), .ZN(
        n7205) );
  OAI22_X1 U21466 ( .A1(n22552), .A2(n1214), .B1(n26189), .B2(n1206), .ZN(
        n72030) );
  OAI22_X1 U21467 ( .A1(n22667), .A2(n1212), .B1(n22147), .B2(n1204), .ZN(
        n72010) );
  OAI22_X1 U21468 ( .A1(n22635), .A2(n1210), .B1(n69), .B2(n1202), .ZN(n71990)
         );
  OAI22_X1 U21469 ( .A1(n25353), .A2(n1208), .B1(n26448), .B2(n1200), .ZN(
        n71970) );
  OAI22_X1 U21470 ( .A1(n22604), .A2(n1206), .B1(n26454), .B2(n1198), .ZN(
        n71950) );
  OAI22_X1 U21471 ( .A1(n22659), .A2(n1204), .B1(n26161), .B2(n1196), .ZN(
        n71930) );
  OAI22_X1 U21472 ( .A1(n22627), .A2(n1202), .B1(n26165), .B2(n1194), .ZN(
        n71910) );
  OAI22_X1 U21473 ( .A1(n24133), .A2(n1200), .B1(n26169), .B2(n1192), .ZN(
        n71890) );
  OAI22_X1 U21474 ( .A1(n22592), .A2(n1198), .B1(n26173), .B2(n1190), .ZN(
        n7187) );
  OAI22_X1 U21475 ( .A1(n22651), .A2(n1196), .B1(n26408), .B2(n1188), .ZN(
        n7185) );
  OAI22_X1 U21476 ( .A1(n22619), .A2(n1194), .B1(n26414), .B2(n1186), .ZN(
        n7183) );
  OAI22_X1 U21477 ( .A1(n24109), .A2(n1192), .B1(n264201), .B2(n1184), .ZN(
        n7181) );
  OAI22_X1 U21478 ( .A1(n22576), .A2(n1190), .B1(n26426), .B2(n1182), .ZN(
        n7179) );
  OAI22_X1 U21479 ( .A1(n23829), .A2(n1188), .B1(n26481), .B2(n1180), .ZN(
        n7177) );
  OAI22_X1 U21480 ( .A1(n25044), .A2(n1186), .B1(n26485), .B2(n1178), .ZN(
        n7175) );
  OAI22_X1 U21481 ( .A1(n25061), .A2(n1184), .B1(n26489), .B2(n1176), .ZN(
        n7173) );
  OAI22_X1 U21482 ( .A1(n24121), .A2(n1182), .B1(n26493), .B2(n1174), .ZN(
        n7171) );
  OAI22_X1 U21483 ( .A1(n22643), .A2(n1180), .B1(n22125), .B2(n27924), .ZN(
        n7169) );
  INV_X1 U21484 ( .A(sram_rdata_d1[24]), .ZN(n27924) );
  OAI22_X1 U21485 ( .A1(n22611), .A2(n1178), .B1(n22169), .B2(n27922), .ZN(
        n7167) );
  INV_X1 U21486 ( .A(sram_rdata_d1[26]), .ZN(n27922) );
  OAI22_X1 U21487 ( .A1(n24127), .A2(n1176), .B1(n22221), .B2(n27920), .ZN(
        n7165) );
  INV_X1 U21488 ( .A(sram_rdata_d1[28]), .ZN(n27920) );
  OAI22_X1 U21489 ( .A1(n22548), .A2(n1174), .B1(n22256), .B2(n27918), .ZN(
        n7163) );
  INV_X1 U21490 ( .A(sram_rdata_d1[30]), .ZN(n27918) );
  OAI22_X1 U21491 ( .A1(n23806), .A2(n15527), .B1(n264801), .B2(n1164), .ZN(
        n7153) );
  OAI22_X1 U21492 ( .A1(n22670), .A2(n15541), .B1(n26484), .B2(n1162), .ZN(
        n7151) );
  OAI22_X1 U21493 ( .A1(n22638), .A2(n15555), .B1(n26488), .B2(n1160), .ZN(
        n71490) );
  OAI22_X1 U21494 ( .A1(n24139), .A2(n15569), .B1(n26492), .B2(n1158), .ZN(
        n71470) );
  OAI22_X1 U21495 ( .A1(n20818), .A2(n1164), .B1(n21982), .B2(n1156), .ZN(
        n71450) );
  OAI22_X1 U21496 ( .A1(n20842), .A2(n1162), .B1(n22018), .B2(n1154), .ZN(
        n71430) );
  OAI22_X1 U21497 ( .A1(n19093), .A2(n1160), .B1(n22054), .B2(n1152), .ZN(
        n71410) );
  OAI22_X1 U21498 ( .A1(n22600), .A2(n1158), .B1(n22090), .B2(n1150), .ZN(
        n71390) );
  OAI22_X1 U21499 ( .A1(n23781), .A2(n1156), .B1(n26208), .B2(n1148), .ZN(
        n71370) );
  OAI22_X1 U21500 ( .A1(n22662), .A2(n1154), .B1(n26216), .B2(n1146), .ZN(
        n71350) );
  OAI22_X1 U21501 ( .A1(n22630), .A2(n1152), .B1(n26224), .B2(n1144), .ZN(
        n71330) );
  OAI22_X1 U21502 ( .A1(n24115), .A2(n1150), .B1(n26232), .B2(n1142), .ZN(
        n71310) );
  OAI22_X1 U21503 ( .A1(n20820), .A2(n1148), .B1(n22133), .B2(n1140), .ZN(
        n7129) );
  OAI22_X1 U21504 ( .A1(n20844), .A2(n1146), .B1(n22177), .B2(n1138), .ZN(
        n7127) );
  OAI22_X1 U21505 ( .A1(n19099), .A2(n1144), .B1(n22216), .B2(n1136), .ZN(
        n7125) );
  OAI22_X1 U21506 ( .A1(n22588), .A2(n1142), .B1(n22252), .B2(n1134), .ZN(
        n7123) );
  OAI22_X1 U21507 ( .A1(n20669), .A2(n1140), .B1(n26176), .B2(n1132), .ZN(
        n7121) );
  OAI22_X1 U21508 ( .A1(n20636), .A2(n1138), .B1(n26180), .B2(n1130), .ZN(
        n7119) );
  OAI22_X1 U21509 ( .A1(n25359), .A2(n1136), .B1(n26184), .B2(n1128), .ZN(
        n7117) );
  OAI22_X1 U21510 ( .A1(n22572), .A2(n1134), .B1(n26188), .B2(n1126), .ZN(
        n7115) );
  OAI22_X1 U21511 ( .A1(n20832), .A2(n1132), .B1(n21988), .B2(n1124), .ZN(
        n7113) );
  OAI22_X1 U21512 ( .A1(n20857), .A2(n1130), .B1(n22024), .B2(n1122), .ZN(
        n71110) );
  OAI22_X1 U21513 ( .A1(n25355), .A2(n1128), .B1(n22060), .B2(n1120), .ZN(
        n71090) );
  OAI22_X1 U21514 ( .A1(n22560), .A2(n1126), .B1(n22096), .B2(n1118), .ZN(
        n71070) );
  OAI22_X1 U21515 ( .A1(n25031), .A2(n1124), .B1(n26160), .B2(n27916), .ZN(
        n71050) );
  INV_X1 U21516 ( .A(sram_rdata_d0[0]), .ZN(n27916) );
  OAI22_X1 U21517 ( .A1(n25048), .A2(n1122), .B1(n26164), .B2(n27914), .ZN(
        n71030) );
  INV_X1 U21518 ( .A(sram_rdata_d0[2]), .ZN(n27914) );
  OAI22_X1 U21519 ( .A1(n25225), .A2(n1120), .B1(n26168), .B2(n27912), .ZN(
        n71010) );
  INV_X1 U21520 ( .A(sram_rdata_d0[4]), .ZN(n27912) );
  OAI22_X1 U21521 ( .A1(n22596), .A2(n1118), .B1(n26172), .B2(n27910), .ZN(
        n70990) );
  INV_X1 U21522 ( .A(sram_rdata_d0[6]), .ZN(n27910) );
  OAI22_X1 U21523 ( .A1(n23752), .A2(n15847), .B1(n26210), .B2(n1108), .ZN(
        n7089) );
  OAI22_X1 U21524 ( .A1(n22654), .A2(n15861), .B1(n26218), .B2(n1106), .ZN(
        n7087) );
  OAI22_X1 U21525 ( .A1(n22622), .A2(n15875), .B1(n26226), .B2(n1104), .ZN(
        n7085) );
  OAI22_X1 U21526 ( .A1(n23966), .A2(n15889), .B1(n26234), .B2(n1102), .ZN(
        n7083) );
  OAI22_X1 U21527 ( .A1(n20823), .A2(n1108), .B1(n22147), .B2(n1100), .ZN(
        n7081) );
  OAI22_X1 U21528 ( .A1(n20847), .A2(n1106), .B1(n22193), .B2(n1098), .ZN(
        n7079) );
  OAI22_X1 U21529 ( .A1(n25234), .A2(n1104), .B1(n22228), .B2(n1096), .ZN(
        n7077) );
  OAI22_X1 U21530 ( .A1(n22584), .A2(n1102), .B1(n22263), .B2(n1094), .ZN(
        n7075) );
  OAI22_X1 U21531 ( .A1(n23823), .A2(n1100), .B1(n22334), .B2(n1092), .ZN(
        n7073) );
  OAI22_X1 U21532 ( .A1(n22646), .A2(n1098), .B1(n22358), .B2(n1090), .ZN(
        n7071) );
  OAI22_X1 U21533 ( .A1(n22614), .A2(n1096), .B1(n22382), .B2(n1088), .ZN(
        n7069) );
  OAI22_X1 U21534 ( .A1(n24981), .A2(n1094), .B1(n22406), .B2(n1086), .ZN(
        n70670) );
  OAI22_X1 U21535 ( .A1(n20825), .A2(n1092), .B1(n22000), .B2(n1084), .ZN(
        n70650) );
  OAI22_X1 U21536 ( .A1(n20849), .A2(n1090), .B1(n22036), .B2(n1082), .ZN(
        n70630) );
  OAI22_X1 U21537 ( .A1(n24977), .A2(n1088), .B1(n22072), .B2(n1080), .ZN(
        n70610) );
  OAI22_X1 U21538 ( .A1(n22568), .A2(n1086), .B1(n22108), .B2(n1078), .ZN(
        n70590) );
  OAI22_X1 U21539 ( .A1(n23800), .A2(n1084), .B1(n22328), .B2(n1076), .ZN(
        n70570) );
  OAI22_X1 U21540 ( .A1(n22666), .A2(n1082), .B1(n22352), .B2(n1074), .ZN(
        n70550) );
  OAI22_X1 U21541 ( .A1(n22634), .A2(n1080), .B1(n22376), .B2(n1072), .ZN(
        n70530) );
  OAI22_X1 U21542 ( .A1(n20757), .A2(n1078), .B1(n22400), .B2(n1070), .ZN(
        n70510) );
  OAI22_X1 U21543 ( .A1(n20835), .A2(n1076), .B1(n22123), .B2(n1068), .ZN(
        n70490) );
  OAI22_X1 U21544 ( .A1(n20860), .A2(n1074), .B1(n22167), .B2(n1066), .ZN(
        n7047) );
  OAI22_X1 U21545 ( .A1(n20778), .A2(n1072), .B1(n22219), .B2(n1064), .ZN(
        n7045) );
  OAI22_X1 U21546 ( .A1(n22554), .A2(n1070), .B1(n22255), .B2(n1062), .ZN(
        n7043) );
  OAI22_X1 U21547 ( .A1(n23933), .A2(n1068), .B1(n22129), .B2(n27908), .ZN(
        n7041) );
  INV_X1 U21548 ( .A(sram_rdata_d0[8]), .ZN(n27908) );
  OAI22_X1 U21549 ( .A1(n23885), .A2(n1066), .B1(n22173), .B2(n27906), .ZN(
        n7039) );
  INV_X1 U21550 ( .A(sram_rdata_d0[10]), .ZN(n27906) );
  OAI22_X1 U21551 ( .A1(n20764), .A2(n1064), .B1(n22213), .B2(n27904), .ZN(
        n7037) );
  INV_X1 U21552 ( .A(sram_rdata_d0[12]), .ZN(n27904) );
  OAI22_X1 U21553 ( .A1(n22606), .A2(n1062), .B1(n22249), .B2(n27902), .ZN(
        n7035) );
  INV_X1 U21554 ( .A(sram_rdata_d0[14]), .ZN(n27902) );
  OAI22_X1 U21555 ( .A1(n23921), .A2(n16167), .B1(n21979), .B2(n1052), .ZN(
        n70250) );
  OAI22_X1 U21556 ( .A1(n23873), .A2(n16181), .B1(n22015), .B2(n1050), .ZN(
        n70230) );
  OAI22_X1 U21557 ( .A1(n25351), .A2(n16195), .B1(n22051), .B2(n1048), .ZN(
        n70210) );
  OAI22_X1 U21558 ( .A1(n22580), .A2(n16209), .B1(n22087), .B2(n1046), .ZN(
        n70190) );
  OAI22_X1 U21559 ( .A1(n23910), .A2(n1052), .B1(n21986), .B2(n1044), .ZN(
        n70170) );
  OAI22_X1 U21560 ( .A1(n23862), .A2(n1050), .B1(n22022), .B2(n1042), .ZN(
        n70150) );
  OAI22_X1 U21561 ( .A1(n20773), .A2(n1048), .B1(n22058), .B2(n1040), .ZN(
        n7013) );
  OAI22_X1 U21562 ( .A1(n22564), .A2(n1046), .B1(n22094), .B2(n1038), .ZN(
        n7011) );
  OAI22_X1 U21563 ( .A1(n23775), .A2(n1044), .B1(n21713), .B2(n1036), .ZN(
        n7009) );
  OAI22_X1 U21564 ( .A1(n22658), .A2(n1042), .B1(n21729), .B2(n1034), .ZN(
        n7007) );
  OAI22_X1 U21565 ( .A1(n22626), .A2(n1040), .B1(n21745), .B2(n1032), .ZN(
        n7005) );
  OAI22_X1 U21566 ( .A1(n17084), .A2(n1038), .B1(n21761), .B2(n1030), .ZN(
        n7003) );
  OAI22_X1 U21567 ( .A1(n23898), .A2(n1036), .B1(n21681), .B2(n1028), .ZN(
        n7001) );
  OAI22_X1 U21568 ( .A1(n23850), .A2(n1034), .B1(n21689), .B2(n1026), .ZN(
        n6999) );
  OAI22_X1 U21569 ( .A1(n25352), .A2(n1032), .B1(n21697), .B2(n1024), .ZN(
        n6997) );
  OAI22_X1 U21570 ( .A1(n22550), .A2(n1030), .B1(n21705), .B2(n1022), .ZN(
        n6995) );
  OAI22_X1 U21571 ( .A1(n23746), .A2(n1028), .B1(n21718), .B2(n1020), .ZN(
        n6993) );
  OAI22_X1 U21572 ( .A1(n22650), .A2(n1026), .B1(n21734), .B2(n1018), .ZN(
        n6991) );
  OAI22_X1 U21573 ( .A1(n22618), .A2(n1024), .B1(n21750), .B2(n1016), .ZN(
        n6989) );
  OAI22_X1 U21574 ( .A1(n23964), .A2(n1022), .B1(n21766), .B2(n1014), .ZN(
        n6987) );
  OAI22_X1 U21575 ( .A1(n23928), .A2(n1020), .B1(n21649), .B2(n1012), .ZN(
        n6985) );
  OAI22_X1 U21576 ( .A1(n23880), .A2(n1018), .B1(n21657), .B2(n1010), .ZN(
        n6983) );
  OAI22_X1 U21577 ( .A1(n19093), .A2(n1016), .B1(n21665), .B2(n1008), .ZN(
        n6981) );
  OAI22_X1 U21578 ( .A1(n22602), .A2(n1014), .B1(n21673), .B2(n1006), .ZN(
        n6979) );
  OAI22_X1 U21579 ( .A1(n23817), .A2(n1012), .B1(n22331), .B2(n27900), .ZN(
        n6977) );
  INV_X1 U21580 ( .A(sram_rdata_d0[16]), .ZN(n27900) );
  OAI22_X1 U21581 ( .A1(n22642), .A2(n1010), .B1(n22355), .B2(n27898), .ZN(
        n69750) );
  INV_X1 U21582 ( .A(sram_rdata_d0[18]), .ZN(n27898) );
  OAI22_X1 U21583 ( .A1(n22610), .A2(n1008), .B1(n22379), .B2(n27896), .ZN(
        n69730) );
  INV_X1 U21584 ( .A(sram_rdata_d0[20]), .ZN(n27896) );
  OAI22_X1 U21585 ( .A1(n25358), .A2(n1006), .B1(n22403), .B2(n27894), .ZN(
        n69710) );
  INV_X1 U21586 ( .A(sram_rdata_d0[22]), .ZN(n27894) );
  OAI22_X1 U21587 ( .A1(n23916), .A2(n16487), .B1(n22144), .B2(n996), .ZN(
        n69610) );
  OAI22_X1 U21588 ( .A1(n23868), .A2(n16501), .B1(n22190), .B2(n994), .ZN(
        n69590) );
  OAI22_X1 U21589 ( .A1(n19099), .A2(n16515), .B1(n22226), .B2(n992), .ZN(
        n69570) );
  OAI22_X1 U21590 ( .A1(n22590), .A2(n16529), .B1(n22261), .B2(n990), .ZN(
        n6955) );
  OAI22_X1 U21591 ( .A1(n23903), .A2(n996), .B1(n22122), .B2(n988), .ZN(n6953)
         );
  OAI22_X1 U21592 ( .A1(n23855), .A2(n994), .B1(n22165), .B2(n986), .ZN(n6951)
         );
  OAI22_X1 U21593 ( .A1(n20763), .A2(n992), .B1(n22218), .B2(n984), .ZN(n6949)
         );
  OAI22_X1 U21594 ( .A1(n22574), .A2(n990), .B1(n22254), .B2(n982), .ZN(n6947)
         );
  OAI22_X1 U21595 ( .A1(n23892), .A2(n988), .B1(n21997), .B2(n980), .ZN(n6945)
         );
  OAI22_X1 U21596 ( .A1(n23844), .A2(n986), .B1(n22033), .B2(n978), .ZN(n6943)
         );
  OAI22_X1 U21597 ( .A1(n20755), .A2(n984), .B1(n22069), .B2(n976), .ZN(n6941)
         );
  OAI22_X1 U21598 ( .A1(n22598), .A2(n982), .B1(n22105), .B2(n974), .ZN(n6939)
         );
  OAI22_X1 U21599 ( .A1(n25035), .A2(n980), .B1(n21977), .B2(n972), .ZN(n69370) );
  OAI22_X1 U21600 ( .A1(n25051), .A2(n978), .B1(n22014), .B2(n970), .ZN(n69350) );
  OAI22_X1 U21601 ( .A1(n24982), .A2(n976), .B1(n22050), .B2(n968), .ZN(n69330) );
  OAI22_X1 U21602 ( .A1(n22586), .A2(n974), .B1(n22086), .B2(n966), .ZN(n69310) );
  OAI22_X1 U21603 ( .A1(n23793), .A2(n972), .B1(n22326), .B2(n964), .ZN(n69290) );
  OAI22_X1 U21604 ( .A1(n24852), .A2(n970), .B1(n22350), .B2(n962), .ZN(n69270) );
  OAI22_X1 U21605 ( .A1(n24836), .A2(n968), .B1(n22374), .B2(n960), .ZN(n69250) );
  OAI22_X1 U21606 ( .A1(n20750), .A2(n966), .B1(n22398), .B2(n958), .ZN(n69230) );
  OAI22_X1 U21607 ( .A1(n25036), .A2(n964), .B1(n22127), .B2(n956), .ZN(n6921)
         );
  OAI22_X1 U21608 ( .A1(n25052), .A2(n962), .B1(n22171), .B2(n954), .ZN(n6919)
         );
  OAI22_X1 U21609 ( .A1(n20759), .A2(n960), .B1(n22212), .B2(n952), .ZN(n6917)
         );
  OAI22_X1 U21610 ( .A1(n22570), .A2(n958), .B1(n22248), .B2(n950), .ZN(n6915)
         );
  OAI22_X1 U21611 ( .A1(n23769), .A2(n956), .B1(n21711), .B2(n27892), .ZN(
        n6913) );
  INV_X1 U21612 ( .A(sram_rdata_d0[24]), .ZN(n27892) );
  OAI22_X1 U21613 ( .A1(n24848), .A2(n954), .B1(n21727), .B2(n27890), .ZN(
        n6911) );
  INV_X1 U21614 ( .A(sram_rdata_d0[26]), .ZN(n27890) );
  OAI22_X1 U21615 ( .A1(n24831), .A2(n952), .B1(n21743), .B2(n27888), .ZN(
        n6909) );
  INV_X1 U21616 ( .A(sram_rdata_d0[28]), .ZN(n27888) );
  OAI22_X1 U21617 ( .A1(n20766), .A2(n950), .B1(n21759), .B2(n27886), .ZN(
        n6907) );
  INV_X1 U21618 ( .A(sram_rdata_d0[30]), .ZN(n27886) );
  OAI22_X1 U21619 ( .A1(n25043), .A2(n11869), .B1(n22019), .B2(n1778), .ZN(
        n6895) );
  OAI22_X1 U21620 ( .A1(n25059), .A2(n11883), .B1(n22055), .B2(n1776), .ZN(
        n68930) );
  OAI22_X1 U21621 ( .A1(n25237), .A2(n11897), .B1(n22091), .B2(n1774), .ZN(
        n68910) );
  OAI22_X1 U21622 ( .A1(n22597), .A2(n11911), .B1(n21715), .B2(n1772), .ZN(
        n68890) );
  OAI22_X1 U21623 ( .A1(n25040), .A2(n11925), .B1(n21731), .B2(n1770), .ZN(
        n68870) );
  OAI22_X1 U21624 ( .A1(n25056), .A2(n11939), .B1(n21747), .B2(n1768), .ZN(
        n68850) );
  OAI22_X1 U21625 ( .A1(n25357), .A2(n11953), .B1(n21763), .B2(n1766), .ZN(
        n68830) );
  OAI22_X1 U21626 ( .A1(n22554), .A2(n11967), .B1(n21679), .B2(n1764), .ZN(
        n68810) );
  OAI22_X1 U21627 ( .A1(n20832), .A2(n11981), .B1(n21687), .B2(n1762), .ZN(
        n68790) );
  OAI22_X1 U21628 ( .A1(n20857), .A2(n11995), .B1(n21695), .B2(n1760), .ZN(
        n68770) );
  OAI22_X1 U21629 ( .A1(n25232), .A2(n12009), .B1(n21703), .B2(n1758), .ZN(
        n68750) );
  OAI22_X1 U21630 ( .A1(n22568), .A2(n12023), .B1(n22142), .B2(n1756), .ZN(
        n6873) );
  OAI22_X1 U21631 ( .A1(n20819), .A2(n12037), .B1(n22188), .B2(n1754), .ZN(
        n6871) );
  OAI22_X1 U21632 ( .A1(n20843), .A2(n12051), .B1(n22223), .B2(n1752), .ZN(
        n6869) );
  OAI22_X1 U21633 ( .A1(n25364), .A2(n12065), .B1(n22258), .B2(n1750), .ZN(
        n6867) );
  OAI22_X1 U21634 ( .A1(n22584), .A2(n12079), .B1(n21983), .B2(n1748), .ZN(
        n6865) );
  OAI22_X1 U21635 ( .A1(n20821), .A2(n12093), .B1(n21655), .B2(n1746), .ZN(
        n6863) );
  OAI22_X1 U21636 ( .A1(n20845), .A2(n12107), .B1(n21663), .B2(n1744), .ZN(
        n6861) );
  OAI22_X1 U21637 ( .A1(n25355), .A2(n12121), .B1(n21671), .B2(n1742), .ZN(
        n6859) );
  OAI22_X1 U21638 ( .A1(n22600), .A2(n12135), .B1(n395), .B2(n1740), .ZN(n6857) );
  OAI22_X1 U21639 ( .A1(n20831), .A2(n12149), .B1(n22032), .B2(n1738), .ZN(
        n68550) );
  OAI22_X1 U21640 ( .A1(n20855), .A2(n12163), .B1(n22068), .B2(n1736), .ZN(
        n68530) );
  OAI22_X1 U21641 ( .A1(n19097), .A2(n12177), .B1(n22104), .B2(n1734), .ZN(
        n68510) );
  OAI22_X1 U21642 ( .A1(n22561), .A2(n12191), .B1(n22330), .B2(n1732), .ZN(
        n68490) );
  OAI22_X1 U21643 ( .A1(n25046), .A2(n12205), .B1(n22354), .B2(n1730), .ZN(
        n68470) );
  OAI22_X1 U21644 ( .A1(n25063), .A2(n12219), .B1(n22378), .B2(n1728), .ZN(
        n68450) );
  OAI22_X1 U21645 ( .A1(n23966), .A2(n12233), .B1(n22402), .B2(n1726), .ZN(
        n68430) );
  OAI22_X1 U21646 ( .A1(n22549), .A2(n12247), .B1(n26429), .B2(n1724), .ZN(
        n68410) );
  OAI22_X1 U21647 ( .A1(n20833), .A2(n12261), .B1(n27114), .B2(n1722), .ZN(
        n6839) );
  OAI22_X1 U21648 ( .A1(n20858), .A2(n12275), .B1(n26447), .B2(n1720), .ZN(
        n6837) );
  OAI22_X1 U21649 ( .A1(n20772), .A2(n12289), .B1(n26453), .B2(n1718), .ZN(
        n6835) );
  OAI22_X1 U21650 ( .A1(n22572), .A2(n1780), .B1(n22324), .B2(n1716), .ZN(
        n6833) );
  OAI22_X1 U21651 ( .A1(n25034), .A2(n1778), .B1(n22348), .B2(n1714), .ZN(
        n6831) );
  OAI22_X1 U21652 ( .A1(n25050), .A2(n1776), .B1(n22372), .B2(n1712), .ZN(
        n6829) );
  OAI22_X1 U21653 ( .A1(n25365), .A2(n1774), .B1(n22396), .B2(n1710), .ZN(
        n6827) );
  OAI22_X1 U21654 ( .A1(n22577), .A2(n1772), .B1(n21996), .B2(n1708), .ZN(
        n6825) );
  OAI22_X1 U21655 ( .A1(n23931), .A2(n1770), .B1(n26411), .B2(n1706), .ZN(
        n6823) );
  OAI22_X1 U21656 ( .A1(n23883), .A2(n1768), .B1(n26417), .B2(n1704), .ZN(
        n6821) );
  OAI22_X1 U21657 ( .A1(n20756), .A2(n1766), .B1(n26423), .B2(n1702), .ZN(
        n6819) );
  OAI22_X1 U21658 ( .A1(n22588), .A2(n1764), .B1(n26209), .B2(n1700), .ZN(
        n6817) );
  OAI22_X1 U21659 ( .A1(n25041), .A2(n1762), .B1(n26217), .B2(n1698), .ZN(
        n6815) );
  OAI22_X1 U21660 ( .A1(n25057), .A2(n1760), .B1(n26225), .B2(n1696), .ZN(
        n6813) );
  OAI22_X1 U21661 ( .A1(n25354), .A2(n1758), .B1(n26233), .B2(n1694), .ZN(
        n6811) );
  OAI22_X1 U21662 ( .A1(n22592), .A2(n1756), .B1(n22170), .B2(n1692), .ZN(
        n6809) );
  OAI22_X1 U21663 ( .A1(n23919), .A2(n1754), .B1(n70), .B2(n1690), .ZN(n6807)
         );
  OAI22_X1 U21664 ( .A1(n23871), .A2(n1752), .B1(n26446), .B2(n1688), .ZN(
        n6805) );
  OAI22_X1 U21665 ( .A1(n20764), .A2(n1750), .B1(n26452), .B2(n1686), .ZN(
        n6803) );
  OAI22_X1 U21666 ( .A1(n22604), .A2(n1748), .B1(n26177), .B2(n1684), .ZN(
        n68010) );
  OAI22_X1 U21667 ( .A1(n23907), .A2(n1746), .B1(n26181), .B2(n1682), .ZN(
        n67990) );
  OAI22_X1 U21668 ( .A1(n23859), .A2(n1744), .B1(n26185), .B2(n1680), .ZN(
        n67970) );
  OAI22_X1 U21669 ( .A1(n20777), .A2(n1742), .B1(n26189), .B2(n1678), .ZN(
        n67950) );
  OAI22_X1 U21670 ( .A1(n22552), .A2(n1740), .B1(n26405), .B2(n1676), .ZN(
        n67930) );
  OAI22_X1 U21671 ( .A1(n23895), .A2(n1738), .B1(n26412), .B2(n1674), .ZN(
        n67910) );
  OAI22_X1 U21672 ( .A1(n23847), .A2(n1736), .B1(n26418), .B2(n1672), .ZN(
        n67890) );
  OAI22_X1 U21673 ( .A1(n24977), .A2(n1734), .B1(n26424), .B2(n1670), .ZN(
        n67870) );
  OAI22_X1 U21674 ( .A1(n23769), .A2(n1732), .B1(n26406), .B2(n1668), .ZN(
        n67850) );
  OAI22_X1 U21675 ( .A1(n23925), .A2(n1730), .B1(n26165), .B2(n1666), .ZN(
        n67830) );
  OAI22_X1 U21676 ( .A1(n23877), .A2(n1728), .B1(n26169), .B2(n1664), .ZN(
        n6781) );
  OAI22_X1 U21677 ( .A1(n24981), .A2(n1726), .B1(n26173), .B2(n1662), .ZN(
        n6779) );
  OAI22_X1 U21678 ( .A1(n22608), .A2(n1724), .B1(n26211), .B2(n1660), .ZN(
        n6777) );
  OAI22_X1 U21679 ( .A1(n20828), .A2(n1722), .B1(n26219), .B2(n1658), .ZN(
        n6775) );
  OAI22_X1 U21680 ( .A1(n20852), .A2(n1720), .B1(n26227), .B2(n1656), .ZN(
        n6773) );
  OAI22_X1 U21681 ( .A1(n24126), .A2(n1718), .B1(n26235), .B2(n1654), .ZN(
        n6771) );
  OAI22_X1 U21682 ( .A1(n23793), .A2(n1716), .B1(n22145), .B2(n1652), .ZN(
        n6769) );
  OAI22_X1 U21683 ( .A1(n23913), .A2(n1714), .B1(n69), .B2(n1650), .ZN(n6767)
         );
  OAI22_X1 U21684 ( .A1(n23865), .A2(n1712), .B1(n26448), .B2(n1648), .ZN(
        n6765) );
  OAI22_X1 U21685 ( .A1(n19101), .A2(n1710), .B1(n26454), .B2(n1646), .ZN(
        n67630) );
  OAI22_X1 U21686 ( .A1(n22556), .A2(n1708), .B1(n26481), .B2(n1644), .ZN(
        n67610) );
  OAI22_X1 U21687 ( .A1(n20838), .A2(n1706), .B1(n26485), .B2(n1642), .ZN(
        n67590) );
  OAI22_X1 U21688 ( .A1(n20864), .A2(n1704), .B1(n26489), .B2(n1640), .ZN(
        n67570) );
  OAI22_X1 U21689 ( .A1(n22674), .A2(n1702), .B1(n26493), .B2(n1638), .ZN(
        n67550) );
  OAI22_X1 U21690 ( .A1(n23818), .A2(n1700), .B1(n26161), .B2(n1636), .ZN(
        n67530) );
  OAI22_X1 U21691 ( .A1(n23901), .A2(n1698), .B1(n26414), .B2(n1634), .ZN(
        n67510) );
  OAI22_X1 U21692 ( .A1(n23853), .A2(n1696), .B1(n264201), .B2(n1632), .ZN(
        n67490) );
  OAI22_X1 U21693 ( .A1(n25351), .A2(n1694), .B1(n26426), .B2(n1630), .ZN(
        n6747) );
  OAI22_X1 U21694 ( .A1(n23775), .A2(n1692), .B1(n264801), .B2(n1628), .ZN(
        n6745) );
  OAI22_X1 U21695 ( .A1(n23933), .A2(n1690), .B1(n26484), .B2(n1626), .ZN(
        n6743) );
  OAI22_X1 U21696 ( .A1(n23885), .A2(n1688), .B1(n26488), .B2(n1624), .ZN(
        n6741) );
  OAI22_X1 U21697 ( .A1(n24114), .A2(n1686), .B1(n26492), .B2(n1622), .ZN(
        n6739) );
  OAI22_X1 U21698 ( .A1(n23763), .A2(n1684), .B1(n22126), .B2(n1620), .ZN(
        n6737) );
  OAI22_X1 U21699 ( .A1(n23889), .A2(n1682), .B1(n22170), .B2(n1618), .ZN(
        n6735) );
  OAI22_X1 U21700 ( .A1(n23841), .A2(n1680), .B1(n22222), .B2(n1616), .ZN(
        n6733) );
  OAI22_X1 U21701 ( .A1(n25228), .A2(n1678), .B1(n22257), .B2(n1614), .ZN(
        n6731) );
  OAI22_X1 U21702 ( .A1(n23781), .A2(n1676), .B1(n22132), .B2(n1612), .ZN(
        n6729) );
  OAI22_X1 U21703 ( .A1(n20816), .A2(n1674), .B1(n22176), .B2(n1610), .ZN(
        n6727) );
  OAI22_X1 U21704 ( .A1(n20840), .A2(n1672), .B1(n22215), .B2(n1608), .ZN(
        n6725) );
  OAI22_X1 U21705 ( .A1(n19059), .A2(n1670), .B1(n22251), .B2(n1606), .ZN(
        n6723) );
  OAI22_X1 U21706 ( .A1(n23799), .A2(n1668), .B1(n26408), .B2(n1604), .ZN(
        n6721) );
  OAI22_X1 U21707 ( .A1(n20827), .A2(n1666), .B1(n22017), .B2(n1602), .ZN(
        n67190) );
  OAI22_X1 U21708 ( .A1(n20851), .A2(n1664), .B1(n22053), .B2(n1600), .ZN(
        n67170) );
  OAI22_X1 U21709 ( .A1(n25240), .A2(n1662), .B1(n22089), .B2(n1598), .ZN(
        n67150) );
  OAI22_X1 U21710 ( .A1(n23823), .A2(n1660), .B1(n21981), .B2(n1596), .ZN(
        n67130) );
  OAI22_X1 U21711 ( .A1(n20829), .A2(n1658), .B1(n22023), .B2(n1594), .ZN(
        n67110) );
  OAI22_X1 U21712 ( .A1(n20853), .A2(n1656), .B1(n22059), .B2(n1592), .ZN(
        n67090) );
  OAI22_X1 U21713 ( .A1(n25231), .A2(n1654), .B1(n22095), .B2(n1590), .ZN(
        n67070) );
  OAI22_X1 U21714 ( .A1(n23806), .A2(n1652), .B1(n26208), .B2(n1588), .ZN(
        n67050) );
  OAI22_X1 U21715 ( .A1(n23922), .A2(n1650), .B1(n26216), .B2(n1586), .ZN(
        n67030) );
  OAI22_X1 U21716 ( .A1(n23874), .A2(n1648), .B1(n26224), .B2(n1584), .ZN(
        n67010) );
  OAI22_X1 U21717 ( .A1(n24138), .A2(n1646), .B1(n26232), .B2(n1582), .ZN(
        n6699) );
  OAI22_X1 U21718 ( .A1(n23746), .A2(n1644), .B1(n26176), .B2(n1580), .ZN(
        n6697) );
  OAI22_X1 U21719 ( .A1(n20839), .A2(n1642), .B1(n26180), .B2(n1578), .ZN(
        n6695) );
  OAI22_X1 U21720 ( .A1(n20865), .A2(n1640), .B1(n26184), .B2(n1576), .ZN(
        n6693) );
  OAI22_X1 U21721 ( .A1(n24115), .A2(n1638), .B1(n26188), .B2(n1574), .ZN(
        n6691) );
  OAI22_X1 U21722 ( .A1(n23830), .A2(n1636), .B1(n26210), .B2(n1572), .ZN(
        n6689) );
  OAI22_X1 U21723 ( .A1(n23909), .A2(n1634), .B1(n26218), .B2(n1570), .ZN(
        n6687) );
  OAI22_X1 U21724 ( .A1(n23861), .A2(n1632), .B1(n26226), .B2(n1568), .ZN(
        n6685) );
  OAI22_X1 U21725 ( .A1(n24120), .A2(n1630), .B1(n26234), .B2(n1566), .ZN(
        n6683) );
  OAI22_X1 U21726 ( .A1(n23787), .A2(n1628), .B1(n21987), .B2(n1564), .ZN(
        n66810) );
  OAI22_X1 U21727 ( .A1(n20817), .A2(n1626), .B1(n26164), .B2(n1562), .ZN(
        n66790) );
  OAI22_X1 U21728 ( .A1(n20841), .A2(n1624), .B1(n26168), .B2(n1560), .ZN(
        n66770) );
  OAI22_X1 U21729 ( .A1(n24139), .A2(n1622), .B1(n26172), .B2(n1558), .ZN(
        n66750) );
  OAI22_X1 U21730 ( .A1(n23752), .A2(n1620), .B1(n22333), .B2(n1556), .ZN(
        n66730) );
  OAI22_X1 U21731 ( .A1(n23897), .A2(n1618), .B1(n22357), .B2(n1554), .ZN(
        n66710) );
  OAI22_X1 U21732 ( .A1(n23849), .A2(n1616), .B1(n22381), .B2(n1552), .ZN(
        n66690) );
  OAI22_X1 U21733 ( .A1(n23962), .A2(n1614), .B1(n22405), .B2(n1550), .ZN(
        n66670) );
  OAI22_X1 U21734 ( .A1(n23811), .A2(n1612), .B1(n22146), .B2(n1548), .ZN(
        n6665) );
  OAI22_X1 U21735 ( .A1(n20826), .A2(n1610), .B1(n22192), .B2(n1546), .ZN(
        n6663) );
  OAI22_X1 U21736 ( .A1(n20850), .A2(n1608), .B1(n22227), .B2(n1544), .ZN(
        n6661) );
  OAI22_X1 U21737 ( .A1(n24128), .A2(n1606), .B1(n22262), .B2(n1542), .ZN(
        n6659) );
  OAI22_X1 U21738 ( .A1(n23836), .A2(n1604), .B1(n22124), .B2(n1540), .ZN(
        n6657) );
  OAI22_X1 U21739 ( .A1(n25042), .A2(n1602), .B1(n22168), .B2(n1538), .ZN(
        n6655) );
  OAI22_X1 U21740 ( .A1(n25058), .A2(n1600), .B1(n22220), .B2(n1536), .ZN(
        n6653) );
  OAI22_X1 U21741 ( .A1(n24109), .A2(n1598), .B1(n22282), .B2(n1534), .ZN(
        n6651) );
  OAI22_X1 U21742 ( .A1(n23757), .A2(n1596), .B1(n26160), .B2(n1532), .ZN(
        n6649) );
  OAI22_X1 U21743 ( .A1(n25049), .A2(n1594), .B1(n22035), .B2(n1530), .ZN(
        n6647) );
  OAI22_X1 U21744 ( .A1(n25066), .A2(n1592), .B1(n22071), .B2(n1528), .ZN(
        n6645) );
  OAI22_X1 U21745 ( .A1(n24133), .A2(n1590), .B1(n22107), .B2(n1526), .ZN(
        n6643) );
  OAI22_X1 U21746 ( .A1(n23771), .A2(n1588), .B1(n21999), .B2(n1524), .ZN(
        n6641) );
  OAI22_X1 U21747 ( .A1(n22673), .A2(n1586), .B1(n22016), .B2(n1522), .ZN(
        n6639) );
  OAI22_X1 U21748 ( .A1(n22641), .A2(n1584), .B1(n22052), .B2(n1520), .ZN(
        n6637) );
  OAI22_X1 U21749 ( .A1(n24121), .A2(n1582), .B1(n22088), .B2(n1518), .ZN(
        n6635) );
  OAI22_X1 U21750 ( .A1(n23777), .A2(n1580), .B1(n22327), .B2(n1516), .ZN(
        n6633) );
  OAI22_X1 U21751 ( .A1(n23927), .A2(n1578), .B1(n22351), .B2(n1514), .ZN(
        n6631) );
  OAI22_X1 U21752 ( .A1(n23879), .A2(n1576), .B1(n22375), .B2(n1512), .ZN(
        n6629) );
  OAI22_X1 U21753 ( .A1(n24108), .A2(n1574), .B1(n22399), .B2(n1510), .ZN(
        n6627) );
  OAI22_X1 U21754 ( .A1(n23795), .A2(n1572), .B1(n22130), .B2(n1508), .ZN(
        n6625) );
  OAI22_X1 U21755 ( .A1(n22665), .A2(n1570), .B1(n22174), .B2(n1506), .ZN(
        n6623) );
  OAI22_X1 U21756 ( .A1(n22633), .A2(n1568), .B1(n22214), .B2(n1504), .ZN(
        n6621) );
  OAI22_X1 U21757 ( .A1(n25225), .A2(n1566), .B1(n22250), .B2(n1502), .ZN(
        n66190) );
  OAI22_X1 U21758 ( .A1(n23801), .A2(n1564), .B1(n21714), .B2(n1500), .ZN(
        n66170) );
  OAI22_X1 U21759 ( .A1(n23915), .A2(n1562), .B1(n21730), .B2(n1498), .ZN(
        n66150) );
  OAI22_X1 U21760 ( .A1(n23867), .A2(n1560), .B1(n21746), .B2(n1496), .ZN(
        n66130) );
  OAI22_X1 U21761 ( .A1(n24132), .A2(n1558), .B1(n21762), .B2(n1494), .ZN(
        n66110) );
  OAI22_X1 U21762 ( .A1(n23820), .A2(n1556), .B1(n21980), .B2(n1492), .ZN(
        n66090) );
  OAI22_X1 U21763 ( .A1(n22657), .A2(n1554), .B1(n22021), .B2(n1490), .ZN(
        n66070) );
  OAI22_X1 U21764 ( .A1(n22625), .A2(n1552), .B1(n22057), .B2(n1488), .ZN(
        n66050) );
  OAI22_X1 U21765 ( .A1(n25238), .A2(n1550), .B1(n22093), .B2(n1486), .ZN(
        n66030) );
  OAI22_X1 U21766 ( .A1(n23826), .A2(n1548), .B1(n21717), .B2(n1484), .ZN(
        n66010) );
  OAI22_X1 U21767 ( .A1(n23904), .A2(n1546), .B1(n21733), .B2(n1482), .ZN(
        n6599) );
  OAI22_X1 U21768 ( .A1(n23856), .A2(n1544), .B1(n21749), .B2(n1480), .ZN(
        n6597) );
  OAI22_X1 U21769 ( .A1(n25227), .A2(n1542), .B1(n21765), .B2(n1478), .ZN(
        n6595) );
  OAI22_X1 U21770 ( .A1(n23765), .A2(n1540), .B1(n21682), .B2(n1476), .ZN(
        n6593) );
  OAI22_X1 U21771 ( .A1(n22649), .A2(n1538), .B1(n21690), .B2(n1474), .ZN(
        n6591) );
  OAI22_X1 U21772 ( .A1(n22617), .A2(n1536), .B1(n21698), .B2(n1472), .ZN(
        n6589) );
  OAI22_X1 U21773 ( .A1(n19095), .A2(n1534), .B1(n21706), .B2(n1470), .ZN(
        n6587) );
  OAI22_X1 U21774 ( .A1(n23784), .A2(n1532), .B1(n22145), .B2(n1468), .ZN(
        n6585) );
  OAI22_X1 U21775 ( .A1(n22668), .A2(n1530), .B1(n22191), .B2(n1466), .ZN(
        n6583) );
  OAI22_X1 U21776 ( .A1(n22636), .A2(n1528), .B1(n22225), .B2(n1464), .ZN(
        n65810) );
  OAI22_X1 U21777 ( .A1(n25226), .A2(n1526), .B1(n22260), .B2(n1462), .ZN(
        n65790) );
  OAI22_X1 U21778 ( .A1(n23808), .A2(n1524), .B1(n21985), .B2(n1460), .ZN(
        n65770) );
  OAI22_X1 U21779 ( .A1(n22661), .A2(n1522), .B1(n21658), .B2(n1458), .ZN(
        n65750) );
  OAI22_X1 U21780 ( .A1(n22629), .A2(n1520), .B1(n21666), .B2(n1456), .ZN(
        n65730) );
  OAI22_X1 U21781 ( .A1(n19063), .A2(n1518), .B1(n21674), .B2(n1454), .ZN(
        n65710) );
  OAI22_X1 U21782 ( .A1(n23832), .A2(n1516), .B1(n21650), .B2(n1452), .ZN(
        n65690) );
  OAI22_X1 U21783 ( .A1(n22653), .A2(n1514), .B1(n22034), .B2(n1450), .ZN(
        n65670) );
  OAI22_X1 U21784 ( .A1(n22621), .A2(n1512), .B1(n22070), .B2(n1448), .ZN(
        n6565) );
  OAI22_X1 U21785 ( .A1(n19058), .A2(n1510), .B1(n22106), .B2(n1446), .ZN(
        n65630) );
  OAI22_X1 U21786 ( .A1(n23747), .A2(n1508), .B1(n22331), .B2(n1444), .ZN(
        n6561) );
  OAI22_X1 U21787 ( .A1(n23891), .A2(n1506), .B1(n22355), .B2(n1442), .ZN(
        n6559) );
  OAI22_X1 U21788 ( .A1(n23843), .A2(n1504), .B1(n22379), .B2(n1440), .ZN(
        n6557) );
  OAI22_X1 U21789 ( .A1(n23963), .A2(n1502), .B1(n22403), .B2(n1438), .ZN(
        n6555) );
  OAI22_X1 U21790 ( .A1(n23754), .A2(n1500), .B1(n22121), .B2(n1436), .ZN(
        n6553) );
  OAI22_X1 U21791 ( .A1(n22644), .A2(n1498), .B1(n22164), .B2(n1434), .ZN(
        n6551) );
  OAI22_X1 U21792 ( .A1(n22612), .A2(n1496), .B1(n22217), .B2(n1432), .ZN(
        n6549) );
  OAI22_X1 U21793 ( .A1(n24113), .A2(n1494), .B1(n22253), .B2(n1430), .ZN(
        n6547) );
  OAI22_X1 U21794 ( .A1(n23790), .A2(n1492), .B1(n22325), .B2(n1428), .ZN(
        n6545) );
  OAI22_X1 U21795 ( .A1(n20812), .A2(n1490), .B1(n22349), .B2(n1426), .ZN(
        n6543) );
  OAI22_X1 U21796 ( .A1(n20836), .A2(n1488), .B1(n22373), .B2(n1424), .ZN(
        n6541) );
  OAI22_X1 U21797 ( .A1(n19056), .A2(n1486), .B1(n22397), .B2(n1422), .ZN(
        n6539) );
  OAI22_X1 U21798 ( .A1(n22563), .A2(n1484), .B1(n21998), .B2(n1420), .ZN(
        n65370) );
  OAI22_X1 U21799 ( .A1(n25034), .A2(n1482), .B1(n22013), .B2(n1418), .ZN(
        n65350) );
  OAI22_X1 U21800 ( .A1(n25050), .A2(n1480), .B1(n22049), .B2(n1416), .ZN(
        n65330) );
  OAI22_X1 U21801 ( .A1(n24137), .A2(n1478), .B1(n22085), .B2(n1414), .ZN(
        n65310) );
  OAI22_X1 U21802 ( .A1(n23814), .A2(n1476), .B1(n21711), .B2(n1412), .ZN(
        n65290) );
  OAI22_X1 U21803 ( .A1(n20826), .A2(n1474), .B1(n21727), .B2(n1410), .ZN(
        n65270) );
  OAI22_X1 U21804 ( .A1(n20850), .A2(n1472), .B1(n21743), .B2(n1408), .ZN(
        n65250) );
  OAI22_X1 U21805 ( .A1(n19096), .A2(n1470), .B1(n21759), .B2(n1406), .ZN(
        n65230) );
  OAI22_X1 U21806 ( .A1(n22579), .A2(n1468), .B1(n22128), .B2(n1404), .ZN(
        n65210) );
  OAI22_X1 U21807 ( .A1(n25041), .A2(n1466), .B1(n22172), .B2(n1402), .ZN(
        n65190) );
  OAI22_X1 U21808 ( .A1(n25057), .A2(n1464), .B1(n22211), .B2(n1400), .ZN(
        n6517) );
  OAI22_X1 U21809 ( .A1(n24125), .A2(n1462), .B1(n22247), .B2(n1398), .ZN(
        n6515) );
  OAI22_X1 U21810 ( .A1(n23837), .A2(n1460), .B1(n21679), .B2(n27884), .ZN(
        n6513) );
  INV_X1 U21811 ( .A(sram_rdata_w1[0]), .ZN(n27884) );
  OAI22_X1 U21812 ( .A1(n20665), .A2(n1458), .B1(n21687), .B2(n27882), .ZN(
        n6511) );
  INV_X1 U21813 ( .A(sram_rdata_w1[2]), .ZN(n27882) );
  OAI22_X1 U21814 ( .A1(n20632), .A2(n1456), .B1(n21695), .B2(n27880), .ZN(
        n6509) );
  INV_X1 U21815 ( .A(sram_rdata_w1[4]), .ZN(n27880) );
  OAI22_X1 U21816 ( .A1(n24107), .A2(n1454), .B1(n21703), .B2(n27878), .ZN(
        n6507) );
  INV_X1 U21817 ( .A(sram_rdata_w1[6]), .ZN(n27878) );
  OAI22_X1 U21818 ( .A1(n23760), .A2(n1452), .B1(n21978), .B2(n27876), .ZN(
        n6505) );
  INV_X1 U21819 ( .A(sram_rdata_w1[8]), .ZN(n27876) );
  OAI22_X1 U21820 ( .A1(n20838), .A2(n1450), .B1(n22019), .B2(n27874), .ZN(
        n6503) );
  INV_X1 U21821 ( .A(sram_rdata_w1[10]), .ZN(n27874) );
  OAI22_X1 U21822 ( .A1(n20864), .A2(n1448), .B1(n22055), .B2(n27872), .ZN(
        n6501) );
  INV_X1 U21823 ( .A(sram_rdata_w1[12]), .ZN(n27872) );
  OAI22_X1 U21824 ( .A1(n24131), .A2(n1446), .B1(n22091), .B2(n27870), .ZN(
        n64990) );
  INV_X1 U21825 ( .A(sram_rdata_w1[14]), .ZN(n27870) );
  OAI22_X1 U21826 ( .A1(n22566), .A2(n1444), .B1(n21983), .B2(n27868), .ZN(
        n64970) );
  INV_X1 U21827 ( .A(sram_rdata_w1[16]), .ZN(n27868) );
  OAI22_X1 U21828 ( .A1(n20685), .A2(n1442), .B1(n21655), .B2(n27866), .ZN(
        n64950) );
  INV_X1 U21829 ( .A(sram_rdata_w1[18]), .ZN(n27866) );
  OAI22_X1 U21830 ( .A1(n20653), .A2(n1440), .B1(n21663), .B2(n27864), .ZN(
        n64930) );
  INV_X1 U21831 ( .A(sram_rdata_w1[20]), .ZN(n27864) );
  OAI22_X1 U21832 ( .A1(n24119), .A2(n1438), .B1(n21671), .B2(n27862), .ZN(
        n64910) );
  INV_X1 U21833 ( .A(sram_rdata_w1[22]), .ZN(n27862) );
  OAI22_X1 U21834 ( .A1(n22594), .A2(n1436), .B1(n21715), .B2(n278601), .ZN(
        n64890) );
  INV_X1 U21835 ( .A(sram_rdata_w1[24]), .ZN(n278601) );
  OAI22_X1 U21836 ( .A1(n20828), .A2(n1434), .B1(n21731), .B2(n27858), .ZN(
        n64870) );
  INV_X1 U21837 ( .A(sram_rdata_w1[26]), .ZN(n27858) );
  OAI22_X1 U21838 ( .A1(n20852), .A2(n1432), .B1(n21747), .B2(n27856), .ZN(
        n64850) );
  INV_X1 U21839 ( .A(sram_rdata_w1[28]), .ZN(n27856) );
  OAI22_X1 U21840 ( .A1(n25231), .A2(n1430), .B1(n21763), .B2(n27854), .ZN(
        n6483) );
  INV_X1 U21841 ( .A(sram_rdata_w1[30]), .ZN(n27854) );
  OAI22_X1 U21842 ( .A1(n22582), .A2(n1428), .B1(n22142), .B2(n27852), .ZN(
        n6481) );
  INV_X1 U21843 ( .A(sram_rdata_w0[0]), .ZN(n27852) );
  OAI22_X1 U21844 ( .A1(n20677), .A2(n1426), .B1(n22188), .B2(n278501), .ZN(
        n6479) );
  INV_X1 U21845 ( .A(sram_rdata_w0[2]), .ZN(n278501) );
  OAI22_X1 U21846 ( .A1(n20645), .A2(n1424), .B1(n22223), .B2(n27848), .ZN(
        n6477) );
  INV_X1 U21847 ( .A(sram_rdata_w0[4]), .ZN(n27848) );
  OAI22_X1 U21848 ( .A1(n19057), .A2(n1422), .B1(n22258), .B2(n27846), .ZN(
        n6475) );
  INV_X1 U21849 ( .A(sram_rdata_w0[6]), .ZN(n27846) );
  OAI22_X1 U21850 ( .A1(n22558), .A2(n1420), .B1(n22329), .B2(n27844), .ZN(
        n6473) );
  INV_X1 U21851 ( .A(sram_rdata_w0[8]), .ZN(n27844) );
  OAI22_X1 U21852 ( .A1(n24840), .A2(n1418), .B1(n22353), .B2(n27842), .ZN(
        n6471) );
  INV_X1 U21853 ( .A(sram_rdata_w0[10]), .ZN(n27842) );
  OAI22_X1 U21854 ( .A1(n24823), .A2(n1416), .B1(n22377), .B2(n278401), .ZN(
        n6469) );
  INV_X1 U21855 ( .A(sram_rdata_w0[12]), .ZN(n278401) );
  OAI22_X1 U21856 ( .A1(n23965), .A2(n1414), .B1(n22401), .B2(n27838), .ZN(
        n6467) );
  INV_X1 U21857 ( .A(sram_rdata_w0[14]), .ZN(n27838) );
  OAI22_X1 U21858 ( .A1(n22598), .A2(n1412), .B1(n395), .B2(n27836), .ZN(n6465) );
  INV_X1 U21859 ( .A(sram_rdata_w0[16]), .ZN(n27836) );
  OAI22_X1 U21860 ( .A1(n20669), .A2(n1410), .B1(n22031), .B2(n27834), .ZN(
        n6463) );
  INV_X1 U21861 ( .A(sram_rdata_w0[18]), .ZN(n27834) );
  OAI22_X1 U21862 ( .A1(n20636), .A2(n1408), .B1(n22067), .B2(n27832), .ZN(
        n6461) );
  INV_X1 U21863 ( .A(sram_rdata_w0[20]), .ZN(n27832) );
  OAI22_X1 U21864 ( .A1(n19062), .A2(n1406), .B1(n22103), .B2(n278301), .ZN(
        n6459) );
  INV_X1 U21865 ( .A(sram_rdata_w0[22]), .ZN(n278301) );
  OAI22_X1 U21866 ( .A1(n22570), .A2(n1404), .B1(n22323), .B2(n27828), .ZN(
        n6457) );
  INV_X1 U21867 ( .A(sram_rdata_w0[24]), .ZN(n27828) );
  OAI22_X1 U21868 ( .A1(n24855), .A2(n1402), .B1(n22347), .B2(n27826), .ZN(
        n6455) );
  INV_X1 U21869 ( .A(sram_rdata_w0[26]), .ZN(n27826) );
  OAI22_X1 U21870 ( .A1(n24839), .A2(n1400), .B1(n22371), .B2(n27824), .ZN(
        n6453) );
  INV_X1 U21871 ( .A(sram_rdata_w0[28]), .ZN(n27824) );
  OAI22_X1 U21872 ( .A1(n25229), .A2(n1398), .B1(n22395), .B2(n27822), .ZN(
        n6451) );
  INV_X1 U21873 ( .A(sram_rdata_w0[30]), .ZN(n27822) );
  OAI22_X1 U21874 ( .A1(n22547), .A2(n14254), .B1(n22135), .B2(n1387), .ZN(
        n74080) );
  OAI22_X1 U21875 ( .A1(n20661), .A2(n14268), .B1(n22180), .B2(n1385), .ZN(
        n74060) );
  OAI22_X1 U21876 ( .A1(n20628), .A2(n14282), .B1(n22230), .B2(n1383), .ZN(
        n74040) );
  OAI22_X1 U21877 ( .A1(n19058), .A2(n14296), .B1(n23582), .B2(n1381), .ZN(
        n74020) );
  OAI22_X1 U21878 ( .A1(n22587), .A2(n1387), .B1(n21723), .B2(n1379), .ZN(
        n74000) );
  OAI22_X1 U21879 ( .A1(n24851), .A2(n1385), .B1(n21739), .B2(n1377), .ZN(
        n73980) );
  OAI22_X1 U21880 ( .A1(n24835), .A2(n1383), .B1(n21755), .B2(n1375), .ZN(
        n73960) );
  OAI22_X1 U21881 ( .A1(n25241), .A2(n1381), .B1(n21771), .B2(n1373), .ZN(
        n73940) );
  OAI22_X1 U21882 ( .A1(n22575), .A2(n1379), .B1(n21659), .B2(n1371), .ZN(
        n7392) );
  OAI22_X1 U21883 ( .A1(n22670), .A2(n1377), .B1(n21667), .B2(n1369), .ZN(
        n7390) );
  OAI22_X1 U21884 ( .A1(n22638), .A2(n1375), .B1(n21675), .B2(n1367), .ZN(
        n7388) );
  OAI22_X1 U21885 ( .A1(n25223), .A2(n1373), .B1(n21683), .B2(n1365), .ZN(
        n7386) );
  OAI22_X1 U21886 ( .A1(n22603), .A2(n1371), .B1(n22341), .B2(n1363), .ZN(
        n7384) );
  OAI22_X1 U21887 ( .A1(n20670), .A2(n1369), .B1(n22365), .B2(n1361), .ZN(
        n7382) );
  OAI22_X1 U21888 ( .A1(n20637), .A2(n1367), .B1(n22389), .B2(n1359), .ZN(
        n7380) );
  OAI22_X1 U21889 ( .A1(n24976), .A2(n1365), .B1(n22413), .B2(n1357), .ZN(
        n7378) );
  OAI22_X1 U21890 ( .A1(n22591), .A2(n1363), .B1(n21691), .B2(n1355), .ZN(
        n7376) );
  OAI22_X1 U21891 ( .A1(n22662), .A2(n1361), .B1(n21699), .B2(n1353), .ZN(
        n73740) );
  OAI22_X1 U21892 ( .A1(n22630), .A2(n1359), .B1(n21707), .B2(n1351), .ZN(
        n73720) );
  OAI22_X1 U21893 ( .A1(n25236), .A2(n1357), .B1(n23585), .B2(n1349), .ZN(
        n73700) );
  OAI22_X1 U21894 ( .A1(n22606), .A2(n1355), .B1(n22150), .B2(n1347), .ZN(
        n73680) );
  OAI22_X1 U21895 ( .A1(n22655), .A2(n1353), .B1(n22195), .B2(n1345), .ZN(
        n73660) );
  OAI22_X1 U21896 ( .A1(n22623), .A2(n1351), .B1(n22241), .B2(n1343), .ZN(
        n73640) );
  OAI22_X1 U21897 ( .A1(n25233), .A2(n1349), .B1(n22275), .B2(n1341), .ZN(
        n73620) );
  OAI22_X1 U21898 ( .A1(n22550), .A2(n1347), .B1(n22001), .B2(n27947), .ZN(
        n73600) );
  INV_X1 U21899 ( .A(sram_rdata_d1[1]), .ZN(n27947) );
  OAI22_X1 U21900 ( .A1(n22646), .A2(n1345), .B1(n22037), .B2(n27945), .ZN(
        n7358) );
  INV_X1 U21901 ( .A(sram_rdata_d1[3]), .ZN(n27945) );
  OAI22_X1 U21902 ( .A1(n22614), .A2(n1343), .B1(n22073), .B2(n27943), .ZN(
        n7356) );
  INV_X1 U21903 ( .A(sram_rdata_d1[5]), .ZN(n27943) );
  OAI22_X1 U21904 ( .A1(n24980), .A2(n1341), .B1(n22109), .B2(n27941), .ZN(
        n7354) );
  INV_X1 U21905 ( .A(sram_rdata_d1[7]), .ZN(n27941) );
  OAI22_X1 U21906 ( .A1(n22565), .A2(n14574), .B1(n264101), .B2(n1331), .ZN(
        n7344) );
  OAI22_X1 U21907 ( .A1(n22666), .A2(n14588), .B1(n26416), .B2(n1329), .ZN(
        n7342) );
  OAI22_X1 U21908 ( .A1(n22634), .A2(n14602), .B1(n27122), .B2(n1327), .ZN(
        n7340) );
  OAI22_X1 U21909 ( .A1(n20750), .A2(n14616), .B1(n26428), .B2(n1325), .ZN(
        n7338) );
  OAI22_X1 U21910 ( .A1(n22555), .A2(n1331), .B1(n22336), .B2(n1323), .ZN(
        n7336) );
  OAI22_X1 U21911 ( .A1(n20662), .A2(n1329), .B1(n22360), .B2(n1321), .ZN(
        n7334) );
  OAI22_X1 U21912 ( .A1(n20629), .A2(n1327), .B1(n22384), .B2(n1319), .ZN(
        n7332) );
  OAI22_X1 U21913 ( .A1(n20767), .A2(n1325), .B1(n22408), .B2(n1317), .ZN(
        n7330) );
  OAI22_X1 U21914 ( .A1(n22581), .A2(n1323), .B1(n27113), .B2(n1315), .ZN(
        n7328) );
  OAI22_X1 U21915 ( .A1(n22658), .A2(n1321), .B1(n26445), .B2(n1313), .ZN(
        n7326) );
  OAI22_X1 U21916 ( .A1(n22626), .A2(n1319), .B1(n264501), .B2(n1311), .ZN(
        n73240) );
  OAI22_X1 U21917 ( .A1(n20758), .A2(n1317), .B1(n68), .B2(n1309), .ZN(n73220)
         );
  OAI22_X1 U21918 ( .A1(n22569), .A2(n1315), .B1(n26213), .B2(n1307), .ZN(
        n73200) );
  OAI22_X1 U21919 ( .A1(n23931), .A2(n1313), .B1(n26221), .B2(n1305), .ZN(
        n73180) );
  OAI22_X1 U21920 ( .A1(n23883), .A2(n1311), .B1(n26229), .B2(n1303), .ZN(
        n73160) );
  OAI22_X1 U21921 ( .A1(n24971), .A2(n1309), .B1(n26237), .B2(n1301), .ZN(
        n73140) );
  OAI22_X1 U21922 ( .A1(n22596), .A2(n1307), .B1(n26407), .B2(n1299), .ZN(
        n73120) );
  OAI22_X1 U21923 ( .A1(n22650), .A2(n1305), .B1(n26413), .B2(n1297), .ZN(
        n73100) );
  OAI22_X1 U21924 ( .A1(n22618), .A2(n1303), .B1(n26419), .B2(n1295), .ZN(
        n73080) );
  OAI22_X1 U21925 ( .A1(n20771), .A2(n1301), .B1(n26425), .B2(n1293), .ZN(
        n73060) );
  OAI22_X1 U21926 ( .A1(n22585), .A2(n1299), .B1(n26215), .B2(n1291), .ZN(
        n73040) );
  OAI22_X1 U21927 ( .A1(n23919), .A2(n1297), .B1(n26223), .B2(n1289), .ZN(
        n7302) );
  OAI22_X1 U21928 ( .A1(n23871), .A2(n1295), .B1(n26231), .B2(n1287), .ZN(
        n7300) );
  OAI22_X1 U21929 ( .A1(n24978), .A2(n1293), .B1(n26239), .B2(n1285), .ZN(
        n7298) );
  OAI22_X1 U21930 ( .A1(n22560), .A2(n1291), .B1(n26431), .B2(n27939), .ZN(
        n7296) );
  INV_X1 U21931 ( .A(sram_rdata_d1[9]), .ZN(n27939) );
  OAI22_X1 U21932 ( .A1(n22642), .A2(n1289), .B1(n26441), .B2(n27937), .ZN(
        n7294) );
  INV_X1 U21933 ( .A(sram_rdata_d1[11]), .ZN(n27937) );
  OAI22_X1 U21934 ( .A1(n22610), .A2(n1287), .B1(n26449), .B2(n27935), .ZN(
        n7292) );
  INV_X1 U21935 ( .A(sram_rdata_d1[13]), .ZN(n27935) );
  OAI22_X1 U21936 ( .A1(n20754), .A2(n1285), .B1(n23586), .B2(n27933), .ZN(
        n7290) );
  INV_X1 U21937 ( .A(sram_rdata_d1[15]), .ZN(n27933) );
  OAI22_X1 U21938 ( .A1(n22573), .A2(n14894), .B1(n26183), .B2(n1275), .ZN(
        n72800) );
  OAI22_X1 U21939 ( .A1(n20685), .A2(n14908), .B1(n26187), .B2(n1273), .ZN(
        n72780) );
  OAI22_X1 U21940 ( .A1(n20653), .A2(n14922), .B1(n26191), .B2(n1271), .ZN(
        n72760) );
  OAI22_X1 U21941 ( .A1(n20762), .A2(n14936), .B1(n22266), .B2(n1269), .ZN(
        n72740) );
  OAI22_X1 U21942 ( .A1(n22589), .A2(n1275), .B1(n26167), .B2(n1267), .ZN(
        n72720) );
  OAI22_X1 U21943 ( .A1(n24851), .A2(n1273), .B1(n26171), .B2(n1265), .ZN(
        n7270) );
  OAI22_X1 U21944 ( .A1(n24835), .A2(n1271), .B1(n26175), .B2(n1263), .ZN(
        n7268) );
  OAI22_X1 U21945 ( .A1(n25365), .A2(n1269), .B1(n26179), .B2(n1261), .ZN(
        n7266) );
  OAI22_X1 U21946 ( .A1(n22601), .A2(n1267), .B1(n26409), .B2(n1259), .ZN(
        n7264) );
  OAI22_X1 U21947 ( .A1(n20830), .A2(n1265), .B1(n26415), .B2(n1257), .ZN(
        n7262) );
  OAI22_X1 U21948 ( .A1(n20854), .A2(n1263), .B1(n26421), .B2(n1255), .ZN(
        n7260) );
  OAI22_X1 U21949 ( .A1(n19094), .A2(n1261), .B1(n26427), .B2(n1253), .ZN(
        n7258) );
  OAI22_X1 U21950 ( .A1(n22605), .A2(n1259), .B1(n26483), .B2(n1251), .ZN(
        n7256) );
  OAI22_X1 U21951 ( .A1(n23907), .A2(n1257), .B1(n26487), .B2(n1249), .ZN(
        n7254) );
  OAI22_X1 U21952 ( .A1(n23859), .A2(n1255), .B1(n26491), .B2(n1247), .ZN(
        n7252) );
  OAI22_X1 U21953 ( .A1(n24982), .A2(n1253), .B1(n26495), .B2(n1245), .ZN(
        n7250) );
  OAI22_X1 U21954 ( .A1(n22548), .A2(n1251), .B1(n26435), .B2(n1243), .ZN(
        n7248) );
  OAI22_X1 U21955 ( .A1(n24841), .A2(n1249), .B1(n26867), .B2(n1241), .ZN(
        n7246) );
  OAI22_X1 U21956 ( .A1(n24824), .A2(n1247), .B1(n26451), .B2(n1239), .ZN(
        n7244) );
  OAI22_X1 U21957 ( .A1(n19060), .A2(n1245), .B1(n26455), .B2(n1237), .ZN(
        n72420) );
  OAI22_X1 U21958 ( .A1(n22553), .A2(n1243), .B1(n26482), .B2(n1235), .ZN(
        n72400) );
  OAI22_X1 U21959 ( .A1(n23895), .A2(n1241), .B1(n26486), .B2(n1233), .ZN(
        n72380) );
  OAI22_X1 U21960 ( .A1(n23847), .A2(n1239), .B1(n264901), .B2(n1231), .ZN(
        n72360) );
  OAI22_X1 U21961 ( .A1(n20754), .A2(n1237), .B1(n26494), .B2(n1229), .ZN(
        n72340) );
  OAI22_X1 U21962 ( .A1(n22576), .A2(n1235), .B1(n22011), .B2(n27931), .ZN(
        n72320) );
  INV_X1 U21963 ( .A(sram_rdata_d1[17]), .ZN(n27931) );
  OAI22_X1 U21964 ( .A1(n20681), .A2(n1233), .B1(n22047), .B2(n27929), .ZN(
        n72300) );
  INV_X1 U21965 ( .A(sram_rdata_d1[19]), .ZN(n27929) );
  OAI22_X1 U21966 ( .A1(n20649), .A2(n1231), .B1(n22083), .B2(n27927), .ZN(
        n72280) );
  INV_X1 U21967 ( .A(sram_rdata_d1[21]), .ZN(n27927) );
  OAI22_X1 U21968 ( .A1(n17084), .A2(n1229), .B1(n22119), .B2(n27925), .ZN(
        n72260) );
  INV_X1 U21969 ( .A(sram_rdata_d1[23]), .ZN(n27925) );
  OAI22_X1 U21970 ( .A1(n23770), .A2(n15214), .B1(n26212), .B2(n1219), .ZN(
        n7216) );
  OAI22_X1 U21971 ( .A1(n23925), .A2(n15228), .B1(n26220), .B2(n1217), .ZN(
        n7214) );
  OAI22_X1 U21972 ( .A1(n23877), .A2(n15242), .B1(n26228), .B2(n1215), .ZN(
        n7212) );
  OAI22_X1 U21973 ( .A1(n19061), .A2(n15256), .B1(n26236), .B2(n1213), .ZN(
        n7210) );
  OAI22_X1 U21974 ( .A1(n22593), .A2(n1219), .B1(n22162), .B2(n1211), .ZN(
        n7208) );
  OAI22_X1 U21975 ( .A1(n24849), .A2(n1217), .B1(n22209), .B2(n1209), .ZN(
        n7206) );
  OAI22_X1 U21976 ( .A1(n24833), .A2(n1215), .B1(n22239), .B2(n1207), .ZN(
        n72040) );
  OAI22_X1 U21977 ( .A1(n19094), .A2(n1213), .B1(n22273), .B2(n1205), .ZN(
        n72020) );
  OAI22_X1 U21978 ( .A1(n22609), .A2(n1211), .B1(n22139), .B2(n1203), .ZN(
        n72000) );
  OAI22_X1 U21979 ( .A1(n24845), .A2(n1209), .B1(n22185), .B2(n1201), .ZN(
        n71980) );
  OAI22_X1 U21980 ( .A1(n24828), .A2(n1207), .B1(n22233), .B2(n1199), .ZN(
        n71960) );
  OAI22_X1 U21981 ( .A1(n25353), .A2(n1205), .B1(n22265), .B2(n1197), .ZN(
        n71940) );
  OAI22_X1 U21982 ( .A1(n22557), .A2(n1203), .B1(n21993), .B2(n1195), .ZN(
        n71920) );
  OAI22_X1 U21983 ( .A1(n24841), .A2(n1201), .B1(n22029), .B2(n1193), .ZN(
        n71900) );
  OAI22_X1 U21984 ( .A1(n24824), .A2(n1199), .B1(n22065), .B2(n1191), .ZN(
        n7188) );
  OAI22_X1 U21985 ( .A1(n20772), .A2(n1197), .B1(n22101), .B2(n1189), .ZN(
        n7186) );
  OAI22_X1 U21986 ( .A1(n23776), .A2(n1195), .B1(n26166), .B2(n1187), .ZN(
        n7184) );
  OAI22_X1 U21987 ( .A1(n23934), .A2(n1193), .B1(n26170), .B2(n1185), .ZN(
        n7182) );
  OAI22_X1 U21988 ( .A1(n23886), .A2(n1191), .B1(n26174), .B2(n1183), .ZN(
        n7180) );
  OAI22_X1 U21989 ( .A1(n20756), .A2(n1189), .B1(n26178), .B2(n1181), .ZN(
        n7178) );
  OAI22_X1 U21990 ( .A1(n23794), .A2(n1187), .B1(n26214), .B2(n1179), .ZN(
        n7176) );
  OAI22_X1 U21991 ( .A1(n23913), .A2(n1185), .B1(n26222), .B2(n1177), .ZN(
        n7174) );
  OAI22_X1 U21992 ( .A1(n23865), .A2(n1183), .B1(n26230), .B2(n1175), .ZN(
        n7172) );
  OAI22_X1 U21993 ( .A1(n19059), .A2(n1181), .B1(n26238), .B2(n1173), .ZN(
        n7170) );
  OAI22_X1 U21994 ( .A1(n23799), .A2(n1179), .B1(n26182), .B2(n27923), .ZN(
        n7168) );
  INV_X1 U21995 ( .A(sram_rdata_d1[25]), .ZN(n27923) );
  OAI22_X1 U21996 ( .A1(n23921), .A2(n1177), .B1(n26186), .B2(n27921), .ZN(
        n7166) );
  INV_X1 U21997 ( .A(sram_rdata_d1[27]), .ZN(n27921) );
  OAI22_X1 U21998 ( .A1(n23873), .A2(n1175), .B1(n26190), .B2(n27919), .ZN(
        n7164) );
  INV_X1 U21999 ( .A(sram_rdata_d1[29]), .ZN(n27919) );
  OAI22_X1 U22000 ( .A1(n24979), .A2(n1173), .B1(n23582), .B2(n27917), .ZN(
        n7162) );
  INV_X1 U22001 ( .A(sram_rdata_d1[31]), .ZN(n27917) );
  OAI22_X1 U22002 ( .A1(n23817), .A2(n15534), .B1(n22345), .B2(n1163), .ZN(
        n7152) );
  OAI22_X1 U22003 ( .A1(n23901), .A2(n15548), .B1(n22369), .B2(n1161), .ZN(
        n71500) );
  OAI22_X1 U22004 ( .A1(n23853), .A2(n15562), .B1(n22393), .B2(n1159), .ZN(
        n71480) );
  OAI22_X1 U22005 ( .A1(n25349), .A2(n15576), .B1(n22417), .B2(n1157), .ZN(
        n71460) );
  OAI22_X1 U22006 ( .A1(n23824), .A2(n1163), .B1(n22005), .B2(n1155), .ZN(
        n71440) );
  OAI22_X1 U22007 ( .A1(n23910), .A2(n1161), .B1(n22041), .B2(n1153), .ZN(
        n71420) );
  OAI22_X1 U22008 ( .A1(n23862), .A2(n1159), .B1(n22077), .B2(n1151), .ZN(
        n71400) );
  OAI22_X1 U22009 ( .A1(n20777), .A2(n1157), .B1(n22113), .B2(n1149), .ZN(
        n71380) );
  OAI22_X1 U22010 ( .A1(n23764), .A2(n1155), .B1(n22339), .B2(n1147), .ZN(
        n71360) );
  OAI22_X1 U22011 ( .A1(n23889), .A2(n1153), .B1(n22363), .B2(n1145), .ZN(
        n71340) );
  OAI22_X1 U22012 ( .A1(n23841), .A2(n1151), .B1(n22387), .B2(n1143), .ZN(
        n71320) );
  OAI22_X1 U22013 ( .A1(n25228), .A2(n1149), .B1(n22411), .B2(n1141), .ZN(
        n71300) );
  OAI22_X1 U22014 ( .A1(n23745), .A2(n1147), .B1(n22155), .B2(n1139), .ZN(
        n7128) );
  OAI22_X1 U22015 ( .A1(n23898), .A2(n1145), .B1(n22200), .B2(n1137), .ZN(
        n7126) );
  OAI22_X1 U22016 ( .A1(n23850), .A2(n1143), .B1(n22245), .B2(n1135), .ZN(
        n7124) );
  OAI22_X1 U22017 ( .A1(n20761), .A2(n1141), .B1(n22281), .B2(n1133), .ZN(
        n7122) );
  OAI22_X1 U22018 ( .A1(n23782), .A2(n1139), .B1(n22160), .B2(n1131), .ZN(
        n7120) );
  OAI22_X1 U22019 ( .A1(n23928), .A2(n1137), .B1(n22206), .B2(n1129), .ZN(
        n7118) );
  OAI22_X1 U22020 ( .A1(n23880), .A2(n1135), .B1(n22238), .B2(n1127), .ZN(
        n7116) );
  OAI22_X1 U22021 ( .A1(n20769), .A2(n1133), .B1(n22271), .B2(n1125), .ZN(
        n7114) );
  OAI22_X1 U22022 ( .A1(n23805), .A2(n1131), .B1(n22009), .B2(n1123), .ZN(
        n71120) );
  OAI22_X1 U22023 ( .A1(n23916), .A2(n1129), .B1(n22045), .B2(n1121), .ZN(
        n71100) );
  OAI22_X1 U22024 ( .A1(n23868), .A2(n1127), .B1(n22081), .B2(n1119), .ZN(
        n71080) );
  OAI22_X1 U22025 ( .A1(n25224), .A2(n1125), .B1(n22117), .B2(n1117), .ZN(
        n71060) );
  OAI22_X1 U22026 ( .A1(n23829), .A2(n1123), .B1(n21991), .B2(n27915), .ZN(
        n71040) );
  INV_X1 U22027 ( .A(sram_rdata_d0[1]), .ZN(n27915) );
  OAI22_X1 U22028 ( .A1(n23903), .A2(n1121), .B1(n22027), .B2(n27913), .ZN(
        n71020) );
  INV_X1 U22029 ( .A(sram_rdata_d0[3]), .ZN(n27913) );
  OAI22_X1 U22030 ( .A1(n23855), .A2(n1119), .B1(n22063), .B2(n27911), .ZN(
        n71000) );
  INV_X1 U22031 ( .A(sram_rdata_d0[5]), .ZN(n27911) );
  OAI22_X1 U22032 ( .A1(n25235), .A2(n1117), .B1(n22099), .B2(n27909), .ZN(
        n70980) );
  INV_X1 U22033 ( .A(sram_rdata_d0[7]), .ZN(n27909) );
  OAI22_X1 U22034 ( .A1(n23788), .A2(n15854), .B1(n21722), .B2(n1107), .ZN(
        n7088) );
  OAI22_X1 U22035 ( .A1(n20816), .A2(n15868), .B1(n21738), .B2(n1105), .ZN(
        n7086) );
  OAI22_X1 U22036 ( .A1(n20840), .A2(n15882), .B1(n21754), .B2(n1103), .ZN(
        n7084) );
  OAI22_X1 U22037 ( .A1(n19057), .A2(n15896), .B1(n21770), .B2(n1101), .ZN(
        n7082) );
  OAI22_X1 U22038 ( .A1(n23751), .A2(n1107), .B1(n22138), .B2(n1099), .ZN(
        n7080) );
  OAI22_X1 U22039 ( .A1(n23892), .A2(n1105), .B1(n22183), .B2(n1097), .ZN(
        n7078) );
  OAI22_X1 U22040 ( .A1(n23844), .A2(n1103), .B1(n22232), .B2(n1095), .ZN(
        n7076) );
  OAI22_X1 U22041 ( .A1(n25234), .A2(n1101), .B1(n23586), .B2(n1093), .ZN(
        n7074) );
  OAI22_X1 U22042 ( .A1(n23812), .A2(n1099), .B1(n21725), .B2(n1091), .ZN(
        n7072) );
  OAI22_X1 U22043 ( .A1(n20678), .A2(n1097), .B1(n21741), .B2(n1089), .ZN(
        n7070) );
  OAI22_X1 U22044 ( .A1(n20646), .A2(n1095), .B1(n21757), .B2(n1087), .ZN(
        n70680) );
  OAI22_X1 U22045 ( .A1(n25238), .A2(n1093), .B1(n21773), .B2(n1085), .ZN(
        n70660) );
  OAI22_X1 U22046 ( .A1(n23772), .A2(n1091), .B1(n21661), .B2(n1083), .ZN(
        n70640) );
  OAI22_X1 U22047 ( .A1(n20818), .A2(n1089), .B1(n21669), .B2(n1081), .ZN(
        n70620) );
  OAI22_X1 U22048 ( .A1(n20842), .A2(n1087), .B1(n21677), .B2(n1079), .ZN(
        n70600) );
  OAI22_X1 U22049 ( .A1(n25360), .A2(n1085), .B1(n21685), .B2(n1077), .ZN(
        n70580) );
  OAI22_X1 U22050 ( .A1(n23835), .A2(n1083), .B1(n22343), .B2(n1075), .ZN(
        n70560) );
  OAI22_X1 U22051 ( .A1(n24845), .A2(n1081), .B1(n22367), .B2(n1073), .ZN(
        n70540) );
  OAI22_X1 U22052 ( .A1(n24828), .A2(n1079), .B1(n22391), .B2(n1071), .ZN(
        n70520) );
  OAI22_X1 U22053 ( .A1(n20765), .A2(n1077), .B1(n22415), .B2(n1069), .ZN(
        n70500) );
  OAI22_X1 U22054 ( .A1(n23796), .A2(n1075), .B1(n21693), .B2(n1067), .ZN(
        n70480) );
  OAI22_X1 U22055 ( .A1(n20820), .A2(n1073), .B1(n21701), .B2(n1065), .ZN(
        n7046) );
  OAI22_X1 U22056 ( .A1(n20844), .A2(n1071), .B1(n21709), .B2(n1063), .ZN(
        n7044) );
  OAI22_X1 U22057 ( .A1(n25348), .A2(n1069), .B1(n24369), .B2(n1061), .ZN(
        n7042) );
  OAI22_X1 U22058 ( .A1(n23819), .A2(n1067), .B1(n22152), .B2(n27907), .ZN(
        n7040) );
  INV_X1 U22059 ( .A(sram_rdata_d0[9]), .ZN(n27907) );
  OAI22_X1 U22060 ( .A1(n24847), .A2(n1065), .B1(n22197), .B2(n27905), .ZN(
        n7038) );
  INV_X1 U22061 ( .A(sram_rdata_d0[11]), .ZN(n27905) );
  OAI22_X1 U22062 ( .A1(n24830), .A2(n1063), .B1(n22244), .B2(n27903), .ZN(
        n7036) );
  INV_X1 U22063 ( .A(sram_rdata_d0[13]), .ZN(n27903) );
  OAI22_X1 U22064 ( .A1(n19098), .A2(n1061), .B1(n22279), .B2(n27901), .ZN(
        n7034) );
  INV_X1 U22065 ( .A(sram_rdata_d0[15]), .ZN(n27901) );
  OAI22_X1 U22066 ( .A1(n23758), .A2(n16174), .B1(n22003), .B2(n1051), .ZN(
        n70240) );
  OAI22_X1 U22067 ( .A1(n20657), .A2(n16188), .B1(n22039), .B2(n1049), .ZN(
        n70220) );
  OAI22_X1 U22068 ( .A1(n20624), .A2(n16202), .B1(n22075), .B2(n1047), .ZN(
        n70200) );
  OAI22_X1 U22069 ( .A1(n24116), .A2(n16216), .B1(n22111), .B2(n1045), .ZN(
        n70180) );
  OAI22_X1 U22070 ( .A1(n23778), .A2(n1051), .B1(n22007), .B2(n1043), .ZN(
        n70160) );
  OAI22_X1 U22071 ( .A1(n24852), .A2(n1049), .B1(n22043), .B2(n1041), .ZN(
        n7014) );
  OAI22_X1 U22072 ( .A1(n24836), .A2(n1047), .B1(n22079), .B2(n1039), .ZN(
        n7012) );
  OAI22_X1 U22073 ( .A1(n24140), .A2(n1045), .B1(n22115), .B2(n1037), .ZN(
        n7010) );
  OAI22_X1 U22074 ( .A1(n23766), .A2(n1043), .B1(n22337), .B2(n1035), .ZN(
        n7008) );
  OAI22_X1 U22075 ( .A1(n20834), .A2(n1041), .B1(n22361), .B2(n1033), .ZN(
        n7006) );
  OAI22_X1 U22076 ( .A1(n20859), .A2(n1039), .B1(n22385), .B2(n1031), .ZN(
        n7004) );
  OAI22_X1 U22077 ( .A1(n24983), .A2(n1037), .B1(n22409), .B2(n1029), .ZN(
        n7002) );
  OAI22_X1 U22078 ( .A1(n23802), .A2(n1035), .B1(n22157), .B2(n1027), .ZN(
        n7000) );
  OAI22_X1 U22079 ( .A1(n24848), .A2(n1033), .B1(n22203), .B2(n1025), .ZN(
        n6998) );
  OAI22_X1 U22080 ( .A1(n24831), .A2(n1031), .B1(n22235), .B2(n1023), .ZN(
        n6996) );
  OAI22_X1 U22081 ( .A1(n24128), .A2(n1029), .B1(n22267), .B2(n1021), .ZN(
        n6994) );
  OAI22_X1 U22082 ( .A1(n23783), .A2(n1027), .B1(n21719), .B2(n1019), .ZN(
        n6992) );
  OAI22_X1 U22083 ( .A1(n24853), .A2(n1025), .B1(n21735), .B2(n1017), .ZN(
        n6990) );
  OAI22_X1 U22084 ( .A1(n24837), .A2(n1023), .B1(n21751), .B2(n1015), .ZN(
        n6988) );
  OAI22_X1 U22085 ( .A1(n24975), .A2(n1021), .B1(n21767), .B2(n1013), .ZN(
        n6986) );
  OAI22_X1 U22086 ( .A1(n23825), .A2(n1019), .B1(n21989), .B2(n1011), .ZN(
        n6984) );
  OAI22_X1 U22087 ( .A1(n20664), .A2(n1017), .B1(n22025), .B2(n1009), .ZN(
        n6982) );
  OAI22_X1 U22088 ( .A1(n20631), .A2(n1015), .B1(n22061), .B2(n1007), .ZN(
        n6980) );
  OAI22_X1 U22089 ( .A1(n24110), .A2(n1013), .B1(n22097), .B2(n1005), .ZN(
        n6978) );
  OAI22_X1 U22090 ( .A1(n23807), .A2(n1011), .B1(n21723), .B2(n27899), .ZN(
        n69760) );
  INV_X1 U22091 ( .A(sram_rdata_d0[17]), .ZN(n27899) );
  OAI22_X1 U22092 ( .A1(n20673), .A2(n1009), .B1(n21739), .B2(n27897), .ZN(
        n69740) );
  INV_X1 U22093 ( .A(sram_rdata_d0[19]), .ZN(n27897) );
  OAI22_X1 U22094 ( .A1(n20641), .A2(n1007), .B1(n21755), .B2(n27895), .ZN(
        n69720) );
  INV_X1 U22095 ( .A(sram_rdata_d0[21]), .ZN(n27895) );
  OAI22_X1 U22096 ( .A1(n20768), .A2(n1005), .B1(n21771), .B2(n27893), .ZN(
        n69700) );
  INV_X1 U22097 ( .A(sram_rdata_d0[23]), .ZN(n27893) );
  OAI22_X1 U22098 ( .A1(n23748), .A2(n16494), .B1(n22134), .B2(n995), .ZN(
        n69600) );
  OAI22_X1 U22099 ( .A1(n24840), .A2(n16508), .B1(n22179), .B2(n993), .ZN(
        n69580) );
  OAI22_X1 U22100 ( .A1(n24823), .A2(n16522), .B1(n22229), .B2(n991), .ZN(
        n69560) );
  OAI22_X1 U22101 ( .A1(n24134), .A2(n16536), .B1(n24368), .B2(n989), .ZN(
        n6954) );
  OAI22_X1 U22102 ( .A1(n23789), .A2(n995), .B1(n21692), .B2(n987), .ZN(n6952)
         );
  OAI22_X1 U22103 ( .A1(n23932), .A2(n993), .B1(n21700), .B2(n985), .ZN(n6950)
         );
  OAI22_X1 U22104 ( .A1(n23884), .A2(n991), .B1(n21708), .B2(n983), .ZN(n6948)
         );
  OAI22_X1 U22105 ( .A1(n24122), .A2(n989), .B1(n24362), .B2(n981), .ZN(n6946)
         );
  OAI22_X1 U22106 ( .A1(n23813), .A2(n987), .B1(n21660), .B2(n979), .ZN(n6944)
         );
  OAI22_X1 U22107 ( .A1(n23920), .A2(n985), .B1(n21668), .B2(n977), .ZN(n6942)
         );
  OAI22_X1 U22108 ( .A1(n23872), .A2(n983), .B1(n21676), .B2(n975), .ZN(n6940)
         );
  OAI22_X1 U22109 ( .A1(n20778), .A2(n981), .B1(n21684), .B2(n973), .ZN(n69380) );
  OAI22_X1 U22110 ( .A1(n23831), .A2(n979), .B1(n22002), .B2(n971), .ZN(n69360) );
  OAI22_X1 U22111 ( .A1(n23908), .A2(n977), .B1(n22038), .B2(n969), .ZN(n69340) );
  OAI22_X1 U22112 ( .A1(n23860), .A2(n975), .B1(n22074), .B2(n967), .ZN(n69320) );
  OAI22_X1 U22113 ( .A1(n25348), .A2(n973), .B1(n22110), .B2(n965), .ZN(n69300) );
  OAI22_X1 U22114 ( .A1(n23838), .A2(n971), .B1(n22342), .B2(n963), .ZN(n69280) );
  OAI22_X1 U22115 ( .A1(n20665), .A2(n969), .B1(n22366), .B2(n961), .ZN(n69260) );
  OAI22_X1 U22116 ( .A1(n20632), .A2(n967), .B1(n22390), .B2(n959), .ZN(n69240) );
  OAI22_X1 U22117 ( .A1(n26674), .A2(n965), .B1(n22414), .B2(n957), .ZN(n6922)
         );
  OAI22_X1 U22118 ( .A1(n23753), .A2(n963), .B1(n22149), .B2(n955), .ZN(n6920)
         );
  OAI22_X1 U22119 ( .A1(n23896), .A2(n961), .B1(n22194), .B2(n953), .ZN(n6918)
         );
  OAI22_X1 U22120 ( .A1(n23848), .A2(n959), .B1(n22242), .B2(n951), .ZN(n6916)
         );
  OAI22_X1 U22121 ( .A1(n25232), .A2(n957), .B1(n22276), .B2(n949), .ZN(n6914)
         );
  OAI22_X1 U22122 ( .A1(n23759), .A2(n955), .B1(n22335), .B2(n27891), .ZN(
        n6912) );
  INV_X1 U22123 ( .A(sram_rdata_d0[25]), .ZN(n27891) );
  OAI22_X1 U22124 ( .A1(n20657), .A2(n953), .B1(n22359), .B2(n27889), .ZN(
        n6910) );
  INV_X1 U22125 ( .A(sram_rdata_d0[27]), .ZN(n27889) );
  OAI22_X1 U22126 ( .A1(n20624), .A2(n951), .B1(n22383), .B2(n27887), .ZN(
        n6908) );
  INV_X1 U22127 ( .A(sram_rdata_d0[29]), .ZN(n27887) );
  OAI22_X1 U22128 ( .A1(n20760), .A2(n949), .B1(n22407), .B2(n27885), .ZN(
        n6906) );
  INV_X1 U22129 ( .A(sram_rdata_d0[31]), .ZN(n27885) );
  NAND2_X1 U22130 ( .A1(n5299), .A2(n884), .ZN(n5297) );
  INV_X1 U22131 ( .A(n53990), .ZN(n27755) );
  AOI22_X1 U22132 ( .A1(n17583), .A2(n25343), .B1(n17595), .B2(n26079), .ZN(
        n53990) );
  INV_X1 U22133 ( .A(n4886), .ZN(n27743) );
  AOI22_X1 U22134 ( .A1(n17751), .A2(n23728), .B1(n17763), .B2(n21466), .ZN(
        n4886) );
  NAND3_X1 U22135 ( .A1(n53960), .A2(n53970), .A3(n53980), .ZN(
        mul_outcome[104]) );
  AOI221_X1 U22136 ( .B1(n26621), .B2(n17571), .C1(n21973), .C2(n17559), .A(
        n27755), .ZN(n53980) );
  AOI22_X1 U22137 ( .A1(n26380), .A2(n17619), .B1(n26369), .B2(n17607), .ZN(
        n53960) );
  AOI22_X1 U22138 ( .A1(n24925), .A2(n17643), .B1(n24934), .B2(n17631), .ZN(
        n53970) );
  NAND3_X1 U22139 ( .A1(n5404), .A2(n5405), .A3(n5406), .ZN(mul_outcome[102])
         );
  AOI221_X1 U22140 ( .B1(n25239), .B2(n17575), .C1(n26399), .C2(n17563), .A(
        n27757), .ZN(n5406) );
  AOI22_X1 U22141 ( .A1(n21599), .A2(n17623), .B1(n21605), .B2(n17611), .ZN(
        n5404) );
  AOI22_X1 U22142 ( .A1(n24927), .A2(n17647), .B1(n24936), .B2(n17635), .ZN(
        n5405) );
  NAND3_X1 U22143 ( .A1(n5412), .A2(n5413), .A3(n5414), .ZN(mul_outcome[100])
         );
  AOI221_X1 U22144 ( .B1(n22679), .B2(n17579), .C1(n23493), .C2(n17567), .A(
        n27759), .ZN(n5414) );
  AOI22_X1 U22145 ( .A1(n17117), .A2(n17627), .B1(n21603), .B2(n17615), .ZN(
        n5412) );
  AOI22_X1 U22146 ( .A1(n19082), .A2(n17651), .B1(n19083), .B2(n17639), .ZN(
        n5413) );
  AOI22_X1 U22147 ( .A1(n24928), .A2(matrix_mul_2D_4__0__0_), .B1(n24937), 
        .B2(matrix_mul_2D_4__1__0_), .ZN(n4780) );
  AOI22_X1 U22148 ( .A1(n24928), .A2(matrix_mul_2D_4__0__1_), .B1(n24937), 
        .B2(matrix_mul_2D_4__1__1_), .ZN(n4776) );
  AOI22_X1 U22149 ( .A1(n19302), .A2(matrix_mul_2D_4__0__2_), .B1(n19300), 
        .B2(matrix_mul_2D_4__1__2_), .ZN(n4772) );
  AOI22_X1 U22150 ( .A1(n25322), .A2(matrix_mul_2D_4__0__3_), .B1(n25324), 
        .B2(matrix_mul_2D_4__1__3_), .ZN(n4768) );
  AOI22_X1 U22151 ( .A1(n24168), .A2(matrix_mul_2D_4__0__4_), .B1(n24164), 
        .B2(matrix_mul_2D_4__1__4_), .ZN(n4764) );
  AOI22_X1 U22152 ( .A1(n19082), .A2(matrix_mul_2D_4__0__5_), .B1(n19083), 
        .B2(matrix_mul_2D_4__1__5_), .ZN(n4760) );
  AOI22_X1 U22153 ( .A1(n24165), .A2(matrix_mul_2D_4__0__6_), .B1(n24161), 
        .B2(matrix_mul_2D_4__1__6_), .ZN(n4752) );
  AOI22_X1 U22154 ( .A1(n25323), .A2(matrix_mul_2D_4__0__7_), .B1(n25325), 
        .B2(matrix_mul_2D_4__1__7_), .ZN(n47480) );
  AOI22_X1 U22155 ( .A1(n24925), .A2(matrix_mul_2D_4__0__8_), .B1(n24934), 
        .B2(matrix_mul_2D_4__1__8_), .ZN(n47440) );
  AOI22_X1 U22156 ( .A1(n24927), .A2(matrix_mul_2D_4__0__9_), .B1(n24936), 
        .B2(matrix_mul_2D_4__1__9_), .ZN(n47400) );
  AOI22_X1 U22157 ( .A1(n26714), .A2(matrix_mul_2D_4__0__10_), .B1(n26710), 
        .B2(matrix_mul_2D_4__1__10_), .ZN(n47360) );
  AOI22_X1 U22158 ( .A1(n24168), .A2(matrix_mul_2D_4__0__11_), .B1(n24164), 
        .B2(matrix_mul_2D_4__1__11_), .ZN(n47320) );
  AOI22_X1 U22159 ( .A1(n24924), .A2(matrix_mul_2D_4__0__12_), .B1(n24933), 
        .B2(matrix_mul_2D_4__1__12_), .ZN(n47280) );
  AOI22_X1 U22160 ( .A1(n25323), .A2(matrix_mul_2D_4__0__13_), .B1(n25325), 
        .B2(matrix_mul_2D_4__1__13_), .ZN(n4724) );
  AOI22_X1 U22161 ( .A1(n24167), .A2(matrix_mul_2D_4__0__14_), .B1(n24163), 
        .B2(matrix_mul_2D_4__1__14_), .ZN(n4718) );
  OAI22_X1 U22162 ( .A1(n11855), .A2(n23763), .B1(n21995), .B2(n1780), .ZN(
        n6897) );
  OAI21_X1 U22163 ( .B1(n24016), .B2(n17020), .A(n45510), .ZN(n6371) );
  AOI22_X1 U22164 ( .A1(N7993), .A2(n25218), .B1(N7960), .B2(n24040), .ZN(
        n45510) );
  OAI21_X1 U22165 ( .B1(n24020), .B2(n17025), .A(n45520), .ZN(n6372) );
  AOI22_X1 U22166 ( .A1(N7992), .A2(n25218), .B1(N7959), .B2(n24044), .ZN(
        n45520) );
  OAI21_X1 U22167 ( .B1(n24022), .B2(n17011), .A(n45530), .ZN(n6373) );
  AOI22_X1 U22168 ( .A1(N7991), .A2(n19055), .B1(N7958), .B2(n24046), .ZN(
        n45530) );
  OAI21_X1 U22169 ( .B1(n24016), .B2(n16794), .A(n45540), .ZN(n6374) );
  AOI22_X1 U22170 ( .A1(N7990), .A2(n19055), .B1(N7957), .B2(n24040), .ZN(
        n45540) );
  OAI21_X1 U22171 ( .B1(n22698), .B2(n16779), .A(n45550), .ZN(n6375) );
  AOI22_X1 U22172 ( .A1(N7989), .A2(n25217), .B1(N7956), .B2(n19282), .ZN(
        n45550) );
  OAI21_X1 U22173 ( .B1(n24019), .B2(n16784), .A(n45560), .ZN(n6376) );
  AOI22_X1 U22174 ( .A1(N7988), .A2(n25217), .B1(N7955), .B2(n24043), .ZN(
        n45560) );
  OAI21_X1 U22175 ( .B1(n24023), .B2(n17060), .A(n45570), .ZN(n6377) );
  AOI22_X1 U22176 ( .A1(N7987), .A2(n24444), .B1(N7954), .B2(n24047), .ZN(
        n45570) );
  OAI21_X1 U22177 ( .B1(n22697), .B2(n17065), .A(n45580), .ZN(n6378) );
  AOI22_X1 U22178 ( .A1(N7986), .A2(n24810), .B1(N7953), .B2(n22707), .ZN(
        n45580) );
  OAI21_X1 U22179 ( .B1(n26639), .B2(n17045), .A(n45590), .ZN(n6379) );
  AOI22_X1 U22180 ( .A1(N7985), .A2(n24811), .B1(N7952), .B2(n22708), .ZN(
        n45590) );
  OAI21_X1 U22181 ( .B1(n24020), .B2(n17050), .A(n45600), .ZN(n6380) );
  AOI22_X1 U22182 ( .A1(N7984), .A2(n24448), .B1(N7951), .B2(n24044), .ZN(
        n45600) );
  OAI21_X1 U22183 ( .B1(n24022), .B2(n17055), .A(n45610), .ZN(n6381) );
  AOI22_X1 U22184 ( .A1(N7983), .A2(n24445), .B1(N7950), .B2(n24046), .ZN(
        n45610) );
  OAI21_X1 U22185 ( .B1(n26639), .B2(n17030), .A(n45620), .ZN(n6382) );
  AOI22_X1 U22186 ( .A1(N7982), .A2(n24442), .B1(N7949), .B2(n26643), .ZN(
        n45620) );
  OAI21_X1 U22187 ( .B1(n19279), .B2(n17035), .A(n45630), .ZN(n6383) );
  AOI22_X1 U22188 ( .A1(N7981), .A2(n24441), .B1(N7948), .B2(n26643), .ZN(
        n45630) );
  OAI21_X1 U22189 ( .B1(n24019), .B2(n17040), .A(n45640), .ZN(n6384) );
  AOI22_X1 U22190 ( .A1(N7980), .A2(n24448), .B1(N7947), .B2(n24043), .ZN(
        n45640) );
  OAI21_X1 U22191 ( .B1(n24023), .B2(n17015), .A(n45650), .ZN(n6385) );
  AOI22_X1 U22192 ( .A1(N7979), .A2(n24447), .B1(N7946), .B2(n24047), .ZN(
        n45650) );
  OAI21_X1 U22193 ( .B1(n22702), .B2(n16799), .A(n3080), .ZN(n54260) );
  AOI22_X1 U22194 ( .A1(N2606), .A2(n25657), .B1(N2573), .B2(n19281), .ZN(
        n3080) );
  OAI21_X1 U22195 ( .B1(n24028), .B2(n16804), .A(n30810), .ZN(n54270) );
  AOI22_X1 U22196 ( .A1(N2605), .A2(n25658), .B1(N2572), .B2(n24036), .ZN(
        n30810) );
  OAI21_X1 U22197 ( .B1(n24030), .B2(n16789), .A(n30820), .ZN(n54280) );
  AOI22_X1 U22198 ( .A1(N2604), .A2(n25654), .B1(N2571), .B2(n24038), .ZN(
        n30820) );
  OAI21_X1 U22199 ( .B1(n24024), .B2(n16814), .A(n30830), .ZN(n54290) );
  AOI22_X1 U22200 ( .A1(N2603), .A2(n21393), .B1(N2570), .B2(n24032), .ZN(
        n30830) );
  OAI21_X1 U22201 ( .B1(n24024), .B2(n16809), .A(n30840), .ZN(n54300) );
  AOI22_X1 U22202 ( .A1(N2602), .A2(n21386), .B1(N2569), .B2(n24032), .ZN(
        n30840) );
  OAI21_X1 U22203 ( .B1(n24027), .B2(n16829), .A(n30850), .ZN(n54310) );
  AOI22_X1 U22204 ( .A1(N2601), .A2(n21386), .B1(N2568), .B2(n24035), .ZN(
        n30850) );
  OAI21_X1 U22205 ( .B1(n24031), .B2(n16824), .A(n30860), .ZN(n54320) );
  AOI22_X1 U22206 ( .A1(N2600), .A2(n19240), .B1(N2567), .B2(n24039), .ZN(
        n30860) );
  OAI21_X1 U22207 ( .B1(n22701), .B2(n16819), .A(n30870), .ZN(n54330) );
  AOI22_X1 U22208 ( .A1(N2599), .A2(n19241), .B1(N2566), .B2(n22704), .ZN(
        n30870) );
  OAI21_X1 U22209 ( .B1(n26641), .B2(n16844), .A(n30880), .ZN(n54340) );
  AOI22_X1 U22210 ( .A1(N2598), .A2(n19239), .B1(N2565), .B2(n22705), .ZN(
        n30880) );
  OAI21_X1 U22211 ( .B1(n24028), .B2(n16849), .A(n30890), .ZN(n54350) );
  AOI22_X1 U22212 ( .A1(N2597), .A2(n25657), .B1(N2564), .B2(n24036), .ZN(
        n30890) );
  OAI21_X1 U22213 ( .B1(n24030), .B2(n16834), .A(n30900), .ZN(n54360) );
  AOI22_X1 U22214 ( .A1(N2596), .A2(n25658), .B1(N2563), .B2(n24038), .ZN(
        n30900) );
  OAI21_X1 U22215 ( .B1(n26641), .B2(n16859), .A(n30910), .ZN(n54370) );
  AOI22_X1 U22216 ( .A1(N2595), .A2(n25654), .B1(N2562), .B2(n26642), .ZN(
        n30910) );
  OAI21_X1 U22217 ( .B1(n19280), .B2(n16864), .A(n30920), .ZN(n54380) );
  AOI22_X1 U22218 ( .A1(N2594), .A2(n21392), .B1(N2561), .B2(n26642), .ZN(
        n30920) );
  OAI21_X1 U22219 ( .B1(n24027), .B2(n16839), .A(n30930), .ZN(n5439) );
  AOI22_X1 U22220 ( .A1(N2593), .A2(n21395), .B1(N2560), .B2(n24035), .ZN(
        n30930) );
  OAI21_X1 U22221 ( .B1(n24031), .B2(n16873), .A(n30940), .ZN(n5440) );
  AOI22_X1 U22222 ( .A1(N2592), .A2(n21385), .B1(N2559), .B2(n24039), .ZN(
        n30940) );
  AOI22_X1 U22223 ( .A1(n17383), .A2(n21495), .B1(n17407), .B2(n23968), .ZN(
        n5216) );
  AOI22_X1 U22224 ( .A1(n17381), .A2(n25910), .B1(n17405), .B2(n23976), .ZN(
        n5212) );
  AOI22_X1 U22225 ( .A1(n17379), .A2(n25911), .B1(n17403), .B2(n17103), .ZN(
        n5208) );
  AOI22_X1 U22226 ( .A1(n17385), .A2(n26066), .B1(n17409), .B2(n26927), .ZN(
        n52200) );
  AOI22_X1 U22227 ( .A1(n17387), .A2(n26756), .B1(n17411), .B2(n22676), .ZN(
        n52240) );
  AOI22_X1 U22228 ( .A1(n17389), .A2(n25908), .B1(n17413), .B2(n23973), .ZN(
        n52280) );
  NOR3_X1 U22229 ( .A1(upper_bound[5]), .A2(upper_bound[4]), .A3(
        upper_bound[3]), .ZN(n54250) );
  XNOR2_X1 U22230 ( .A(n26967), .B(n536), .ZN(upper_bound[3]) );
  XNOR2_X1 U22231 ( .A(n458), .B(sub_127_aco_carry[4]), .ZN(upper_bound[4]) );
  XNOR2_X1 U22232 ( .A(n462), .B(sub_127_aco_carry[5]), .ZN(upper_bound[5]) );
  OAI22_X1 U22233 ( .A1(n2024), .A2(n21246), .B1(n2003), .B2(n21243), .ZN(
        n50010) );
  OAI22_X1 U22234 ( .A1(n2023), .A2(n20487), .B1(n2002), .B2(n21232), .ZN(
        n4993) );
  OAI22_X1 U22235 ( .A1(n2022), .A2(n19202), .B1(n2001), .B2(n19201), .ZN(
        n4984) );
  OAI22_X1 U22236 ( .A1(n2025), .A2(n21239), .B1(n2004), .B2(n21236), .ZN(
        n50050) );
  OAI22_X1 U22237 ( .A1(n2026), .A2(n19204), .B1(n2005), .B2(n19200), .ZN(
        n50090) );
  OAI22_X1 U22238 ( .A1(n2027), .A2(n19203), .B1(n2006), .B2(n21241), .ZN(
        n50130) );
  AOI22_X1 U22239 ( .A1(n17299), .A2(n22830), .B1(n17311), .B2(n24424), .ZN(
        n5117) );
  AOI22_X1 U22240 ( .A1(n17297), .A2(n26075), .B1(n17309), .B2(n20814), .ZN(
        n5113) );
  AOI22_X1 U22241 ( .A1(n17295), .A2(n26068), .B1(n17307), .B2(n26404), .ZN(
        n5109) );
  AOI22_X1 U22242 ( .A1(n17301), .A2(n17077), .B1(n17313), .B2(n26399), .ZN(
        n5121) );
  AOI22_X1 U22243 ( .A1(n17303), .A2(n26067), .B1(n17315), .B2(n24401), .ZN(
        n5125) );
  AOI22_X1 U22244 ( .A1(n17305), .A2(n19249), .B1(n17317), .B2(n21967), .ZN(
        n5129) );
  AND2_X1 U22245 ( .A1(n549), .A2(n54250), .ZN(n54220) );
  INV_X1 U22246 ( .A(n50840), .ZN(n27783) );
  AOI22_X1 U22247 ( .A1(n17895), .A2(n21510), .B1(n17919), .B2(n21875), .ZN(
        n50840) );
  INV_X1 U22248 ( .A(n51440), .ZN(n27788) );
  AOI22_X1 U22249 ( .A1(n17905), .A2(n21508), .B1(n17929), .B2(n21872), .ZN(
        n51440) );
  AOI22_X1 U22250 ( .A1(n27016), .A2(matrix_mul_2D_5__0__0_), .B1(n25185), 
        .B2(matrix_mul_2D_5__1__0_), .ZN(n53920) );
  AOI22_X1 U22251 ( .A1(n27017), .A2(matrix_mul_2D_5__0__1_), .B1(n25186), 
        .B2(matrix_mul_2D_5__1__1_), .ZN(n53880) );
  AOI22_X1 U22252 ( .A1(n27018), .A2(matrix_mul_2D_5__0__2_), .B1(n22895), 
        .B2(matrix_mul_2D_5__1__2_), .ZN(n5384) );
  AOI22_X1 U22253 ( .A1(n27019), .A2(matrix_mul_2D_5__0__3_), .B1(n25183), 
        .B2(matrix_mul_2D_5__1__3_), .ZN(n5380) );
  AOI22_X1 U22254 ( .A1(n27020), .A2(matrix_mul_2D_5__0__4_), .B1(n24746), 
        .B2(matrix_mul_2D_5__1__4_), .ZN(n5376) );
  AOI22_X1 U22255 ( .A1(n27021), .A2(matrix_mul_2D_5__0__5_), .B1(n24747), 
        .B2(matrix_mul_2D_5__1__5_), .ZN(n5368) );
  AOI22_X1 U22256 ( .A1(n27022), .A2(matrix_mul_2D_5__0__6_), .B1(n19052), 
        .B2(matrix_mul_2D_5__1__6_), .ZN(n5364) );
  AOI22_X1 U22257 ( .A1(n27023), .A2(matrix_mul_2D_5__0__7_), .B1(n27029), 
        .B2(matrix_mul_2D_5__1__7_), .ZN(n5360) );
  AOI22_X1 U22258 ( .A1(n27024), .A2(matrix_mul_2D_5__0__8_), .B1(n25187), 
        .B2(matrix_mul_2D_5__1__8_), .ZN(n53560) );
  AOI22_X1 U22259 ( .A1(n27022), .A2(matrix_mul_2D_5__0__9_), .B1(n25184), 
        .B2(matrix_mul_2D_5__1__9_), .ZN(n53520) );
  AOI22_X1 U22260 ( .A1(n27023), .A2(matrix_mul_2D_5__0__10_), .B1(n24746), 
        .B2(matrix_mul_2D_5__1__10_), .ZN(n53480) );
  AOI22_X1 U22261 ( .A1(n27024), .A2(matrix_mul_2D_5__0__11_), .B1(n25187), 
        .B2(matrix_mul_2D_5__1__11_), .ZN(n53440) );
  AOI22_X1 U22262 ( .A1(n27025), .A2(matrix_mul_2D_5__0__12_), .B1(n27027), 
        .B2(matrix_mul_2D_5__1__12_), .ZN(n53400) );
  AOI22_X1 U22263 ( .A1(n27025), .A2(matrix_mul_2D_5__0__13_), .B1(n22896), 
        .B2(matrix_mul_2D_5__1__13_), .ZN(n5336) );
  AOI22_X1 U22264 ( .A1(n27026), .A2(matrix_mul_2D_5__0__14_), .B1(n25185), 
        .B2(matrix_mul_2D_5__1__14_), .ZN(n5332) );
  AOI22_X1 U22265 ( .A1(n27100), .A2(matrix_mul_2D_3__0__0_), .B1(n21187), 
        .B2(matrix_mul_2D_3__1__0_), .ZN(n48770) );
  AOI22_X1 U22266 ( .A1(n27063), .A2(matrix_mul_2D_2__0__0_), .B1(n27076), 
        .B2(matrix_mul_2D_2__1__0_), .ZN(n49760) );
  AOI22_X1 U22267 ( .A1(n27101), .A2(matrix_mul_2D_3__0__1_), .B1(n19184), 
        .B2(matrix_mul_2D_3__1__1_), .ZN(n48730) );
  AOI22_X1 U22268 ( .A1(n27064), .A2(matrix_mul_2D_2__0__1_), .B1(n27077), 
        .B2(matrix_mul_2D_2__1__1_), .ZN(n49720) );
  AOI22_X1 U22269 ( .A1(n27102), .A2(matrix_mul_2D_3__0__2_), .B1(n25748), 
        .B2(matrix_mul_2D_3__1__2_), .ZN(n48690) );
  AOI22_X1 U22270 ( .A1(n27065), .A2(matrix_mul_2D_2__0__2_), .B1(n27078), 
        .B2(matrix_mul_2D_2__1__2_), .ZN(n49680) );
  AOI22_X1 U22271 ( .A1(n27103), .A2(matrix_mul_2D_3__0__3_), .B1(n25749), 
        .B2(matrix_mul_2D_3__1__3_), .ZN(n4865) );
  AOI22_X1 U22272 ( .A1(n27066), .A2(matrix_mul_2D_2__0__3_), .B1(n27079), 
        .B2(matrix_mul_2D_2__1__3_), .ZN(n49640) );
  AOI22_X1 U22273 ( .A1(n27104), .A2(matrix_mul_2D_3__0__4_), .B1(n21190), 
        .B2(matrix_mul_2D_3__1__4_), .ZN(n4861) );
  AOI22_X1 U22274 ( .A1(n27067), .A2(matrix_mul_2D_2__0__4_), .B1(n27082), 
        .B2(matrix_mul_2D_2__1__4_), .ZN(n4960) );
  AOI22_X1 U22275 ( .A1(n27105), .A2(matrix_mul_2D_3__0__5_), .B1(n25541), 
        .B2(matrix_mul_2D_3__1__5_), .ZN(n4857) );
  AOI22_X1 U22276 ( .A1(n27068), .A2(matrix_mul_2D_2__0__5_), .B1(n27080), 
        .B2(matrix_mul_2D_2__1__5_), .ZN(n4956) );
  AOI22_X1 U22277 ( .A1(n27106), .A2(matrix_mul_2D_3__0__6_), .B1(n25536), 
        .B2(matrix_mul_2D_3__1__6_), .ZN(n4853) );
  AOI22_X1 U22278 ( .A1(n27069), .A2(matrix_mul_2D_2__0__6_), .B1(n22963), 
        .B2(matrix_mul_2D_2__1__6_), .ZN(n4952) );
  AOI22_X1 U22279 ( .A1(n27107), .A2(matrix_mul_2D_3__0__7_), .B1(n25749), 
        .B2(matrix_mul_2D_3__1__7_), .ZN(n4845) );
  AOI22_X1 U22280 ( .A1(n27070), .A2(matrix_mul_2D_2__0__7_), .B1(n22962), 
        .B2(matrix_mul_2D_2__1__7_), .ZN(n4948) );
  AOI22_X1 U22281 ( .A1(n27108), .A2(matrix_mul_2D_3__0__8_), .B1(n21179), 
        .B2(matrix_mul_2D_3__1__8_), .ZN(n4841) );
  AOI22_X1 U22282 ( .A1(n27071), .A2(matrix_mul_2D_2__0__8_), .B1(n27081), 
        .B2(matrix_mul_2D_2__1__8_), .ZN(n4940) );
  AOI22_X1 U22283 ( .A1(n27106), .A2(matrix_mul_2D_3__0__9_), .B1(n21190), 
        .B2(matrix_mul_2D_3__1__9_), .ZN(n48370) );
  AOI22_X1 U22284 ( .A1(n27069), .A2(matrix_mul_2D_2__0__9_), .B1(n27084), 
        .B2(matrix_mul_2D_2__1__9_), .ZN(n4936) );
  AOI22_X1 U22285 ( .A1(n27107), .A2(matrix_mul_2D_3__0__10_), .B1(n21178), 
        .B2(matrix_mul_2D_3__1__10_), .ZN(n48330) );
  AOI22_X1 U22286 ( .A1(n27070), .A2(matrix_mul_2D_2__0__10_), .B1(n22962), 
        .B2(matrix_mul_2D_2__1__10_), .ZN(n4932) );
  AOI22_X1 U22287 ( .A1(n27108), .A2(matrix_mul_2D_3__0__11_), .B1(n25747), 
        .B2(matrix_mul_2D_3__1__11_), .ZN(n48290) );
  AOI22_X1 U22288 ( .A1(n27071), .A2(matrix_mul_2D_2__0__11_), .B1(n27081), 
        .B2(matrix_mul_2D_2__1__11_), .ZN(n4928) );
  AOI22_X1 U22289 ( .A1(n22965), .A2(matrix_mul_2D_3__0__12_), .B1(n25746), 
        .B2(matrix_mul_2D_3__1__12_), .ZN(n48250) );
  AOI22_X1 U22290 ( .A1(n22966), .A2(matrix_mul_2D_3__0__13_), .B1(n25541), 
        .B2(matrix_mul_2D_3__1__13_), .ZN(n48210) );
  AOI22_X1 U22291 ( .A1(n22965), .A2(matrix_mul_2D_3__0__14_), .B1(n21189), 
        .B2(matrix_mul_2D_3__1__14_), .ZN(n4815) );
  OAI21_X1 U22292 ( .B1(n26355), .B2(n7419), .A(n4415), .ZN(n6294) );
  AOI22_X1 U22293 ( .A1(N7473), .A2(n21849), .B1(N7440), .B2(n25884), .ZN(
        n4415) );
  OAI21_X1 U22294 ( .B1(n21583), .B2(n7857), .A(n4255), .ZN(n61890) );
  AOI22_X1 U22295 ( .A1(N6875), .A2(n25997), .B1(N6842), .B2(n21276), .ZN(
        n4255) );
  OAI21_X1 U22296 ( .B1(n26346), .B2(n8018), .A(n42070), .ZN(n61590) );
  AOI22_X1 U22297 ( .A1(N6701), .A2(n21858), .B1(N6668), .B2(n25858), .ZN(
        n42070) );
  OAI21_X1 U22298 ( .B1(n21585), .B2(n8392), .A(n4094), .ZN(n6084) );
  AOI22_X1 U22299 ( .A1(N6262), .A2(n24265), .B1(N6229), .B2(n25889), .ZN(
        n4094) );
  OAI21_X1 U22300 ( .B1(n21555), .B2(n8552), .A(n40500), .ZN(n6054) );
  AOI22_X1 U22301 ( .A1(N6094), .A2(n21469), .B1(N6061), .B2(n25580), .ZN(
        n40500) );
  OAI21_X1 U22302 ( .B1(n21557), .B2(n9086), .A(n38890), .ZN(n5949) );
  AOI22_X1 U22303 ( .A1(N5508), .A2(n24253), .B1(N5475), .B2(n25862), .ZN(
        n38890) );
  OAI21_X1 U22304 ( .B1(n21917), .B2(n9486), .A(n3773), .ZN(n5874) );
  AOI22_X1 U22305 ( .A1(N5077), .A2(n21845), .B1(N5044), .B2(n24788), .ZN(
        n3773) );
  OAI21_X1 U22306 ( .B1(n21902), .B2(n9619), .A(n3729), .ZN(n58440) );
  AOI22_X1 U22307 ( .A1(N4903), .A2(n26071), .B1(N4870), .B2(n21261), .ZN(
        n3729) );
  OAI21_X1 U22308 ( .B1(n26123), .B2(n9993), .A(n3614), .ZN(n57690) );
  AOI22_X1 U22309 ( .A1(N4465), .A2(n22852), .B1(N4432), .B2(n25897), .ZN(
        n3614) );
  OAI21_X1 U22310 ( .B1(n21905), .B2(n10154), .A(n3570), .ZN(n5739) );
  AOI22_X1 U22311 ( .A1(N4297), .A2(n21853), .B1(N4264), .B2(n22891), .ZN(
        n3570) );
  OAI21_X1 U22312 ( .B1(n26124), .B2(n10554), .A(n34570), .ZN(n5664) );
  AOI22_X1 U22313 ( .A1(N3872), .A2(n21483), .B1(N3839), .B2(n22882), .ZN(
        n34570) );
  OAI21_X1 U22314 ( .B1(n26109), .B2(n10712), .A(n3410), .ZN(n5634) );
  AOI22_X1 U22315 ( .A1(N3701), .A2(n22845), .B1(N3668), .B2(n25878), .ZN(
        n3410) );
  OAI21_X1 U22316 ( .B1(n261101), .B2(n11257), .A(n3250), .ZN(n5529) );
  AOI22_X1 U22317 ( .A1(N3115), .A2(n21493), .B1(N3082), .B2(n24751), .ZN(
        n3250) );
  AOI22_X1 U22318 ( .A1(n26377), .A2(matrix_mul_2D_4__2__0_), .B1(n26366), 
        .B2(matrix_mul_2D_4__3__0_), .ZN(n4779) );
  AOI22_X1 U22319 ( .A1(n26130), .A2(matrix_mul_2D_4__2__1_), .B1(n26133), 
        .B2(matrix_mul_2D_4__3__1_), .ZN(n4775) );
  AOI22_X1 U22320 ( .A1(n26131), .A2(matrix_mul_2D_4__2__2_), .B1(n26134), 
        .B2(matrix_mul_2D_4__3__2_), .ZN(n4771) );
  AOI22_X1 U22321 ( .A1(n21948), .A2(matrix_mul_2D_4__2__3_), .B1(n21939), 
        .B2(matrix_mul_2D_4__3__3_), .ZN(n4767) );
  AOI22_X1 U22322 ( .A1(n17117), .A2(matrix_mul_2D_4__2__4_), .B1(n21606), 
        .B2(matrix_mul_2D_4__3__4_), .ZN(n4763) );
  AOI22_X1 U22323 ( .A1(n21597), .A2(matrix_mul_2D_4__2__5_), .B1(n21603), 
        .B2(matrix_mul_2D_4__3__5_), .ZN(n4759) );
  AOI22_X1 U22324 ( .A1(n21599), .A2(matrix_mul_2D_4__2__6_), .B1(n21605), 
        .B2(matrix_mul_2D_4__3__6_), .ZN(n4751) );
  AOI22_X1 U22325 ( .A1(n26380), .A2(matrix_mul_2D_4__2__7_), .B1(n26369), 
        .B2(matrix_mul_2D_4__3__7_), .ZN(n47470) );
  AOI22_X1 U22326 ( .A1(n26379), .A2(matrix_mul_2D_4__2__8_), .B1(n26368), 
        .B2(matrix_mul_2D_4__3__8_), .ZN(n47430) );
  AOI22_X1 U22327 ( .A1(n26130), .A2(matrix_mul_2D_4__2__9_), .B1(n26133), 
        .B2(matrix_mul_2D_4__3__9_), .ZN(n47390) );
  AOI22_X1 U22328 ( .A1(n26131), .A2(matrix_mul_2D_4__2__10_), .B1(n26134), 
        .B2(matrix_mul_2D_4__3__10_), .ZN(n47350) );
  AOI22_X1 U22329 ( .A1(n21947), .A2(matrix_mul_2D_4__2__11_), .B1(n21938), 
        .B2(matrix_mul_2D_4__3__11_), .ZN(n47310) );
  AOI22_X1 U22330 ( .A1(n21597), .A2(matrix_mul_2D_4__2__12_), .B1(n21939), 
        .B2(matrix_mul_2D_4__3__12_), .ZN(n4727) );
  AOI22_X1 U22331 ( .A1(n21596), .A2(matrix_mul_2D_4__2__13_), .B1(n21602), 
        .B2(matrix_mul_2D_4__3__13_), .ZN(n4723) );
  AOI22_X1 U22332 ( .A1(n21600), .A2(matrix_mul_2D_4__2__14_), .B1(n21606), 
        .B2(matrix_mul_2D_4__3__14_), .ZN(n4717) );
  OAI21_X1 U22333 ( .B1(n23705), .B2(n2986), .A(n4427), .ZN(n6296) );
  AOI22_X1 U22334 ( .A1(N7575), .A2(n25796), .B1(N7542), .B2(n23298), .ZN(
        n4427) );
  OAI21_X1 U22335 ( .B1(n25162), .B2(n29900), .A(n4428), .ZN(n6297) );
  AOI22_X1 U22336 ( .A1(N7574), .A2(n25801), .B1(N7541), .B2(n23141), .ZN(
        n4428) );
  OAI21_X1 U22337 ( .B1(n19104), .B2(n29940), .A(n4429), .ZN(n6298) );
  AOI22_X1 U22338 ( .A1(N7573), .A2(n25808), .B1(N7540), .B2(n24455), .ZN(
        n4429) );
  OAI21_X1 U22339 ( .B1(n25150), .B2(n29980), .A(n4430), .ZN(n6299) );
  AOI22_X1 U22340 ( .A1(N7572), .A2(n25825), .B1(N7539), .B2(n21635), .ZN(
        n4430) );
  OAI21_X1 U22341 ( .B1(n25147), .B2(n30020), .A(n44310), .ZN(n6300) );
  AOI22_X1 U22342 ( .A1(N7571), .A2(n25829), .B1(N7538), .B2(n20602), .ZN(
        n44310) );
  OAI21_X1 U22343 ( .B1(n23710), .B2(n3006), .A(n44320), .ZN(n6301) );
  AOI22_X1 U22344 ( .A1(N7570), .A2(n27186), .B1(N7537), .B2(n21645), .ZN(
        n44320) );
  OAI21_X1 U22345 ( .B1(n23716), .B2(n3010), .A(n44330), .ZN(n6302) );
  AOI22_X1 U22346 ( .A1(N7569), .A2(n25817), .B1(N7536), .B2(n21654), .ZN(
        n44330) );
  OAI21_X1 U22347 ( .B1(n26576), .B2(n3018), .A(n44350), .ZN(n6304) );
  AOI22_X1 U22348 ( .A1(N7567), .A2(n25814), .B1(N7534), .B2(n25992), .ZN(
        n44350) );
  OAI21_X1 U22349 ( .B1(n26571), .B2(n30220), .A(n44360), .ZN(n6305) );
  AOI22_X1 U22350 ( .A1(N7566), .A2(n27182), .B1(N7533), .B2(n24800), .ZN(
        n44360) );
  OAI21_X1 U22351 ( .B1(n19105), .B2(n30260), .A(n44370), .ZN(n6306) );
  AOI22_X1 U22352 ( .A1(N7565), .A2(n27179), .B1(N7532), .B2(n24453), .ZN(
        n44370) );
  OAI21_X1 U22353 ( .B1(n19038), .B2(n30300), .A(n44380), .ZN(n6307) );
  AOI22_X1 U22354 ( .A1(N7564), .A2(n25844), .B1(N7531), .B2(n25076), .ZN(
        n44380) );
  OAI21_X1 U22355 ( .B1(n19043), .B2(n30340), .A(n44390), .ZN(n6308) );
  AOI22_X1 U22356 ( .A1(N7563), .A2(n25850), .B1(N7530), .B2(n24449), .ZN(
        n44390) );
  OAI21_X1 U22357 ( .B1(n26575), .B2(n30380), .A(n44400), .ZN(n6309) );
  AOI22_X1 U22358 ( .A1(N7562), .A2(n25856), .B1(N7529), .B2(n26157), .ZN(
        n44400) );
  OAI21_X1 U22359 ( .B1(n26582), .B2(n3043), .A(n44410), .ZN(n6310) );
  AOI22_X1 U22360 ( .A1(N7561), .A2(n19316), .B1(N7528), .B2(n21652), .ZN(
        n44410) );
  OAI21_X1 U22361 ( .B1(n25159), .B2(n77380), .A(n42640), .ZN(n61910) );
  AOI22_X1 U22362 ( .A1(N6970), .A2(n25824), .B1(N6937), .B2(n23297), .ZN(
        n42640) );
  OAI21_X1 U22363 ( .B1(n25154), .B2(n77420), .A(n42650), .ZN(n61920) );
  AOI22_X1 U22364 ( .A1(N6969), .A2(n25828), .B1(N6936), .B2(n24802), .ZN(
        n42650) );
  OAI21_X1 U22365 ( .B1(n25153), .B2(n77460), .A(n42660), .ZN(n61930) );
  AOI22_X1 U22366 ( .A1(N6968), .A2(n22910), .B1(N6935), .B2(n21648), .ZN(
        n42660) );
  OAI21_X1 U22367 ( .B1(n19038), .B2(n7750), .A(n42670), .ZN(n61940) );
  AOI22_X1 U22368 ( .A1(N6967), .A2(n27183), .B1(N6934), .B2(n26163), .ZN(
        n42670) );
  OAI21_X1 U22369 ( .B1(n22524), .B2(n7754), .A(n42680), .ZN(n61950) );
  AOI22_X1 U22370 ( .A1(N6966), .A2(n25811), .B1(N6933), .B2(n24455), .ZN(
        n42680) );
  OAI21_X1 U22371 ( .B1(n26579), .B2(n7758), .A(n42690), .ZN(n61960) );
  AOI22_X1 U22372 ( .A1(N6965), .A2(n25813), .B1(N6932), .B2(n21459), .ZN(
        n42690) );
  OAI21_X1 U22373 ( .B1(n26570), .B2(n7766), .A(n42710), .ZN(n61980) );
  AOI22_X1 U22374 ( .A1(N6963), .A2(n25799), .B1(N6930), .B2(n21653), .ZN(
        n42710) );
  OAI21_X1 U22375 ( .B1(n25155), .B2(n7770), .A(n42720), .ZN(n61990) );
  AOI22_X1 U22376 ( .A1(N6962), .A2(n25849), .B1(N6929), .B2(n24456), .ZN(
        n42720) );
  OAI21_X1 U22377 ( .B1(n25157), .B2(n7774), .A(n42730), .ZN(n62000) );
  AOI22_X1 U22378 ( .A1(N6961), .A2(n25853), .B1(N6928), .B2(n21458), .ZN(
        n42730) );
  OAI21_X1 U22379 ( .B1(n19043), .B2(n77780), .A(n42740), .ZN(n62010) );
  AOI22_X1 U22380 ( .A1(N6960), .A2(n25857), .B1(N6927), .B2(n23139), .ZN(
        n42740) );
  OAI21_X1 U22381 ( .B1(n25369), .B2(n77820), .A(n42750), .ZN(n62020) );
  AOI22_X1 U22382 ( .A1(N6959), .A2(n22900), .B1(N6926), .B2(n23138), .ZN(
        n42750) );
  OAI21_X1 U22383 ( .B1(n23711), .B2(n77860), .A(n42760), .ZN(n6203) );
  AOI22_X1 U22384 ( .A1(N6958), .A2(n25553), .B1(N6925), .B2(n21635), .ZN(
        n42760) );
  OAI21_X1 U22385 ( .B1(n22527), .B2(n77900), .A(n42770), .ZN(n6204) );
  AOI22_X1 U22386 ( .A1(N6957), .A2(n24526), .B1(N6924), .B2(n23296), .ZN(
        n42770) );
  OAI21_X1 U22387 ( .B1(n25123), .B2(n8259), .A(n41030), .ZN(n6086) );
  AOI22_X1 U22388 ( .A1(N6364), .A2(n25821), .B1(N6331), .B2(n21651), .ZN(
        n41030) );
  OAI21_X1 U22389 ( .B1(n25371), .B2(n8263), .A(n41040), .ZN(n6087) );
  AOI22_X1 U22390 ( .A1(N6363), .A2(n25812), .B1(N6330), .B2(n23142), .ZN(
        n41040) );
  OAI21_X1 U22391 ( .B1(n26578), .B2(n8267), .A(n41050), .ZN(n6088) );
  AOI22_X1 U22392 ( .A1(N6362), .A2(n25815), .B1(N6329), .B2(n25993), .ZN(
        n41050) );
  OAI21_X1 U22393 ( .B1(n23715), .B2(n8275), .A(n41070), .ZN(n6090) );
  AOI22_X1 U22394 ( .A1(N6360), .A2(n25797), .B1(N6327), .B2(n24454), .ZN(
        n41070) );
  OAI21_X1 U22395 ( .B1(n22521), .B2(n8283), .A(n41090), .ZN(n6092) );
  AOI22_X1 U22396 ( .A1(N6358), .A2(n25852), .B1(N6325), .B2(n25991), .ZN(
        n41090) );
  OAI21_X1 U22397 ( .B1(n19045), .B2(n8287), .A(n41100), .ZN(n60930) );
  AOI22_X1 U22398 ( .A1(N6357), .A2(n25854), .B1(N6324), .B2(n20594), .ZN(
        n41100) );
  OAI21_X1 U22399 ( .B1(n25368), .B2(n8291), .A(n4111), .ZN(n60940) );
  AOI22_X1 U22400 ( .A1(N6356), .A2(n25848), .B1(N6323), .B2(n20593), .ZN(
        n4111) );
  OAI21_X1 U22401 ( .B1(n19044), .B2(n8295), .A(n4112), .ZN(n60950) );
  AOI22_X1 U22402 ( .A1(N6355), .A2(n24528), .B1(N6322), .B2(n21636), .ZN(
        n4112) );
  OAI21_X1 U22403 ( .B1(n23706), .B2(n8299), .A(n4113), .ZN(n60960) );
  AOI22_X1 U22404 ( .A1(N6354), .A2(n24529), .B1(N6321), .B2(n23299), .ZN(
        n4113) );
  OAI21_X1 U22405 ( .B1(n26575), .B2(n8303), .A(n4114), .ZN(n60970) );
  AOI22_X1 U22406 ( .A1(N6353), .A2(n25804), .B1(N6320), .B2(n21633), .ZN(
        n4114) );
  OAI21_X1 U22407 ( .B1(n26580), .B2(n8307), .A(n4115), .ZN(n60980) );
  AOI22_X1 U22408 ( .A1(N6352), .A2(n25808), .B1(N6319), .B2(n24450), .ZN(
        n4115) );
  OAI21_X1 U22409 ( .B1(n26573), .B2(n8316), .A(n4117), .ZN(n61000) );
  AOI22_X1 U22410 ( .A1(N6350), .A2(n25816), .B1(N6317), .B2(n20875), .ZN(
        n4117) );
  OAI21_X1 U22411 ( .B1(n23690), .B2(n8567), .A(n40110), .ZN(n60260) );
  AOI22_X1 U22412 ( .A1(N6028), .A2(n25762), .B1(N5995), .B2(n23284), .ZN(
        n40110) );
  OAI21_X1 U22413 ( .B1(n25144), .B2(n8572), .A(n40120), .ZN(n60270) );
  AOI22_X1 U22414 ( .A1(N6027), .A2(n25767), .B1(N5994), .B2(n23132), .ZN(
        n40120) );
  OAI21_X1 U22415 ( .B1(n19106), .B2(n8577), .A(n40130), .ZN(n60280) );
  AOI22_X1 U22416 ( .A1(N6026), .A2(n25774), .B1(N5993), .B2(n24462), .ZN(
        n40130) );
  OAI21_X1 U22417 ( .B1(n25132), .B2(n8582), .A(n40140), .ZN(n60290) );
  AOI22_X1 U22418 ( .A1(N6025), .A2(n25791), .B1(N5992), .B2(n21628), .ZN(
        n40140) );
  OAI21_X1 U22419 ( .B1(n25129), .B2(n8587), .A(n40150), .ZN(n60300) );
  AOI22_X1 U22420 ( .A1(N6024), .A2(n25795), .B1(N5991), .B2(n20603), .ZN(
        n40150) );
  OAI21_X1 U22421 ( .B1(n23695), .B2(n8592), .A(n40160), .ZN(n60310) );
  AOI22_X1 U22422 ( .A1(N6023), .A2(n27241), .B1(N5990), .B2(n21643), .ZN(
        n40160) );
  OAI21_X1 U22423 ( .B1(n23701), .B2(n8597), .A(n40170), .ZN(n60320) );
  AOI22_X1 U22424 ( .A1(N6022), .A2(n25783), .B1(N5989), .B2(n26152), .ZN(
        n40170) );
  OAI21_X1 U22425 ( .B1(n26563), .B2(n8607), .A(n40190), .ZN(n60340) );
  AOI22_X1 U22426 ( .A1(N6020), .A2(n25779), .B1(N5987), .B2(n25988), .ZN(
        n40190) );
  OAI21_X1 U22427 ( .B1(n26557), .B2(n8612), .A(n40200), .ZN(n6035) );
  AOI22_X1 U22428 ( .A1(N6019), .A2(n25765), .B1(N5986), .B2(n23128), .ZN(
        n40200) );
  OAI21_X1 U22429 ( .B1(n19107), .B2(n8617), .A(n40210), .ZN(n6036) );
  AOI22_X1 U22430 ( .A1(N6018), .A2(n27236), .B1(N5985), .B2(n24459), .ZN(
        n40210) );
  OAI21_X1 U22431 ( .B1(n19039), .B2(n8622), .A(n4022), .ZN(n6037) );
  AOI22_X1 U22432 ( .A1(N6017), .A2(n25830), .B1(N5984), .B2(n25082), .ZN(
        n4022) );
  OAI21_X1 U22433 ( .B1(n19040), .B2(n8627), .A(n4023), .ZN(n6038) );
  AOI22_X1 U22434 ( .A1(N6016), .A2(n25836), .B1(N5983), .B2(n24451), .ZN(
        n4023) );
  OAI21_X1 U22435 ( .B1(n26562), .B2(n8632), .A(n4024), .ZN(n6039) );
  AOI22_X1 U22436 ( .A1(N6015), .A2(n25842), .B1(N5982), .B2(n21642), .ZN(
        n4024) );
  OAI21_X1 U22437 ( .B1(n26569), .B2(n8636), .A(n4025), .ZN(n6040) );
  AOI22_X1 U22438 ( .A1(N6014), .A2(n27233), .B1(N5981), .B2(n21639), .ZN(
        n4025) );
  OAI21_X1 U22439 ( .B1(n25154), .B2(n8806), .A(n39420), .ZN(n59810) );
  AOI22_X1 U22440 ( .A1(N5768), .A2(n22916), .B1(N5735), .B2(n26156), .ZN(
        n39420) );
  OAI21_X1 U22441 ( .B1(n22524), .B2(n8810), .A(n3943), .ZN(n59820) );
  AOI22_X1 U22442 ( .A1(N5767), .A2(n27180), .B1(N5734), .B2(n26162), .ZN(
        n3943) );
  OAI21_X1 U22443 ( .B1(n26581), .B2(n8814), .A(n3944), .ZN(n59830) );
  AOI22_X1 U22444 ( .A1(N5766), .A2(n21419), .B1(N5733), .B2(n24800), .ZN(
        n3944) );
  OAI21_X1 U22445 ( .B1(n23711), .B2(n8822), .A(n3946), .ZN(n59850) );
  AOI22_X1 U22446 ( .A1(N5764), .A2(n25855), .B1(N5731), .B2(n23139), .ZN(
        n3946) );
  OAI21_X1 U22447 ( .B1(n26570), .B2(n8826), .A(n3947), .ZN(n59860) );
  AOI22_X1 U22448 ( .A1(N5763), .A2(n25845), .B1(N5730), .B2(n23142), .ZN(
        n3947) );
  OAI21_X1 U22449 ( .B1(n25148), .B2(n8830), .A(n3948), .ZN(n59870) );
  AOI22_X1 U22450 ( .A1(N5762), .A2(n25554), .B1(N5729), .B2(n23298), .ZN(
        n3948) );
  OAI21_X1 U22451 ( .B1(n25371), .B2(n8834), .A(n3949), .ZN(n59880) );
  AOI22_X1 U22452 ( .A1(N5761), .A2(n25551), .B1(N5728), .B2(n20600), .ZN(
        n3949) );
  OAI21_X1 U22453 ( .B1(n25156), .B2(n8838), .A(n3950), .ZN(n59890) );
  AOI22_X1 U22454 ( .A1(N5760), .A2(n25803), .B1(N5727), .B2(n26157), .ZN(
        n3950) );
  OAI21_X1 U22455 ( .B1(n26578), .B2(n8842), .A(n3951), .ZN(n59900) );
  AOI22_X1 U22456 ( .A1(N5759), .A2(n25807), .B1(N5726), .B2(n26163), .ZN(
        n3951) );
  OAI21_X1 U22457 ( .B1(n22528), .B2(n8846), .A(n3952), .ZN(n59910) );
  AOI22_X1 U22458 ( .A1(N5758), .A2(n25824), .B1(N5725), .B2(n26150), .ZN(
        n3952) );
  OAI21_X1 U22459 ( .B1(n23716), .B2(n8850), .A(n3953), .ZN(n59920) );
  AOI22_X1 U22460 ( .A1(N5757), .A2(n25828), .B1(N5724), .B2(n25076), .ZN(
        n3953) );
  OAI21_X1 U22461 ( .B1(n22521), .B2(n8858), .A(n3955), .ZN(n59940) );
  AOI22_X1 U22462 ( .A1(N5755), .A2(n25820), .B1(N5722), .B2(n23296), .ZN(
        n3955) );
  OAI21_X1 U22463 ( .B1(n25149), .B2(n8863), .A(n3956), .ZN(n59950) );
  AOI22_X1 U22464 ( .A1(N5754), .A2(n22907), .B1(N5721), .B2(n21646), .ZN(
        n3956) );
  OAI21_X1 U22465 ( .B1(n25141), .B2(n9101), .A(n3854), .ZN(n5921) );
  AOI22_X1 U22466 ( .A1(N5432), .A2(n25790), .B1(N5399), .B2(n23285), .ZN(
        n3854) );
  OAI21_X1 U22467 ( .B1(n25136), .B2(n9106), .A(n3855), .ZN(n5922) );
  AOI22_X1 U22468 ( .A1(N5431), .A2(n25794), .B1(N5398), .B2(n24801), .ZN(
        n3855) );
  OAI21_X1 U22469 ( .B1(n25135), .B2(n9111), .A(n3856), .ZN(n5923) );
  AOI22_X1 U22470 ( .A1(N5430), .A2(n22921), .B1(N5397), .B2(n21644), .ZN(
        n3856) );
  OAI21_X1 U22471 ( .B1(n19039), .B2(n9116), .A(n3857), .ZN(n5924) );
  AOI22_X1 U22472 ( .A1(N5429), .A2(n27238), .B1(N5396), .B2(n26153), .ZN(
        n3857) );
  OAI21_X1 U22473 ( .B1(n22515), .B2(n9121), .A(n3858), .ZN(n59250) );
  AOI22_X1 U22474 ( .A1(N5428), .A2(n25778), .B1(N5395), .B2(n24464), .ZN(
        n3858) );
  OAI21_X1 U22475 ( .B1(n26566), .B2(n9126), .A(n3859), .ZN(n59260) );
  AOI22_X1 U22476 ( .A1(N5427), .A2(n25780), .B1(N5394), .B2(n25989), .ZN(
        n3859) );
  OAI21_X1 U22477 ( .B1(n26556), .B2(n9136), .A(n3861), .ZN(n59280) );
  AOI22_X1 U22478 ( .A1(N5425), .A2(n27237), .B1(N5392), .B2(n26153), .ZN(
        n3861) );
  OAI21_X1 U22479 ( .B1(n25137), .B2(n9141), .A(n3862), .ZN(n59290) );
  AOI22_X1 U22480 ( .A1(N5424), .A2(n25835), .B1(N5391), .B2(n24461), .ZN(
        n3862) );
  OAI21_X1 U22481 ( .B1(n25139), .B2(n9146), .A(n3863), .ZN(n59300) );
  AOI22_X1 U22482 ( .A1(N5423), .A2(n25839), .B1(N5390), .B2(n21457), .ZN(
        n3863) );
  OAI21_X1 U22483 ( .B1(n19040), .B2(n9151), .A(n3864), .ZN(n59310) );
  AOI22_X1 U22484 ( .A1(N5422), .A2(n25843), .B1(N5389), .B2(n23130), .ZN(
        n3864) );
  OAI21_X1 U22485 ( .B1(n25373), .B2(n9156), .A(n3865), .ZN(n59320) );
  AOI22_X1 U22486 ( .A1(N5421), .A2(n22903), .B1(N5388), .B2(n23129), .ZN(
        n3865) );
  OAI21_X1 U22487 ( .B1(n23696), .B2(n9161), .A(n3866), .ZN(n59330) );
  AOI22_X1 U22488 ( .A1(N5420), .A2(n24532), .B1(N5387), .B2(n21627), .ZN(
        n3866) );
  OAI21_X1 U22489 ( .B1(n22518), .B2(n9166), .A(n3867), .ZN(n59340) );
  AOI22_X1 U22490 ( .A1(N5419), .A2(n24534), .B1(N5386), .B2(n20879), .ZN(
        n3867) );
  OAI21_X1 U22491 ( .B1(n26577), .B2(n9341), .A(n3782), .ZN(n5876) );
  AOI22_X1 U22492 ( .A1(N5182), .A2(n25853), .B1(N5149), .B2(n21458), .ZN(
        n3782) );
  OAI21_X1 U22493 ( .B1(n26582), .B2(n9346), .A(n3783), .ZN(n5877) );
  AOI22_X1 U22494 ( .A1(N5181), .A2(n25857), .B1(N5148), .B2(n21647), .ZN(
        n3783) );
  OAI21_X1 U22495 ( .B1(n23706), .B2(n9356), .A(n3785), .ZN(n5879) );
  AOI22_X1 U22496 ( .A1(N5179), .A2(n25554), .B1(N5146), .B2(n23137), .ZN(
        n3785) );
  OAI21_X1 U22497 ( .B1(n25124), .B2(n9361), .A(n3786), .ZN(n5880) );
  AOI22_X1 U22498 ( .A1(N5178), .A2(n24527), .B1(N5145), .B2(n25992), .ZN(
        n3786) );
  OAI21_X1 U22499 ( .B1(n25158), .B2(n9366), .A(n3787), .ZN(n5881) );
  AOI22_X1 U22500 ( .A1(N5177), .A2(n25804), .B1(N5144), .B2(n24456), .ZN(
        n3787) );
  OAI21_X1 U22501 ( .B1(n25161), .B2(n9371), .A(n3788), .ZN(n5882) );
  AOI22_X1 U22502 ( .A1(N5176), .A2(n25805), .B1(N5143), .B2(n24458), .ZN(
        n3788) );
  OAI21_X1 U22503 ( .B1(n25161), .B2(n9376), .A(n37890), .ZN(n5883) );
  AOI22_X1 U22504 ( .A1(N5175), .A2(n25822), .B1(N5142), .B2(n26150), .ZN(
        n37890) );
  OAI21_X1 U22505 ( .B1(n22525), .B2(n9381), .A(n37900), .ZN(n5884) );
  AOI22_X1 U22506 ( .A1(N5174), .A2(n25829), .B1(N5141), .B2(n20874), .ZN(
        n37900) );
  OAI21_X1 U22507 ( .B1(n26579), .B2(n9386), .A(n37910), .ZN(n5885) );
  AOI22_X1 U22508 ( .A1(N5173), .A2(n25818), .B1(N5140), .B2(n24806), .ZN(
        n37910) );
  OAI21_X1 U22509 ( .B1(n26573), .B2(n9396), .A(n37930), .ZN(n5887) );
  AOI22_X1 U22510 ( .A1(N5171), .A2(n25825), .B1(N5138), .B2(n23136), .ZN(
        n37930) );
  OAI21_X1 U22511 ( .B1(n25146), .B2(n9401), .A(n37940), .ZN(n58880) );
  AOI22_X1 U22512 ( .A1(N5170), .A2(n25826), .B1(N5137), .B2(n23137), .ZN(
        n37940) );
  OAI21_X1 U22513 ( .B1(n19104), .B2(n9406), .A(n37950), .ZN(n5889) );
  AOI22_X1 U22514 ( .A1(N5169), .A2(n25809), .B1(N5136), .B2(n26151), .ZN(
        n37950) );
  OAI21_X1 U22515 ( .B1(n25148), .B2(n9410), .A(n37960), .ZN(n5890) );
  AOI22_X1 U22516 ( .A1(N5168), .A2(n25815), .B1(N5135), .B2(n20597), .ZN(
        n37960) );
  OAI21_X1 U22517 ( .B1(n25125), .B2(n9635), .A(n3694), .ZN(n58160) );
  AOI22_X1 U22518 ( .A1(N4834), .A2(n25787), .B1(N4801), .B2(n21637), .ZN(
        n3694) );
  OAI21_X1 U22519 ( .B1(n25375), .B2(n9640), .A(n3695), .ZN(n58170) );
  AOI22_X1 U22520 ( .A1(N4833), .A2(n25778), .B1(N4800), .B2(n23133), .ZN(
        n3695) );
  OAI21_X1 U22521 ( .B1(n26565), .B2(n9645), .A(n3696), .ZN(n58180) );
  AOI22_X1 U22522 ( .A1(N4832), .A2(n25781), .B1(N4799), .B2(n21456), .ZN(
        n3696) );
  OAI21_X1 U22523 ( .B1(n23700), .B2(n9655), .A(n3698), .ZN(n58200) );
  AOI22_X1 U22524 ( .A1(N4830), .A2(n27235), .B1(N4797), .B2(n23127), .ZN(
        n3698) );
  OAI21_X1 U22525 ( .B1(n22512), .B2(n9665), .A(n37000), .ZN(n58220) );
  AOI22_X1 U22526 ( .A1(N4828), .A2(n25839), .B1(N4795), .B2(n25987), .ZN(
        n37000) );
  OAI21_X1 U22527 ( .B1(n19042), .B2(n9670), .A(n37010), .ZN(n58230) );
  AOI22_X1 U22528 ( .A1(N4827), .A2(n25840), .B1(N4794), .B2(n24798), .ZN(
        n37010) );
  OAI21_X1 U22529 ( .B1(n25372), .B2(n9675), .A(n37020), .ZN(n58240) );
  AOI22_X1 U22530 ( .A1(N4826), .A2(n25834), .B1(N4793), .B2(n20591), .ZN(
        n37020) );
  OAI21_X1 U22531 ( .B1(n19041), .B2(n9680), .A(n37030), .ZN(n58250) );
  AOI22_X1 U22532 ( .A1(N4825), .A2(n24535), .B1(N4792), .B2(n21627), .ZN(
        n37030) );
  OAI21_X1 U22533 ( .B1(n23691), .B2(n9685), .A(n37040), .ZN(n5826) );
  AOI22_X1 U22534 ( .A1(N4824), .A2(n24561), .B1(N4791), .B2(n24808), .ZN(
        n37040) );
  OAI21_X1 U22535 ( .B1(n26562), .B2(n9690), .A(n37050), .ZN(n5827) );
  AOI22_X1 U22536 ( .A1(N4823), .A2(n25770), .B1(N4790), .B2(n26146), .ZN(
        n37050) );
  OAI21_X1 U22537 ( .B1(n26567), .B2(n9695), .A(n37060), .ZN(n5828) );
  AOI22_X1 U22538 ( .A1(N4822), .A2(n25773), .B1(N4789), .B2(n23284), .ZN(
        n37060) );
  OAI21_X1 U22539 ( .B1(n26559), .B2(n9704), .A(n37080), .ZN(n5830) );
  AOI22_X1 U22540 ( .A1(N4820), .A2(n25782), .B1(N4787), .B2(n23287), .ZN(
        n37080) );
  OAI21_X1 U22541 ( .B1(n22527), .B2(n9874), .A(n36260), .ZN(n57710) );
  AOI22_X1 U22542 ( .A1(N4560), .A2(n25552), .B1(N4527), .B2(n24458), .ZN(
        n36260) );
  OAI21_X1 U22543 ( .B1(n26572), .B2(n9882), .A(n36280), .ZN(n57730) );
  AOI22_X1 U22544 ( .A1(N4558), .A2(n25802), .B1(N4525), .B2(n24457), .ZN(
        n36280) );
  OAI21_X1 U22545 ( .B1(n25370), .B2(n9886), .A(n36290), .ZN(n57740) );
  AOI22_X1 U22546 ( .A1(N4557), .A2(n25806), .B1(N4524), .B2(n23138), .ZN(
        n36290) );
  OAI21_X1 U22547 ( .B1(n25368), .B2(n9890), .A(n36300), .ZN(n5775) );
  AOI22_X1 U22548 ( .A1(N4556), .A2(n25823), .B1(N4523), .B2(n21634), .ZN(
        n36300) );
  OAI21_X1 U22549 ( .B1(n25150), .B2(n9894), .A(n36310), .ZN(n5776) );
  AOI22_X1 U22550 ( .A1(N4555), .A2(n25827), .B1(N4522), .B2(n20599), .ZN(
        n36310) );
  OAI21_X1 U22551 ( .B1(n22522), .B2(n9898), .A(n36320), .ZN(n5777) );
  AOI22_X1 U22552 ( .A1(N4554), .A2(n27185), .B1(N4521), .B2(n26151), .ZN(
        n36320) );
  OAI21_X1 U22553 ( .B1(n23710), .B2(n9902), .A(n36330), .ZN(n5778) );
  AOI22_X1 U22554 ( .A1(N4553), .A2(n27184), .B1(N4520), .B2(n24806), .ZN(
        n36330) );
  OAI21_X1 U22555 ( .B1(n23715), .B2(n9906), .A(n36340), .ZN(n5779) );
  AOI22_X1 U22556 ( .A1(N4552), .A2(n25812), .B1(N4519), .B2(n24802), .ZN(
        n36340) );
  OAI21_X1 U22557 ( .B1(n23705), .B2(n9914), .A(n36360), .ZN(n5781) );
  AOI22_X1 U22558 ( .A1(N4550), .A2(n25803), .B1(N4517), .B2(n24804), .ZN(
        n36360) );
  OAI21_X1 U22559 ( .B1(n25159), .B2(n9918), .A(n36370), .ZN(n5782) );
  AOI22_X1 U22560 ( .A1(N4549), .A2(n25807), .B1(N4516), .B2(n24804), .ZN(
        n36370) );
  OAI21_X1 U22561 ( .B1(n19105), .B2(n9922), .A(n36380), .ZN(n5783) );
  AOI22_X1 U22562 ( .A1(N4548), .A2(n22915), .B1(N4515), .B2(n21647), .ZN(
        n36380) );
  OAI21_X1 U22563 ( .B1(n25152), .B2(n9926), .A(n36390), .ZN(n5784) );
  AOI22_X1 U22564 ( .A1(N4547), .A2(n22913), .B1(N4514), .B2(n26162), .ZN(
        n36390) );
  OAI21_X1 U22565 ( .B1(n25123), .B2(n9931), .A(n36400), .ZN(n5785) );
  AOI22_X1 U22566 ( .A1(N4546), .A2(n27178), .B1(N4513), .B2(n24457), .ZN(
        n36400) );
  OAI21_X1 U22567 ( .B1(n25136), .B2(n10169), .A(n35350), .ZN(n5711) );
  AOI22_X1 U22568 ( .A1(N4221), .A2(n22927), .B1(N4188), .B2(n26154), .ZN(
        n35350) );
  OAI21_X1 U22569 ( .B1(n22515), .B2(n10174), .A(n35360), .ZN(n5712) );
  AOI22_X1 U22570 ( .A1(N4220), .A2(n25763), .B1(N4187), .B2(n21638), .ZN(
        n35360) );
  OAI21_X1 U22571 ( .B1(n26568), .B2(n10179), .A(n35370), .ZN(n5713) );
  AOI22_X1 U22572 ( .A1(N4219), .A2(n19317), .B1(N4186), .B2(n24462), .ZN(
        n35370) );
  OAI21_X1 U22573 ( .B1(n23696), .B2(n10189), .A(n35390), .ZN(n5715) );
  AOI22_X1 U22574 ( .A1(N4217), .A2(n25843), .B1(N4184), .B2(n23130), .ZN(
        n35390) );
  OAI21_X1 U22575 ( .B1(n26556), .B2(n10194), .A(n35400), .ZN(n5716) );
  AOI22_X1 U22576 ( .A1(N4216), .A2(n21416), .B1(N4183), .B2(n24459), .ZN(
        n35400) );
  OAI21_X1 U22577 ( .B1(n25130), .B2(n10199), .A(n35410), .ZN(n5717) );
  AOI22_X1 U22578 ( .A1(N4215), .A2(n24562), .B1(N4182), .B2(n23286), .ZN(
        n35410) );
  OAI21_X1 U22579 ( .B1(n25375), .B2(n10204), .A(n35420), .ZN(n5718) );
  AOI22_X1 U22580 ( .A1(N4214), .A2(n25549), .B1(N4181), .B2(n20595), .ZN(
        n35420) );
  OAI21_X1 U22581 ( .B1(n25138), .B2(n10209), .A(n35430), .ZN(n5719) );
  AOI22_X1 U22582 ( .A1(N4213), .A2(n25769), .B1(N4180), .B2(n26155), .ZN(
        n35430) );
  OAI21_X1 U22583 ( .B1(n26565), .B2(n10214), .A(n35440), .ZN(n5720) );
  AOI22_X1 U22584 ( .A1(N4212), .A2(n25774), .B1(N4179), .B2(n21640), .ZN(
        n35440) );
  OAI21_X1 U22585 ( .B1(n22519), .B2(n10219), .A(n35450), .ZN(n57210) );
  AOI22_X1 U22586 ( .A1(N4211), .A2(n25791), .B1(N4178), .B2(n21625), .ZN(
        n35450) );
  OAI21_X1 U22587 ( .B1(n23701), .B2(n10224), .A(n35460), .ZN(n57220) );
  AOI22_X1 U22588 ( .A1(N4210), .A2(n25795), .B1(N4177), .B2(n23286), .ZN(
        n35460) );
  OAI21_X1 U22589 ( .B1(n22512), .B2(n10234), .A(n35480), .ZN(n57240) );
  AOI22_X1 U22590 ( .A1(N4208), .A2(n25784), .B1(N4175), .B2(n20589), .ZN(
        n35480) );
  OAI21_X1 U22591 ( .B1(n25131), .B2(n10238), .A(n35490), .ZN(n57250) );
  AOI22_X1 U22592 ( .A1(N4207), .A2(n22919), .B1(N4174), .B2(n21641), .ZN(
        n35490) );
  OAI21_X1 U22593 ( .B1(n26564), .B2(n10739), .A(n33750), .ZN(n56060) );
  AOI22_X1 U22594 ( .A1(N3635), .A2(n25838), .B1(N3602), .B2(n21456), .ZN(
        n33750) );
  OAI21_X1 U22595 ( .B1(n26569), .B2(n10743), .A(n33760), .ZN(n5607) );
  AOI22_X1 U22596 ( .A1(N3634), .A2(n25841), .B1(N3601), .B2(n26155), .ZN(
        n33760) );
  OAI21_X1 U22597 ( .B1(n23691), .B2(n10751), .A(n33780), .ZN(n5609) );
  AOI22_X1 U22598 ( .A1(N3632), .A2(n24562), .B1(N3599), .B2(n24798), .ZN(
        n33780) );
  OAI21_X1 U22599 ( .B1(n25126), .B2(n10755), .A(n33790), .ZN(n5610) );
  AOI22_X1 U22600 ( .A1(N3631), .A2(n24531), .B1(N3598), .B2(n25988), .ZN(
        n33790) );
  OAI21_X1 U22601 ( .B1(n25140), .B2(n10759), .A(n33800), .ZN(n5611) );
  AOI22_X1 U22602 ( .A1(N3630), .A2(n25770), .B1(N3597), .B2(n24461), .ZN(
        n33800) );
  OAI21_X1 U22603 ( .B1(n25143), .B2(n10763), .A(n33810), .ZN(n5612) );
  AOI22_X1 U22604 ( .A1(N3629), .A2(n25771), .B1(N3596), .B2(n24464), .ZN(
        n33810) );
  OAI21_X1 U22605 ( .B1(n25143), .B2(n10767), .A(n33820), .ZN(n5613) );
  AOI22_X1 U22606 ( .A1(N3628), .A2(n25788), .B1(N3595), .B2(n26145), .ZN(
        n33820) );
  OAI21_X1 U22607 ( .B1(n22516), .B2(n10771), .A(n33830), .ZN(n5614) );
  AOI22_X1 U22608 ( .A1(N3627), .A2(n25794), .B1(N3594), .B2(n25082), .ZN(
        n33830) );
  OAI21_X1 U22609 ( .B1(n26566), .B2(n10775), .A(n33840), .ZN(n5615) );
  AOI22_X1 U22610 ( .A1(N3626), .A2(n27240), .B1(N3593), .B2(n20596), .ZN(
        n33840) );
  OAI21_X1 U22611 ( .B1(n26559), .B2(n10783), .A(n3386), .ZN(n5617) );
  AOI22_X1 U22612 ( .A1(N3624), .A2(n25790), .B1(N3591), .B2(n20592), .ZN(
        n3386) );
  OAI21_X1 U22613 ( .B1(n25128), .B2(n10787), .A(n3387), .ZN(n5618) );
  AOI22_X1 U22614 ( .A1(N3623), .A2(n25792), .B1(N3590), .B2(n23127), .ZN(
        n3387) );
  OAI21_X1 U22615 ( .B1(n19106), .B2(n10791), .A(n3388), .ZN(n5619) );
  AOI22_X1 U22616 ( .A1(N3622), .A2(n25775), .B1(N3589), .B2(n26146), .ZN(
        n3388) );
  OAI21_X1 U22617 ( .B1(n25130), .B2(n10796), .A(n3389), .ZN(n5620) );
  AOI22_X1 U22618 ( .A1(N3621), .A2(n25781), .B1(N3588), .B2(n24801), .ZN(
        n3389) );
  OAI21_X1 U22619 ( .B1(n22518), .B2(n11271), .A(n32120), .ZN(n5501) );
  AOI22_X1 U22620 ( .A1(N3036), .A2(n25550), .B1(N3003), .B2(n23133), .ZN(
        n32120) );
  OAI21_X1 U22621 ( .B1(n26558), .B2(n11279), .A(n32140), .ZN(n5503) );
  AOI22_X1 U22622 ( .A1(N3034), .A2(n25768), .B1(N3001), .B2(n24463), .ZN(
        n32140) );
  OAI21_X1 U22623 ( .B1(n25374), .B2(n11283), .A(n32150), .ZN(n5504) );
  AOI22_X1 U22624 ( .A1(N3033), .A2(n25772), .B1(N3000), .B2(n23129), .ZN(
        n32150) );
  OAI21_X1 U22625 ( .B1(n25372), .B2(n11287), .A(n32160), .ZN(n5505) );
  AOI22_X1 U22626 ( .A1(N3032), .A2(n25789), .B1(N2999), .B2(n21626), .ZN(
        n32160) );
  OAI21_X1 U22627 ( .B1(n25132), .B2(n11291), .A(n3217), .ZN(n5506) );
  AOI22_X1 U22628 ( .A1(N3031), .A2(n25793), .B1(N2998), .B2(n24796), .ZN(
        n3217) );
  OAI21_X1 U22629 ( .B1(n22513), .B2(n11295), .A(n3218), .ZN(n55070) );
  AOI22_X1 U22630 ( .A1(N3030), .A2(n25786), .B1(N2997), .B2(n26145), .ZN(
        n3218) );
  OAI21_X1 U22631 ( .B1(n23695), .B2(n11299), .A(n3219), .ZN(n55080) );
  AOI22_X1 U22632 ( .A1(N3029), .A2(n27239), .B1(N2996), .B2(n24808), .ZN(
        n3219) );
  OAI21_X1 U22633 ( .B1(n23700), .B2(n11303), .A(n3220), .ZN(n55090) );
  AOI22_X1 U22634 ( .A1(N3028), .A2(n25777), .B1(N2995), .B2(n24796), .ZN(
        n3220) );
  OAI21_X1 U22635 ( .B1(n23690), .B2(n11311), .A(n3222), .ZN(n55110) );
  AOI22_X1 U22636 ( .A1(N3026), .A2(n25769), .B1(N2993), .B2(n24452), .ZN(
        n3222) );
  OAI21_X1 U22637 ( .B1(n25141), .B2(n11315), .A(n3223), .ZN(n55120) );
  AOI22_X1 U22638 ( .A1(N3025), .A2(n25773), .B1(N2992), .B2(n20590), .ZN(
        n3223) );
  OAI21_X1 U22639 ( .B1(n19107), .B2(n11319), .A(n3224), .ZN(n55130) );
  AOI22_X1 U22640 ( .A1(N3024), .A2(n22928), .B1(N2991), .B2(n21643), .ZN(
        n3224) );
  OAI21_X1 U22641 ( .B1(n25134), .B2(n11323), .A(n3225), .ZN(n55140) );
  AOI22_X1 U22642 ( .A1(N3023), .A2(n22925), .B1(N2990), .B2(n26152), .ZN(
        n3225) );
  OAI21_X1 U22643 ( .B1(n25125), .B2(n11328), .A(n3226), .ZN(n55150) );
  AOI22_X1 U22644 ( .A1(N3022), .A2(n25831), .B1(N2989), .B2(n24463), .ZN(
        n3226) );
  OAI21_X1 U22645 ( .B1(n25157), .B2(n3014), .A(n44340), .ZN(n6303) );
  AOI22_X1 U22646 ( .A1(N7568), .A2(n25811), .B1(N7535), .B2(n24453), .ZN(
        n44340) );
  OAI21_X1 U22647 ( .B1(n25162), .B2(n7762), .A(n42700), .ZN(n61970) );
  AOI22_X1 U22648 ( .A1(N6964), .A2(n22912), .B1(N6931), .B2(n26156), .ZN(
        n42700) );
  OAI21_X1 U22649 ( .B1(n25147), .B2(n7795), .A(n42780), .ZN(n6205) );
  AOI22_X1 U22650 ( .A1(N6956), .A2(n27181), .B1(N6923), .B2(n24450), .ZN(
        n42780) );
  OAI21_X1 U22651 ( .B1(n25149), .B2(n8271), .A(n41060), .ZN(n6089) );
  AOI22_X1 U22652 ( .A1(N6361), .A2(n25800), .B1(N6328), .B2(n24454), .ZN(
        n41060) );
  OAI21_X1 U22653 ( .B1(n25124), .B2(n8279), .A(n41080), .ZN(n6091) );
  AOI22_X1 U22654 ( .A1(N6359), .A2(n22897), .B1(N6326), .B2(n23136), .ZN(
        n41080) );
  OAI21_X1 U22655 ( .B1(n25369), .B2(n8311), .A(n4116), .ZN(n60990) );
  AOI22_X1 U22656 ( .A1(N6351), .A2(n25810), .B1(N6318), .B2(n23297), .ZN(
        n4116) );
  OAI21_X1 U22657 ( .B1(n25139), .B2(n8602), .A(n40180), .ZN(n60330) );
  AOI22_X1 U22658 ( .A1(N6021), .A2(n25777), .B1(N5988), .B2(n24460), .ZN(
        n40180) );
  OAI21_X1 U22659 ( .B1(n25370), .B2(n8818), .A(n3945), .ZN(n59840) );
  AOI22_X1 U22660 ( .A1(N5765), .A2(n25851), .B1(N5732), .B2(n25991), .ZN(
        n3945) );
  OAI21_X1 U22661 ( .B1(n19044), .B2(n8854), .A(n3954), .ZN(n59930) );
  AOI22_X1 U22662 ( .A1(N5756), .A2(n22906), .B1(N5723), .B2(n23299), .ZN(
        n3954) );
  OAI21_X1 U22663 ( .B1(n25144), .B2(n9131), .A(n3860), .ZN(n59270) );
  AOI22_X1 U22664 ( .A1(N5426), .A2(n22924), .B1(N5393), .B2(n26154), .ZN(
        n3860) );
  OAI21_X1 U22665 ( .B1(n25129), .B2(n9170), .A(n3868), .ZN(n59350) );
  AOI22_X1 U22666 ( .A1(N5418), .A2(n27234), .B1(N5385), .B2(n24452), .ZN(
        n3868) );
  OAI21_X1 U22667 ( .B1(n25153), .B2(n9351), .A(n3784), .ZN(n5878) );
  AOI22_X1 U22668 ( .A1(N5180), .A2(n22899), .B1(N5147), .B2(n21653), .ZN(
        n3784) );
  OAI21_X1 U22669 ( .B1(n25156), .B2(n9391), .A(n37920), .ZN(n5886) );
  AOI22_X1 U22670 ( .A1(N5172), .A2(n22909), .B1(N5139), .B2(n20601), .ZN(
        n37920) );
  OAI21_X1 U22671 ( .B1(n25131), .B2(n9650), .A(n3697), .ZN(n58190) );
  AOI22_X1 U22672 ( .A1(N4831), .A2(n25766), .B1(N4798), .B2(n24460), .ZN(
        n3697) );
  OAI21_X1 U22673 ( .B1(n25126), .B2(n9660), .A(n3699), .ZN(n58210) );
  AOI22_X1 U22674 ( .A1(N4829), .A2(n22901), .B1(N4796), .B2(n23128), .ZN(
        n3699) );
  OAI21_X1 U22675 ( .B1(n25373), .B2(n9700), .A(n37070), .ZN(n5829) );
  AOI22_X1 U22676 ( .A1(N4821), .A2(n25776), .B1(N4788), .B2(n23285), .ZN(
        n37070) );
  OAI21_X1 U22677 ( .B1(n19045), .B2(n9878), .A(n36270), .ZN(n57720) );
  AOI22_X1 U22678 ( .A1(N4559), .A2(n24529), .B1(N4526), .B2(n25993), .ZN(
        n36270) );
  OAI21_X1 U22679 ( .B1(n25146), .B2(n9910), .A(n36350), .ZN(n5780) );
  AOI22_X1 U22680 ( .A1(N4551), .A2(n25816), .B1(N4518), .B2(n20598), .ZN(
        n36350) );
  OAI21_X1 U22681 ( .B1(n25374), .B2(n10184), .A(n35380), .ZN(n5714) );
  AOI22_X1 U22682 ( .A1(N4218), .A2(n25837), .B1(N4185), .B2(n25987), .ZN(
        n35380) );
  OAI21_X1 U22683 ( .B1(n19041), .B2(n10229), .A(n35470), .ZN(n57230) );
  AOI22_X1 U22684 ( .A1(N4209), .A2(n22918), .B1(N4176), .B2(n23287), .ZN(
        n35470) );
  OAI21_X1 U22685 ( .B1(n25135), .B2(n10747), .A(n33770), .ZN(n5608) );
  AOI22_X1 U22686 ( .A1(N3633), .A2(n22904), .B1(N3600), .B2(n21639), .ZN(
        n33770) );
  OAI21_X1 U22687 ( .B1(n25138), .B2(n10779), .A(n3385), .ZN(n5616) );
  AOI22_X1 U22688 ( .A1(N3625), .A2(n22922), .B1(N3592), .B2(n20880), .ZN(
        n3385) );
  OAI21_X1 U22689 ( .B1(n19042), .B2(n11275), .A(n32130), .ZN(n5502) );
  AOI22_X1 U22690 ( .A1(N3035), .A2(n24535), .B1(N3002), .B2(n25989), .ZN(
        n32130) );
  OAI21_X1 U22691 ( .B1(n25128), .B2(n11307), .A(n3221), .ZN(n55100) );
  AOI22_X1 U22692 ( .A1(N3027), .A2(n25782), .B1(N2994), .B2(n20604), .ZN(
        n3221) );
  AND3_X1 U22693 ( .A1(n27741), .A2(n25664), .A3(n457), .ZN(n5299) );
  NAND3_X1 U22694 ( .A1(n49110), .A2(n49120), .A3(n49130), .ZN(mul_outcome[57]) );
  AOI22_X1 U22695 ( .A1(n27060), .A2(n17821), .B1(n19230), .B2(n17809), .ZN(
        n49110) );
  AOI22_X1 U22696 ( .A1(n27063), .A2(n17845), .B1(n27076), .B2(n17833), .ZN(
        n49120) );
  AOI221_X1 U22697 ( .B1(n27087), .B2(n17797), .C1(n21356), .C2(n17785), .A(
        n27748), .ZN(n49130) );
  NAND3_X1 U22698 ( .A1(n47090), .A2(n47100), .A3(n4711), .ZN(mul_outcome[99])
         );
  AOI221_X1 U22699 ( .B1(n26620), .B2(n17581), .C1(n21970), .C2(n17569), .A(
        n27742), .ZN(n4711) );
  AOI22_X1 U22700 ( .A1(n26377), .A2(n17629), .B1(n26366), .B2(n17617), .ZN(
        n47090) );
  AOI22_X1 U22701 ( .A1(n25322), .A2(n17653), .B1(n25324), .B2(n17641), .ZN(
        n47100) );
  OR2_X1 U22702 ( .A1(n26967), .A2(n537), .ZN(sub_127_aco_carry[4]) );
  AND2_X1 U22703 ( .A1(n537), .A2(add_124_aco_B_3_), .ZN(n26969) );
  OAI21_X1 U22704 ( .B1(n21801), .B2(n7434), .A(n43770), .ZN(n62660) );
  AOI22_X1 U22705 ( .A1(N7407), .A2(n22316), .B1(N7374), .B2(n27208), .ZN(
        n43770) );
  OAI21_X1 U22706 ( .B1(n21825), .B2(n74390), .A(n43780), .ZN(n62670) );
  AOI22_X1 U22707 ( .A1(N7406), .A2(n22306), .B1(N7373), .B2(n25251), .ZN(
        n43780) );
  OAI21_X1 U22708 ( .B1(n21817), .B2(n74440), .A(n43790), .ZN(n62680) );
  AOI22_X1 U22709 ( .A1(N7405), .A2(n22296), .B1(N7372), .B2(n26737), .ZN(
        n43790) );
  OAI21_X1 U22710 ( .B1(n21805), .B2(n74490), .A(n43800), .ZN(n62690) );
  AOI22_X1 U22711 ( .A1(N7404), .A2(n22286), .B1(N7371), .B2(n25254), .ZN(
        n43800) );
  OAI21_X1 U22712 ( .B1(n21829), .B2(n74540), .A(n43810), .ZN(n62700) );
  AOI22_X1 U22713 ( .A1(N7403), .A2(n22321), .B1(N7370), .B2(n25267), .ZN(
        n43810) );
  OAI21_X1 U22714 ( .B1(n21821), .B2(n7459), .A(n43820), .ZN(n62710) );
  AOI22_X1 U22715 ( .A1(N7402), .A2(n22311), .B1(N7369), .B2(n22815), .ZN(
        n43820) );
  OAI21_X1 U22716 ( .B1(n26271), .B2(n7464), .A(n43830), .ZN(n62720) );
  AOI22_X1 U22717 ( .A1(N7401), .A2(n22301), .B1(N7368), .B2(n24187), .ZN(
        n43830) );
  OAI21_X1 U22718 ( .B1(n26296), .B2(n7469), .A(n43840), .ZN(n62730) );
  AOI22_X1 U22719 ( .A1(N7400), .A2(n22291), .B1(N7367), .B2(n24191), .ZN(
        n43840) );
  OAI21_X1 U22720 ( .B1(n26287), .B2(n74740), .A(n43850), .ZN(n62740) );
  AOI22_X1 U22721 ( .A1(N7399), .A2(n24340), .B1(N7366), .B2(n22815), .ZN(
        n43850) );
  OAI21_X1 U22722 ( .B1(n26796), .B2(n74790), .A(n43860), .ZN(n62750) );
  AOI22_X1 U22723 ( .A1(N7398), .A2(n24345), .B1(N7365), .B2(n24471), .ZN(
        n43860) );
  OAI21_X1 U22724 ( .B1(n26785), .B2(n74840), .A(n43870), .ZN(n62760) );
  AOI22_X1 U22725 ( .A1(N7397), .A2(n24352), .B1(N7364), .B2(n21282), .ZN(
        n43870) );
  OAI21_X1 U22726 ( .B1(n26789), .B2(n74890), .A(n43880), .ZN(n62770) );
  AOI22_X1 U22727 ( .A1(N7396), .A2(n23333), .B1(N7363), .B2(n25621), .ZN(
        n43880) );
  OAI21_X1 U22728 ( .B1(n21799), .B2(n7494), .A(n43890), .ZN(n62780) );
  AOI22_X1 U22729 ( .A1(N7395), .A2(n26207), .B1(N7362), .B2(n21287), .ZN(
        n43890) );
  OAI21_X1 U22730 ( .B1(n21823), .B2(n7499), .A(n43900), .ZN(n62790) );
  AOI22_X1 U22731 ( .A1(N7394), .A2(n24348), .B1(N7361), .B2(n24783), .ZN(
        n43900) );
  OAI21_X1 U22732 ( .B1(n21815), .B2(n7503), .A(n43910), .ZN(n62800) );
  AOI22_X1 U22733 ( .A1(N7393), .A2(n26199), .B1(N7360), .B2(n21283), .ZN(
        n43910) );
  OAI21_X1 U22734 ( .B1(n21803), .B2(n78730), .A(n42200), .ZN(n61610) );
  AOI22_X1 U22735 ( .A1(N6796), .A2(n22304), .B1(N6763), .B2(n25254), .ZN(
        n42200) );
  OAI21_X1 U22736 ( .B1(n21827), .B2(n78780), .A(n42210), .ZN(n61620) );
  AOI22_X1 U22737 ( .A1(N6795), .A2(n22294), .B1(N6762), .B2(n21303), .ZN(
        n42210) );
  OAI21_X1 U22738 ( .B1(n21819), .B2(n7883), .A(n42220), .ZN(n61630) );
  AOI22_X1 U22739 ( .A1(N6794), .A2(n26195), .B1(N6761), .B2(n21291), .ZN(
        n42220) );
  OAI21_X1 U22740 ( .B1(n19264), .B2(n7888), .A(n42230), .ZN(n61640) );
  AOI22_X1 U22741 ( .A1(N6793), .A2(n22314), .B1(N6760), .B2(n20582), .ZN(
        n42230) );
  OAI21_X1 U22742 ( .B1(n26783), .B2(n7893), .A(n42240), .ZN(n6165) );
  AOI22_X1 U22743 ( .A1(N6792), .A2(n22308), .B1(N6759), .B2(n26747), .ZN(
        n42240) );
  OAI21_X1 U22744 ( .B1(n19265), .B2(n78980), .A(n42250), .ZN(n6166) );
  AOI22_X1 U22745 ( .A1(N6791), .A2(n22299), .B1(N6758), .B2(n21426), .ZN(
        n42250) );
  OAI21_X1 U22746 ( .B1(n26795), .B2(n79030), .A(n42260), .ZN(n6167) );
  AOI22_X1 U22747 ( .A1(N6790), .A2(n22284), .B1(N6757), .B2(n25882), .ZN(
        n42260) );
  OAI21_X1 U22748 ( .B1(n26784), .B2(n79080), .A(n42270), .ZN(n6168) );
  AOI22_X1 U22749 ( .A1(N6789), .A2(n22319), .B1(N6756), .B2(n21282), .ZN(
        n42270) );
  OAI21_X1 U22750 ( .B1(n26788), .B2(n79130), .A(n4228), .ZN(n6169) );
  AOI22_X1 U22751 ( .A1(N6788), .A2(n23340), .B1(N6755), .B2(n22812), .ZN(
        n4228) );
  OAI21_X1 U22752 ( .B1(n26276), .B2(n7918), .A(n4229), .ZN(n6170) );
  AOI22_X1 U22753 ( .A1(N6787), .A2(n23337), .B1(N6754), .B2(n25256), .ZN(
        n4229) );
  OAI21_X1 U22754 ( .B1(n26302), .B2(n7923), .A(n4230), .ZN(n6171) );
  AOI22_X1 U22755 ( .A1(N6786), .A2(n22288), .B1(N6753), .B2(n26736), .ZN(
        n4230) );
  OAI21_X1 U22756 ( .B1(n26293), .B2(n7928), .A(n4231), .ZN(n6172) );
  AOI22_X1 U22757 ( .A1(N6785), .A2(n23343), .B1(N6752), .B2(n22816), .ZN(
        n4231) );
  OAI21_X1 U22758 ( .B1(n26278), .B2(n7933), .A(n4232), .ZN(n6173) );
  AOI22_X1 U22759 ( .A1(N6784), .A2(n26203), .B1(N6751), .B2(n25880), .ZN(
        n4232) );
  OAI21_X1 U22760 ( .B1(n26304), .B2(n7938), .A(n4233), .ZN(n6174) );
  AOI22_X1 U22761 ( .A1(N6783), .A2(n24354), .B1(N6750), .B2(n23070), .ZN(
        n4233) );
  OAI21_X1 U22762 ( .B1(n26295), .B2(n79420), .A(n4234), .ZN(n6175) );
  AOI22_X1 U22763 ( .A1(N6782), .A2(n24361), .B1(N6749), .B2(n25882), .ZN(
        n4234) );
  OAI21_X1 U22764 ( .B1(n26796), .B2(n8407), .A(n40590), .ZN(n6056) );
  AOI22_X1 U22765 ( .A1(N6196), .A2(n26462), .B1(N6163), .B2(n21299), .ZN(
        n40590) );
  OAI21_X1 U22766 ( .B1(n26785), .B2(n8412), .A(n4060), .ZN(n6057) );
  AOI22_X1 U22767 ( .A1(N6195), .A2(n24358), .B1(N6162), .B2(n25616), .ZN(
        n4060) );
  OAI21_X1 U22768 ( .B1(n26789), .B2(n8417), .A(n4061), .ZN(n6058) );
  AOI22_X1 U22769 ( .A1(N6194), .A2(n24342), .B1(N6161), .B2(n26729), .ZN(
        n4061) );
  OAI21_X1 U22770 ( .B1(n24285), .B2(n8422), .A(n4062), .ZN(n6059) );
  AOI22_X1 U22771 ( .A1(N6193), .A2(n26468), .B1(N6160), .B2(n24780), .ZN(
        n4062) );
  OAI21_X1 U22772 ( .B1(n24267), .B2(n8427), .A(n4063), .ZN(n60600) );
  AOI22_X1 U22773 ( .A1(N6192), .A2(n26465), .B1(N6159), .B2(n20584), .ZN(
        n4063) );
  OAI21_X1 U22774 ( .B1(n24273), .B2(n8432), .A(n4064), .ZN(n60610) );
  AOI22_X1 U22775 ( .A1(N6191), .A2(n26456), .B1(N6158), .B2(n24783), .ZN(
        n4064) );
  OAI21_X1 U22776 ( .B1(n26275), .B2(n8437), .A(n4065), .ZN(n60620) );
  AOI22_X1 U22777 ( .A1(N6190), .A2(n26474), .B1(N6157), .B2(n17120), .ZN(
        n4065) );
  OAI21_X1 U22778 ( .B1(n26301), .B2(n8442), .A(n4066), .ZN(n60630) );
  AOI22_X1 U22779 ( .A1(N6189), .A2(n26472), .B1(N6156), .B2(n25622), .ZN(
        n4066) );
  OAI21_X1 U22780 ( .B1(n26292), .B2(n8447), .A(n4067), .ZN(n60640) );
  AOI22_X1 U22781 ( .A1(N6188), .A2(n24351), .B1(N6155), .B2(n21010), .ZN(
        n4067) );
  OAI21_X1 U22782 ( .B1(n26277), .B2(n8452), .A(n4068), .ZN(n60650) );
  AOI22_X1 U22783 ( .A1(N6187), .A2(n264601), .B1(N6154), .B2(n25265), .ZN(
        n4068) );
  OAI21_X1 U22784 ( .B1(n26303), .B2(n8457), .A(n4069), .ZN(n60660) );
  AOI22_X1 U22785 ( .A1(N6186), .A2(n26478), .B1(N6153), .B2(n25618), .ZN(
        n4069) );
  OAI21_X1 U22786 ( .B1(n26294), .B2(n8462), .A(n4070), .ZN(n60670) );
  AOI22_X1 U22787 ( .A1(N6185), .A2(n24346), .B1(N6152), .B2(n24188), .ZN(
        n4070) );
  OAI21_X1 U22788 ( .B1(n26794), .B2(n8467), .A(n4071), .ZN(n60680) );
  AOI22_X1 U22789 ( .A1(N6184), .A2(n26198), .B1(N6151), .B2(n20580), .ZN(
        n4071) );
  OAI21_X1 U22790 ( .B1(n26783), .B2(n8472), .A(n4072), .ZN(n60690) );
  AOI22_X1 U22791 ( .A1(N6183), .A2(n23334), .B1(N6150), .B2(n25258), .ZN(
        n4072) );
  OAI21_X1 U22792 ( .B1(n26787), .B2(n8476), .A(n4073), .ZN(n60700) );
  AOI22_X1 U22793 ( .A1(N6182), .A2(n24339), .B1(N6149), .B2(n19303), .ZN(
        n4073) );
  OAI21_X1 U22794 ( .B1(n26274), .B2(n8941), .A(n3898), .ZN(n5951) );
  AOI22_X1 U22795 ( .A1(N5600), .A2(n26194), .B1(N5567), .B2(n26743), .ZN(
        n3898) );
  OAI21_X1 U22796 ( .B1(n26300), .B2(n8946), .A(n3899), .ZN(n5952) );
  AOI22_X1 U22797 ( .A1(N5599), .A2(n26206), .B1(N5566), .B2(n20583), .ZN(
        n3899) );
  OAI21_X1 U22798 ( .B1(n26291), .B2(n8951), .A(n3900), .ZN(n5953) );
  AOI22_X1 U22799 ( .A1(N5598), .A2(n24349), .B1(N5565), .B2(n27207), .ZN(
        n3900) );
  OAI21_X1 U22800 ( .B1(n21801), .B2(n8956), .A(n3901), .ZN(n5954) );
  AOI22_X1 U22801 ( .A1(N5597), .A2(n26464), .B1(N5564), .B2(n19213), .ZN(
        n3901) );
  OAI21_X1 U22802 ( .B1(n21825), .B2(n8961), .A(n3902), .ZN(n5955) );
  AOI22_X1 U22803 ( .A1(N5596), .A2(n26458), .B1(N5563), .B2(n24778), .ZN(
        n3902) );
  OAI21_X1 U22804 ( .B1(n21817), .B2(n8966), .A(n3903), .ZN(n5956) );
  AOI22_X1 U22805 ( .A1(N5595), .A2(n26476), .B1(N5562), .B2(n25255), .ZN(
        n3903) );
  OAI21_X1 U22806 ( .B1(n21806), .B2(n8971), .A(n3904), .ZN(n5957) );
  AOI22_X1 U22807 ( .A1(N5594), .A2(n264701), .B1(N5561), .B2(n22813), .ZN(
        n3904) );
  OAI21_X1 U22808 ( .B1(n21830), .B2(n8976), .A(n3905), .ZN(n5958) );
  AOI22_X1 U22809 ( .A1(N5593), .A2(n26467), .B1(N5560), .B2(n19214), .ZN(
        n3905) );
  OAI21_X1 U22810 ( .B1(n21822), .B2(n8981), .A(n3906), .ZN(n5959) );
  AOI22_X1 U22811 ( .A1(N5592), .A2(n26461), .B1(N5559), .B2(n26729), .ZN(
        n3906) );
  OAI21_X1 U22812 ( .B1(n24285), .B2(n8986), .A(n3907), .ZN(n5960) );
  AOI22_X1 U22813 ( .A1(N5591), .A2(n26479), .B1(N5558), .B2(n25611), .ZN(
        n3907) );
  OAI21_X1 U22814 ( .B1(n24267), .B2(n8991), .A(n3908), .ZN(n5961) );
  AOI22_X1 U22815 ( .A1(N5590), .A2(n26473), .B1(N5557), .B2(n20584), .ZN(
        n3908) );
  OAI21_X1 U22816 ( .B1(n24273), .B2(n8996), .A(n3909), .ZN(n5962) );
  AOI22_X1 U22817 ( .A1(N5589), .A2(n26196), .B1(N5556), .B2(n20579), .ZN(
        n3909) );
  OAI21_X1 U22818 ( .B1(n24286), .B2(n9001), .A(n3910), .ZN(n5963) );
  AOI22_X1 U22819 ( .A1(N5588), .A2(n26192), .B1(N5555), .B2(n25614), .ZN(
        n3910) );
  OAI21_X1 U22820 ( .B1(n24268), .B2(n9006), .A(n3911), .ZN(n5964) );
  AOI22_X1 U22821 ( .A1(N5587), .A2(n26844), .B1(N5554), .B2(n19217), .ZN(
        n3911) );
  OAI21_X1 U22822 ( .B1(n24274), .B2(n9010), .A(n3912), .ZN(n5965) );
  AOI22_X1 U22823 ( .A1(N5586), .A2(n26848), .B1(N5553), .B2(n21427), .ZN(
        n3912) );
  OAI21_X1 U22824 ( .B1(n21799), .B2(n9500), .A(n3738), .ZN(n58460) );
  AOI22_X1 U22825 ( .A1(N5008), .A2(n26204), .B1(N4975), .B2(n24187), .ZN(
        n3738) );
  OAI21_X1 U22826 ( .B1(n21823), .B2(n9504), .A(n3739), .ZN(n58470) );
  AOI22_X1 U22827 ( .A1(N5007), .A2(n26200), .B1(N4974), .B2(n23069), .ZN(
        n3739) );
  OAI21_X1 U22828 ( .B1(n21815), .B2(n9508), .A(n3740), .ZN(n58480) );
  AOI22_X1 U22829 ( .A1(N5006), .A2(n26849), .B1(N4973), .B2(n21010), .ZN(
        n3740) );
  OAI21_X1 U22830 ( .B1(n21804), .B2(n9512), .A(n3741), .ZN(n58490) );
  AOI22_X1 U22831 ( .A1(N5005), .A2(n26853), .B1(N4972), .B2(n25622), .ZN(
        n3741) );
  OAI21_X1 U22832 ( .B1(n21828), .B2(n9516), .A(n3742), .ZN(n58500) );
  AOI22_X1 U22833 ( .A1(N5004), .A2(n22317), .B1(N4971), .B2(n25256), .ZN(
        n3742) );
  OAI21_X1 U22834 ( .B1(n21820), .B2(n9520), .A(n3743), .ZN(n58510) );
  AOI22_X1 U22835 ( .A1(N5003), .A2(n22307), .B1(N4970), .B2(n25267), .ZN(
        n3743) );
  OAI21_X1 U22836 ( .B1(n26274), .B2(n9524), .A(n3744), .ZN(n58520) );
  AOI22_X1 U22837 ( .A1(N5002), .A2(n22297), .B1(N4969), .B2(n25616), .ZN(
        n3744) );
  OAI21_X1 U22838 ( .B1(n26300), .B2(n9528), .A(n3745), .ZN(n58530) );
  AOI22_X1 U22839 ( .A1(N5001), .A2(n22287), .B1(N4968), .B2(n23070), .ZN(
        n3745) );
  OAI21_X1 U22840 ( .B1(n26291), .B2(n9532), .A(n3746), .ZN(n58540) );
  AOI22_X1 U22841 ( .A1(N5000), .A2(n22322), .B1(N4967), .B2(n24188), .ZN(
        n3746) );
  OAI21_X1 U22842 ( .B1(n26273), .B2(n9536), .A(n3747), .ZN(n58550) );
  AOI22_X1 U22843 ( .A1(N4999), .A2(n22312), .B1(N4966), .B2(n19303), .ZN(
        n3747) );
  OAI21_X1 U22844 ( .B1(n26299), .B2(n9540), .A(n3748), .ZN(n58560) );
  AOI22_X1 U22845 ( .A1(N4998), .A2(n22302), .B1(N4965), .B2(n24191), .ZN(
        n3748) );
  OAI21_X1 U22846 ( .B1(n26290), .B2(n9544), .A(n3749), .ZN(n58570) );
  AOI22_X1 U22847 ( .A1(N4997), .A2(n22292), .B1(N4964), .B2(n25251), .ZN(
        n3749) );
  OAI21_X1 U22848 ( .B1(n26276), .B2(n9548), .A(n3750), .ZN(n58580) );
  AOI22_X1 U22849 ( .A1(N4996), .A2(n26842), .B1(N4963), .B2(n22812), .ZN(
        n3750) );
  OAI21_X1 U22850 ( .B1(n26302), .B2(n9552), .A(n3751), .ZN(n58590) );
  AOI22_X1 U22851 ( .A1(N4995), .A2(n26846), .B1(N4962), .B2(n25612), .ZN(
        n3751) );
  OAI21_X1 U22852 ( .B1(n26293), .B2(n9557), .A(n3752), .ZN(n58600) );
  AOI22_X1 U22853 ( .A1(N4994), .A2(n26199), .B1(N4961), .B2(n21300), .ZN(
        n3752) );
  OAI21_X1 U22854 ( .B1(n26278), .B2(n10009), .A(n3579), .ZN(n5741) );
  AOI22_X1 U22855 ( .A1(N4389), .A2(n26202), .B1(N4356), .B2(n24776), .ZN(
        n3579) );
  OAI21_X1 U22856 ( .B1(n26304), .B2(n10014), .A(n3580), .ZN(n5742) );
  AOI22_X1 U22857 ( .A1(N4388), .A2(n24355), .B1(N4355), .B2(n25615), .ZN(
        n3580) );
  OAI21_X1 U22858 ( .B1(n26295), .B2(n10019), .A(n3581), .ZN(n5743) );
  AOI22_X1 U22859 ( .A1(N4387), .A2(n19258), .B1(N4354), .B2(n19218), .ZN(
        n3581) );
  OAI21_X1 U22860 ( .B1(n24286), .B2(n10024), .A(n3582), .ZN(n5744) );
  AOI22_X1 U22861 ( .A1(N4386), .A2(n24343), .B1(N4353), .B2(n26746), .ZN(
        n3582) );
  OAI21_X1 U22862 ( .B1(n24268), .B2(n10029), .A(n3583), .ZN(n5745) );
  AOI22_X1 U22863 ( .A1(N4385), .A2(n22303), .B1(N4352), .B2(n26738), .ZN(
        n3583) );
  OAI21_X1 U22864 ( .B1(n24274), .B2(n10034), .A(n3584), .ZN(n5746) );
  AOI22_X1 U22865 ( .A1(N4384), .A2(n22293), .B1(N4351), .B2(n21290), .ZN(
        n3584) );
  OAI21_X1 U22866 ( .B1(n24289), .B2(n10039), .A(n3585), .ZN(n5747) );
  AOI22_X1 U22867 ( .A1(N4383), .A2(n24357), .B1(N4350), .B2(n25881), .ZN(
        n3585) );
  OAI21_X1 U22868 ( .B1(n24271), .B2(n10044), .A(n3586), .ZN(n5748) );
  AOI22_X1 U22869 ( .A1(N4382), .A2(n22313), .B1(N4349), .B2(n25881), .ZN(
        n3586) );
  OAI21_X1 U22870 ( .B1(n24277), .B2(n10049), .A(n3587), .ZN(n5749) );
  AOI22_X1 U22871 ( .A1(N4381), .A2(n22309), .B1(N4348), .B2(n26745), .ZN(
        n3587) );
  OAI21_X1 U22872 ( .B1(n26275), .B2(n10054), .A(n35880), .ZN(n5750) );
  AOI22_X1 U22873 ( .A1(N4380), .A2(n22298), .B1(N4347), .B2(n21424), .ZN(
        n35880) );
  OAI21_X1 U22874 ( .B1(n26301), .B2(n10059), .A(n35890), .ZN(n5751) );
  AOI22_X1 U22875 ( .A1(N4379), .A2(n22283), .B1(N4346), .B2(n21011), .ZN(
        n35890) );
  OAI21_X1 U22876 ( .B1(n26292), .B2(n10064), .A(n35900), .ZN(n5752) );
  AOI22_X1 U22877 ( .A1(N4378), .A2(n22318), .B1(N4345), .B2(n25268), .ZN(
        n35900) );
  OAI21_X1 U22878 ( .B1(n26277), .B2(n10069), .A(n35910), .ZN(n5753) );
  AOI22_X1 U22879 ( .A1(N4377), .A2(n19260), .B1(N4344), .B2(n25258), .ZN(
        n35910) );
  OAI21_X1 U22880 ( .B1(n26303), .B2(n10074), .A(n35920), .ZN(n57540) );
  AOI22_X1 U22881 ( .A1(N4376), .A2(n19259), .B1(N4343), .B2(n20578), .ZN(
        n35920) );
  OAI21_X1 U22882 ( .B1(n26294), .B2(n10078), .A(n35930), .ZN(n57550) );
  AOI22_X1 U22883 ( .A1(N4375), .A2(n22289), .B1(N4342), .B2(n25612), .ZN(
        n35930) );
  OAI21_X1 U22884 ( .B1(n26273), .B2(n10569), .A(n3419), .ZN(n5636) );
  AOI22_X1 U22885 ( .A1(N3803), .A2(n23336), .B1(N3770), .B2(n25614), .ZN(
        n3419) );
  OAI21_X1 U22886 ( .B1(n26299), .B2(n10574), .A(n34200), .ZN(n5637) );
  AOI22_X1 U22887 ( .A1(N3802), .A2(n26854), .B1(N3769), .B2(n25621), .ZN(
        n34200) );
  OAI21_X1 U22888 ( .B1(n26290), .B2(n10579), .A(n34210), .ZN(n5638) );
  AOI22_X1 U22889 ( .A1(N3801), .A2(n19261), .B1(N3768), .B2(n21286), .ZN(
        n34210) );
  OAI21_X1 U22890 ( .B1(n23404), .B2(n10584), .A(n34220), .ZN(n5639) );
  AOI22_X1 U22891 ( .A1(N3800), .A2(n23339), .B1(N3767), .B2(n24780), .ZN(
        n34220) );
  OAI21_X1 U22892 ( .B1(n20506), .B2(n10589), .A(n34230), .ZN(n5640) );
  AOI22_X1 U22893 ( .A1(N3799), .A2(n26463), .B1(N3766), .B2(n22817), .ZN(
        n34230) );
  OAI21_X1 U22894 ( .B1(n23418), .B2(n10594), .A(n34240), .ZN(n5641) );
  AOI22_X1 U22895 ( .A1(N3798), .A2(n24360), .B1(N3765), .B2(n21426), .ZN(
        n34240) );
  OAI21_X1 U22896 ( .B1(n21802), .B2(n10599), .A(n34250), .ZN(n56420) );
  AOI22_X1 U22897 ( .A1(N3797), .A2(n23342), .B1(N3764), .B2(n24190), .ZN(
        n34250) );
  OAI21_X1 U22898 ( .B1(n21826), .B2(n10604), .A(n34260), .ZN(n56430) );
  AOI22_X1 U22899 ( .A1(N3796), .A2(n26469), .B1(N3763), .B2(n22818), .ZN(
        n34260) );
  OAI21_X1 U22900 ( .B1(n21818), .B2(n10609), .A(n34270), .ZN(n56440) );
  AOI22_X1 U22901 ( .A1(N3795), .A2(n26466), .B1(N3762), .B2(n21302), .ZN(
        n34270) );
  OAI21_X1 U22902 ( .B1(n21805), .B2(n10614), .A(n34280), .ZN(n56450) );
  AOI22_X1 U22903 ( .A1(N3794), .A2(n26457), .B1(N3761), .B2(n25618), .ZN(
        n34280) );
  OAI21_X1 U22904 ( .B1(n21829), .B2(n10619), .A(n34290), .ZN(n56460) );
  AOI22_X1 U22905 ( .A1(N3793), .A2(n26475), .B1(N3760), .B2(n25265), .ZN(
        n34290) );
  OAI21_X1 U22906 ( .B1(n21821), .B2(n10624), .A(n34300), .ZN(n56470) );
  AOI22_X1 U22907 ( .A1(N3792), .A2(n26471), .B1(N3759), .B2(n26744), .ZN(
        n34300) );
  OAI21_X1 U22908 ( .B1(n24289), .B2(n10629), .A(n34310), .ZN(n56480) );
  AOI22_X1 U22909 ( .A1(N3791), .A2(n26851), .B1(N3758), .B2(n24190), .ZN(
        n34310) );
  OAI21_X1 U22910 ( .B1(n24271), .B2(n10634), .A(n34320), .ZN(n56490) );
  AOI22_X1 U22911 ( .A1(N3790), .A2(n26459), .B1(N3757), .B2(n23069), .ZN(
        n34320) );
  OAI21_X1 U22912 ( .B1(n24277), .B2(n10638), .A(n34330), .ZN(n56500) );
  AOI22_X1 U22913 ( .A1(N3789), .A2(n26477), .B1(N3756), .B2(n24470), .ZN(
        n34330) );
  OAI21_X1 U22914 ( .B1(n24288), .B2(n11124), .A(n32620), .ZN(n5531) );
  AOI22_X1 U22915 ( .A1(N3210), .A2(n24358), .B1(N3177), .B2(n19306), .ZN(
        n32620) );
  OAI21_X1 U22916 ( .B1(n24270), .B2(n11128), .A(n32630), .ZN(n5532) );
  AOI22_X1 U22917 ( .A1(N3209), .A2(n24343), .B1(N3176), .B2(n25259), .ZN(
        n32630) );
  OAI21_X1 U22918 ( .B1(n24276), .B2(n11132), .A(n32640), .ZN(n5533) );
  AOI22_X1 U22919 ( .A1(N3208), .A2(n26203), .B1(N3175), .B2(n24778), .ZN(
        n32640) );
  OAI21_X1 U22920 ( .B1(n21800), .B2(n11136), .A(n32650), .ZN(n5534) );
  AOI22_X1 U22921 ( .A1(N3207), .A2(n24355), .B1(N3174), .B2(n22800), .ZN(
        n32650) );
  OAI21_X1 U22922 ( .B1(n21824), .B2(n11140), .A(n32660), .ZN(n5535) );
  AOI22_X1 U22923 ( .A1(N3206), .A2(n26195), .B1(N3173), .B2(n22799), .ZN(
        n32660) );
  OAI21_X1 U22924 ( .B1(n21816), .B2(n11144), .A(n32670), .ZN(n5536) );
  AOI22_X1 U22925 ( .A1(N3205), .A2(n26207), .B1(N3172), .B2(n20581), .ZN(
        n32670) );
  OAI21_X1 U22926 ( .B1(n21803), .B2(n11148), .A(n3268), .ZN(n5537) );
  AOI22_X1 U22927 ( .A1(N3204), .A2(n24349), .B1(N3171), .B2(n25611), .ZN(
        n3268) );
  OAI21_X1 U22928 ( .B1(n21827), .B2(n11152), .A(n3269), .ZN(n5538) );
  AOI22_X1 U22929 ( .A1(N3203), .A2(n26464), .B1(N3170), .B2(n19217), .ZN(
        n3269) );
  OAI21_X1 U22930 ( .B1(n21819), .B2(n11156), .A(n3270), .ZN(n5539) );
  AOI22_X1 U22931 ( .A1(N3202), .A2(n26458), .B1(N3169), .B2(n25615), .ZN(
        n3270) );
  OAI21_X1 U22932 ( .B1(n23404), .B2(n11160), .A(n3271), .ZN(n5540) );
  AOI22_X1 U22933 ( .A1(N3201), .A2(n26476), .B1(N3168), .B2(n19218), .ZN(
        n3271) );
  OAI21_X1 U22934 ( .B1(n20505), .B2(n11164), .A(n3272), .ZN(n5541) );
  AOI22_X1 U22935 ( .A1(N3200), .A2(n264701), .B1(N3167), .B2(n19213), .ZN(
        n3272) );
  OAI21_X1 U22936 ( .B1(n23418), .B2(n11168), .A(n3273), .ZN(n5542) );
  AOI22_X1 U22937 ( .A1(N3199), .A2(n26467), .B1(N3166), .B2(n24776), .ZN(
        n3273) );
  OAI21_X1 U22938 ( .B1(n23403), .B2(n11172), .A(n3274), .ZN(n5543) );
  AOI22_X1 U22939 ( .A1(N3198), .A2(n26461), .B1(N3165), .B2(n25880), .ZN(
        n3274) );
  OAI21_X1 U22940 ( .B1(n23424), .B2(n11176), .A(n3275), .ZN(n5544) );
  AOI22_X1 U22941 ( .A1(N3197), .A2(n26479), .B1(N3164), .B2(n19214), .ZN(
        n3275) );
  OAI21_X1 U22942 ( .B1(n23417), .B2(n11181), .A(n3276), .ZN(n5545) );
  AOI22_X1 U22943 ( .A1(N3196), .A2(n26473), .B1(N3163), .B2(n24471), .ZN(
        n3276) );
  NAND3_X1 U22944 ( .A1(n4783), .A2(n4784), .A3(n4785), .ZN(mul_outcome[83])
         );
  AOI22_X1 U22945 ( .A1(n25756), .A2(n17715), .B1(n26592), .B2(n17667), .ZN(
        n4783) );
  AOI22_X1 U22946 ( .A1(n27105), .A2(n17739), .B1(n25748), .B2(n17727), .ZN(
        n4784) );
  AOI221_X1 U22947 ( .B1(n21832), .B2(n17679), .C1(n26623), .C2(n17655), .A(
        n277601), .ZN(n4785) );
  NAND2_X1 U22948 ( .A1(n50110), .A2(n50120), .ZN(mul_outcome[36]) );
  AOI221_X1 U22949 ( .B1(n26105), .B2(n17869), .C1(n26057), .C2(n17857), .A(
        n50140), .ZN(n50110) );
  AOI221_X1 U22950 ( .B1(n26107), .B2(n17893), .C1(n261001), .C2(n17881), .A(
        n50130), .ZN(n50120) );
  OAI22_X1 U22951 ( .A1(n2069), .A2(n19206), .B1(n2048), .B2(n19196), .ZN(
        n50140) );
  NAND3_X1 U22952 ( .A1(n5300), .A2(n5301), .A3(n5302), .ZN(mul_outcome[125])
         );
  AOI221_X1 U22953 ( .B1(n21968), .B2(n17475), .C1(n26757), .C2(n17463), .A(
        n27774), .ZN(n5302) );
  AOI22_X1 U22954 ( .A1(n27021), .A2(n17547), .B1(n24747), .B2(n17535), .ZN(
        n5301) );
  AOI22_X1 U22955 ( .A1(n27007), .A2(n17523), .B1(n260601), .B2(n17511), .ZN(
        n5300) );
  OAI21_X1 U22956 ( .B1(n20723), .B2(n2923), .A(n4452), .ZN(n6312) );
  AOI22_X1 U22957 ( .A1(N7653), .A2(n25180), .B1(N7620), .B2(n26249), .ZN(
        n4452) );
  OAI21_X1 U22958 ( .B1(n25336), .B2(n2927), .A(n4453), .ZN(n6313) );
  AOI22_X1 U22959 ( .A1(N7652), .A2(n25168), .B1(N7619), .B2(n26245), .ZN(
        n4453) );
  OAI21_X1 U22960 ( .B1(n24954), .B2(n2935), .A(n4455), .ZN(n6315) );
  AOI22_X1 U22961 ( .A1(N7650), .A2(n25170), .B1(N7617), .B2(n26257), .ZN(
        n4455) );
  OAI21_X1 U22962 ( .B1(n20725), .B2(n29430), .A(n4457), .ZN(n63170) );
  AOI22_X1 U22963 ( .A1(N7648), .A2(n25182), .B1(N7615), .B2(n21776), .ZN(
        n4457) );
  OAI21_X1 U22964 ( .B1(n26699), .B2(n29470), .A(n4458), .ZN(n63180) );
  AOI22_X1 U22965 ( .A1(N7647), .A2(n22934), .B1(N7614), .B2(n26258), .ZN(
        n4458) );
  OAI21_X1 U22966 ( .B1(n25334), .B2(n29510), .A(n4459), .ZN(n63190) );
  AOI22_X1 U22967 ( .A1(N7646), .A2(n25558), .B1(N7613), .B2(n26261), .ZN(
        n4459) );
  OAI21_X1 U22968 ( .B1(n24951), .B2(n29550), .A(n4460), .ZN(n63200) );
  AOI22_X1 U22969 ( .A1(N7645), .A2(n21207), .B1(N7612), .B2(n26253), .ZN(
        n4460) );
  OAI21_X1 U22970 ( .B1(n25531), .B2(n2963), .A(n4462), .ZN(n63220) );
  AOI22_X1 U22971 ( .A1(N7643), .A2(n24550), .B1(N7610), .B2(n24297), .ZN(
        n4462) );
  OAI21_X1 U22972 ( .B1(n26698), .B2(n2967), .A(n4463), .ZN(n63230) );
  AOI22_X1 U22973 ( .A1(N7642), .A2(n24551), .B1(N7609), .B2(n26802), .ZN(
        n4463) );
  OAI21_X1 U22974 ( .B1(n25120), .B2(n2971), .A(n44640), .ZN(n63240) );
  AOI22_X1 U22975 ( .A1(N7641), .A2(n24536), .B1(N7608), .B2(n26249), .ZN(
        n44640) );
  OAI21_X1 U22976 ( .B1(n26697), .B2(n2976), .A(n44650), .ZN(n63250) );
  AOI22_X1 U22977 ( .A1(N7640), .A2(n24559), .B1(N7607), .B2(n26248), .ZN(
        n44650) );
  OAI21_X1 U22978 ( .B1(n24947), .B2(n7671), .A(n4286), .ZN(n6206) );
  AOI22_X1 U22979 ( .A1(N7062), .A2(n21202), .B1(N7029), .B2(n26250), .ZN(
        n4286) );
  OAI21_X1 U22980 ( .B1(n25532), .B2(n7675), .A(n4287), .ZN(n6207) );
  AOI22_X1 U22981 ( .A1(N7061), .A2(n24551), .B1(N7028), .B2(n26252), .ZN(
        n4287) );
  OAI21_X1 U22982 ( .B1(n19297), .B2(n7683), .A(n4289), .ZN(n6209) );
  AOI22_X1 U22983 ( .A1(N7059), .A2(n24558), .B1(N7026), .B2(n26259), .ZN(
        n4289) );
  OAI21_X1 U22984 ( .B1(n24949), .B2(n7691), .A(n4291), .ZN(n6211) );
  AOI22_X1 U22985 ( .A1(N7057), .A2(n24539), .B1(N7024), .B2(n24307), .ZN(
        n4291) );
  OAI21_X1 U22986 ( .B1(n22776), .B2(n7695), .A(n4292), .ZN(n6212) );
  AOI22_X1 U22987 ( .A1(N7056), .A2(n25562), .B1(N7023), .B2(n21787), .ZN(
        n4292) );
  OAI21_X1 U22988 ( .B1(n19088), .B2(n76990), .A(n4293), .ZN(n6213) );
  AOI22_X1 U22989 ( .A1(N7055), .A2(n21225), .B1(N7022), .B2(n26254), .ZN(
        n4293) );
  OAI21_X1 U22990 ( .B1(n20729), .B2(n77030), .A(n4294), .ZN(n6214) );
  AOI22_X1 U22991 ( .A1(N7054), .A2(n21216), .B1(N7021), .B2(n24306), .ZN(
        n4294) );
  OAI21_X1 U22992 ( .B1(n19087), .B2(n77110), .A(n42960), .ZN(n6216) );
  AOI22_X1 U22993 ( .A1(N7052), .A2(n19047), .B1(N7019), .B2(n23388), .ZN(
        n42960) );
  OAI21_X1 U22994 ( .B1(n22777), .B2(n7715), .A(n42970), .ZN(n6217) );
  AOI22_X1 U22995 ( .A1(N7051), .A2(n25170), .B1(N7018), .B2(n21784), .ZN(
        n42970) );
  OAI21_X1 U22996 ( .B1(n25335), .B2(n7719), .A(n42980), .ZN(n6218) );
  AOI22_X1 U22997 ( .A1(N7050), .A2(n24578), .B1(N7017), .B2(n26251), .ZN(
        n42980) );
  OAI21_X1 U22998 ( .B1(n20727), .B2(n7723), .A(n42990), .ZN(n6219) );
  AOI22_X1 U22999 ( .A1(N7049), .A2(n25175), .B1(N7016), .B2(n21782), .ZN(
        n42990) );
  OAI21_X1 U23000 ( .B1(n26697), .B2(n7728), .A(n43000), .ZN(n6220) );
  AOI22_X1 U23001 ( .A1(N7048), .A2(n19197), .B1(N7015), .B2(n26260), .ZN(
        n43000) );
  OAI21_X1 U23002 ( .B1(n21180), .B2(n8192), .A(n4125), .ZN(n61010) );
  AOI22_X1 U23003 ( .A1(N6443), .A2(n27170), .B1(N6410), .B2(n24303), .ZN(
        n4125) );
  OAI21_X1 U23004 ( .B1(n19297), .B2(n8200), .A(n4127), .ZN(n61030) );
  AOI22_X1 U23005 ( .A1(N6441), .A2(n19051), .B1(N6408), .B2(n268001), .ZN(
        n4127) );
  OAI21_X1 U23006 ( .B1(n20723), .B2(n8208), .A(n41290), .ZN(n61050) );
  AOI22_X1 U23007 ( .A1(N6439), .A2(n24579), .B1(N6406), .B2(n26802), .ZN(
        n41290) );
  OAI21_X1 U23008 ( .B1(n20726), .B2(n8212), .A(n41300), .ZN(n61060) );
  AOI22_X1 U23009 ( .A1(N6438), .A2(n27167), .B1(N6405), .B2(n24301), .ZN(
        n41300) );
  OAI21_X1 U23010 ( .B1(n25533), .B2(n8216), .A(n41310), .ZN(n61070) );
  AOI22_X1 U23011 ( .A1(N6437), .A2(n25181), .B1(N6404), .B2(n26259), .ZN(
        n41310) );
  OAI21_X1 U23012 ( .B1(n20729), .B2(n8220), .A(n41320), .ZN(n61080) );
  AOI22_X1 U23013 ( .A1(N6436), .A2(n27165), .B1(N6403), .B2(n26251), .ZN(
        n41320) );
  OAI21_X1 U23014 ( .B1(n21171), .B2(n8228), .A(n41340), .ZN(n61100) );
  AOI22_X1 U23015 ( .A1(N6434), .A2(n25559), .B1(N6401), .B2(n26260), .ZN(
        n41340) );
  OAI21_X1 U23016 ( .B1(n24943), .B2(n8232), .A(n41350), .ZN(n61110) );
  AOI22_X1 U23017 ( .A1(N6433), .A2(n19190), .B1(N6400), .B2(n20500), .ZN(
        n41350) );
  OAI21_X1 U23018 ( .B1(n21182), .B2(n8236), .A(n41360), .ZN(n61120) );
  AOI22_X1 U23019 ( .A1(N6432), .A2(n24556), .B1(N6399), .B2(n21781), .ZN(
        n41360) );
  OAI21_X1 U23020 ( .B1(n20728), .B2(n8240), .A(n41370), .ZN(n61130) );
  AOI22_X1 U23021 ( .A1(N6431), .A2(n24555), .B1(N6398), .B2(n24304), .ZN(
        n41370) );
  OAI21_X1 U23022 ( .B1(n21182), .B2(n8244), .A(n41380), .ZN(n6114) );
  AOI22_X1 U23023 ( .A1(N6430), .A2(n19191), .B1(N6397), .B2(n24298), .ZN(
        n41380) );
  OAI21_X1 U23024 ( .B1(n26690), .B2(n8732), .A(n39650), .ZN(n5997) );
  AOI22_X1 U23025 ( .A1(N5856), .A2(n21224), .B1(N5823), .B2(n21785), .ZN(
        n39650) );
  OAI21_X1 U23026 ( .B1(n24943), .B2(n8742), .A(n39670), .ZN(n5999) );
  AOI22_X1 U23027 ( .A1(N5854), .A2(n24556), .B1(N5821), .B2(n26245), .ZN(
        n39670) );
  OAI21_X1 U23028 ( .B1(n24947), .B2(n8747), .A(n39680), .ZN(n6000) );
  AOI22_X1 U23029 ( .A1(N5853), .A2(n25556), .B1(N5820), .B2(n26261), .ZN(
        n39680) );
  OAI21_X1 U23030 ( .B1(n21168), .B2(n8752), .A(n39690), .ZN(n6001) );
  AOI22_X1 U23031 ( .A1(N5852), .A2(n25561), .B1(N5819), .B2(n26257), .ZN(
        n39690) );
  OAI21_X1 U23032 ( .B1(n24954), .B2(n8757), .A(n39700), .ZN(n6002) );
  AOI22_X1 U23033 ( .A1(N5851), .A2(n24537), .B1(N5818), .B2(n21777), .ZN(
        n39700) );
  OAI21_X1 U23034 ( .B1(n25537), .B2(n8767), .A(n39720), .ZN(n6004) );
  AOI22_X1 U23035 ( .A1(N5849), .A2(n21215), .B1(N5816), .B2(n24300), .ZN(
        n39720) );
  OAI21_X1 U23036 ( .B1(n24949), .B2(n8772), .A(n39730), .ZN(n6005) );
  AOI22_X1 U23037 ( .A1(N5848), .A2(n19050), .B1(N5815), .B2(n21786), .ZN(
        n39730) );
  OAI21_X1 U23038 ( .B1(n21167), .B2(n8777), .A(n39740), .ZN(n6006) );
  AOI22_X1 U23039 ( .A1(N5847), .A2(n19047), .B1(N5814), .B2(n21779), .ZN(
        n39740) );
  OAI21_X1 U23040 ( .B1(n24951), .B2(n8782), .A(n39750), .ZN(n6007) );
  AOI22_X1 U23041 ( .A1(N5846), .A2(n22931), .B1(N5813), .B2(n23380), .ZN(
        n39750) );
  OAI21_X1 U23042 ( .B1(n22773), .B2(n8787), .A(n39760), .ZN(n6008) );
  AOI22_X1 U23043 ( .A1(N5845), .A2(n25179), .B1(N5812), .B2(n21789), .ZN(
        n39760) );
  OAI21_X1 U23044 ( .B1(n26701), .B2(n8796), .A(n39780), .ZN(n6010) );
  AOI22_X1 U23045 ( .A1(N5843), .A2(n22930), .B1(N5810), .B2(n23381), .ZN(
        n39780) );
  OAI21_X1 U23046 ( .B1(n20736), .B2(n9186), .A(n3830), .ZN(n59070) );
  AOI22_X1 U23047 ( .A1(N5352), .A2(n25178), .B1(N5319), .B2(n26266), .ZN(
        n3830) );
  OAI21_X1 U23048 ( .B1(n25342), .B2(n9191), .A(n3831), .ZN(n5908) );
  AOI22_X1 U23049 ( .A1(N5351), .A2(n25164), .B1(N5318), .B2(n26798), .ZN(
        n3831) );
  OAI21_X1 U23050 ( .B1(n20731), .B2(n9201), .A(n3833), .ZN(n5910) );
  AOI22_X1 U23051 ( .A1(N5349), .A2(n25166), .B1(N5316), .B2(n26282), .ZN(
        n3833) );
  OAI21_X1 U23052 ( .B1(n17090), .B2(n9211), .A(n3835), .ZN(n5912) );
  AOI22_X1 U23053 ( .A1(N5347), .A2(n25172), .B1(N5314), .B2(n21791), .ZN(
        n3835) );
  OAI21_X1 U23054 ( .B1(n19296), .B2(n9216), .A(n3836), .ZN(n5913) );
  AOI22_X1 U23055 ( .A1(N5346), .A2(n22940), .B1(N5313), .B2(n26283), .ZN(
        n3836) );
  OAI21_X1 U23056 ( .B1(n25339), .B2(n9221), .A(n3837), .ZN(n5914) );
  AOI22_X1 U23057 ( .A1(N5345), .A2(n25545), .B1(N5312), .B2(n26286), .ZN(
        n3837) );
  OAI21_X1 U23058 ( .B1(n20732), .B2(n9226), .A(n38380), .ZN(n5915) );
  AOI22_X1 U23059 ( .A1(N5344), .A2(n21198), .B1(N5311), .B2(n26270), .ZN(
        n38380) );
  OAI21_X1 U23060 ( .B1(n25526), .B2(n9236), .A(n38400), .ZN(n5917) );
  AOI22_X1 U23061 ( .A1(N5342), .A2(n24568), .B1(N5309), .B2(n24280), .ZN(
        n38400) );
  OAI21_X1 U23062 ( .B1(n26686), .B2(n9241), .A(n38410), .ZN(n5918) );
  AOI22_X1 U23063 ( .A1(N5341), .A2(n24572), .B1(N5308), .B2(n26792), .ZN(
        n38410) );
  OAI21_X1 U23064 ( .B1(n25122), .B2(n9246), .A(n38420), .ZN(n5919) );
  AOI22_X1 U23065 ( .A1(N5340), .A2(n24542), .B1(N5307), .B2(n26266), .ZN(
        n38420) );
  OAI21_X1 U23066 ( .B1(n26693), .B2(n9250), .A(n38430), .ZN(n5920) );
  AOI22_X1 U23067 ( .A1(N5339), .A2(n24575), .B1(N5306), .B2(n26265), .ZN(
        n38430) );
  OAI21_X1 U23068 ( .B1(n22774), .B2(n9261), .A(n38070), .ZN(n5891) );
  AOI22_X1 U23069 ( .A1(N5264), .A2(n21204), .B1(N5231), .B2(n20501), .ZN(
        n38070) );
  OAI21_X1 U23070 ( .B1(n26701), .B2(n9271), .A(n38090), .ZN(n58930) );
  AOI22_X1 U23071 ( .A1(N5262), .A2(n25167), .B1(N5229), .B2(n21778), .ZN(
        n38090) );
  OAI21_X1 U23072 ( .B1(n20724), .B2(n9276), .A(n3810), .ZN(n58940) );
  AOI22_X1 U23073 ( .A1(N5261), .A2(n27168), .B1(N5228), .B2(n26256), .ZN(
        n3810) );
  OAI21_X1 U23074 ( .B1(n19036), .B2(n9281), .A(n3811), .ZN(n58950) );
  AOI22_X1 U23075 ( .A1(N5260), .A2(n24579), .B1(N5227), .B2(n21783), .ZN(
        n3811) );
  OAI21_X1 U23076 ( .B1(n20730), .B2(n9286), .A(n3812), .ZN(n58960) );
  AOI22_X1 U23077 ( .A1(N5259), .A2(n24548), .B1(N5226), .B2(n21780), .ZN(
        n3812) );
  OAI21_X1 U23078 ( .B1(n25119), .B2(n9296), .A(n3814), .ZN(n58980) );
  AOI22_X1 U23079 ( .A1(N5257), .A2(n22933), .B1(N5224), .B2(n21789), .ZN(
        n3814) );
  OAI21_X1 U23080 ( .B1(n20725), .B2(n9301), .A(n3815), .ZN(n58990) );
  AOI22_X1 U23081 ( .A1(N5256), .A2(n25558), .B1(N5223), .B2(n24298), .ZN(
        n3815) );
  OAI21_X1 U23082 ( .B1(n19183), .B2(n9306), .A(n3816), .ZN(n59000) );
  AOI22_X1 U23083 ( .A1(N5255), .A2(n19192), .B1(N5222), .B2(n24307), .ZN(
        n3816) );
  OAI21_X1 U23084 ( .B1(n20727), .B2(n9311), .A(n3817), .ZN(n59010) );
  AOI22_X1 U23085 ( .A1(N5254), .A2(n25555), .B1(N5221), .B2(n24304), .ZN(
        n3817) );
  OAI21_X1 U23086 ( .B1(n26696), .B2(n9316), .A(n3818), .ZN(n59020) );
  AOI22_X1 U23087 ( .A1(N5253), .A2(n21201), .B1(N5220), .B2(n24301), .ZN(
        n3818) );
  OAI21_X1 U23088 ( .B1(n26698), .B2(n9326), .A(n3820), .ZN(n59040) );
  AOI22_X1 U23089 ( .A1(N5251), .A2(n24553), .B1(N5218), .B2(n21775), .ZN(
        n3820) );
  OAI21_X1 U23090 ( .B1(n25333), .B2(n9330), .A(n3821), .ZN(n59050) );
  AOI22_X1 U23091 ( .A1(N5250), .A2(n24540), .B1(N5217), .B2(n26252), .ZN(
        n3821) );
  OAI21_X1 U23092 ( .B1(n20738), .B2(n9715), .A(n36720), .ZN(n5801) );
  AOI22_X1 U23093 ( .A1(N4742), .A2(n21193), .B1(N4709), .B2(n26267), .ZN(
        n36720) );
  OAI21_X1 U23094 ( .B1(n25529), .B2(n9720), .A(n36730), .ZN(n5802) );
  AOI22_X1 U23095 ( .A1(N4741), .A2(n24567), .B1(N4708), .B2(n26269), .ZN(
        n36730) );
  OAI21_X1 U23096 ( .B1(n26692), .B2(n9730), .A(n36750), .ZN(n5804) );
  AOI22_X1 U23097 ( .A1(N4739), .A2(n24576), .B1(N4706), .B2(n21807), .ZN(
        n36750) );
  OAI21_X1 U23098 ( .B1(n20735), .B2(n9740), .A(n36770), .ZN(n5806) );
  AOI22_X1 U23099 ( .A1(N4737), .A2(n24545), .B1(N4704), .B2(n24295), .ZN(
        n36770) );
  OAI21_X1 U23100 ( .B1(n26686), .B2(n9745), .A(n36780), .ZN(n5807) );
  AOI22_X1 U23101 ( .A1(N4736), .A2(n25548), .B1(N4703), .B2(n21812), .ZN(
        n36780) );
  OAI21_X1 U23102 ( .B1(n19090), .B2(n9750), .A(n36790), .ZN(n5808) );
  AOI22_X1 U23103 ( .A1(N4735), .A2(n21218), .B1(N4702), .B2(n20503), .ZN(
        n36790) );
  OAI21_X1 U23104 ( .B1(n24956), .B2(n9755), .A(n36800), .ZN(n5809) );
  AOI22_X1 U23105 ( .A1(N4734), .A2(n21211), .B1(N4701), .B2(n24295), .ZN(
        n36800) );
  OAI21_X1 U23106 ( .B1(n19089), .B2(n9765), .A(n36820), .ZN(n58110) );
  AOI22_X1 U23107 ( .A1(N4732), .A2(n19046), .B1(N4699), .B2(n20503), .ZN(
        n36820) );
  OAI21_X1 U23108 ( .B1(n19296), .B2(n9770), .A(n3683), .ZN(n58120) );
  AOI22_X1 U23109 ( .A1(N4731), .A2(n27258), .B1(N4698), .B2(n21809), .ZN(
        n3683) );
  OAI21_X1 U23110 ( .B1(n25341), .B2(n9775), .A(n3684), .ZN(n58130) );
  AOI22_X1 U23111 ( .A1(N4730), .A2(n25165), .B1(N4697), .B2(n26268), .ZN(
        n3684) );
  OAI21_X1 U23112 ( .B1(n24958), .B2(n9780), .A(n3685), .ZN(n58140) );
  AOI22_X1 U23113 ( .A1(N4729), .A2(n25173), .B1(N4696), .B2(n21797), .ZN(
        n3685) );
  OAI21_X1 U23114 ( .B1(n26695), .B2(n9784), .A(n3686), .ZN(n58150) );
  AOI22_X1 U23115 ( .A1(N4728), .A2(n19195), .B1(N4695), .B2(n26285), .ZN(
        n3686) );
  OAI21_X1 U23116 ( .B1(n21173), .B2(n10249), .A(n35130), .ZN(n5696) );
  AOI22_X1 U23117 ( .A1(N4142), .A2(n24581), .B1(N4109), .B2(n24292), .ZN(
        n35130) );
  OAI21_X1 U23118 ( .B1(n26695), .B2(n10259), .A(n3515), .ZN(n5698) );
  AOI22_X1 U23119 ( .A1(N4140), .A2(n19048), .B1(N4107), .B2(n20504), .ZN(
        n3515) );
  OAI21_X1 U23120 ( .B1(n20738), .B2(n10269), .A(n3517), .ZN(n5700) );
  AOI22_X1 U23121 ( .A1(N4138), .A2(n24582), .B1(N4105), .B2(n26792), .ZN(
        n3517) );
  OAI21_X1 U23122 ( .B1(n20736), .B2(n10274), .A(n3518), .ZN(n5701) );
  AOI22_X1 U23123 ( .A1(N4137), .A2(n27255), .B1(N4104), .B2(n24282), .ZN(
        n3518) );
  OAI21_X1 U23124 ( .B1(n25530), .B2(n10279), .A(n3519), .ZN(n5702) );
  AOI22_X1 U23125 ( .A1(N4136), .A2(n25171), .B1(N4103), .B2(n26284), .ZN(
        n3519) );
  OAI21_X1 U23126 ( .B1(n21165), .B2(n10284), .A(n3520), .ZN(n5703) );
  AOI22_X1 U23127 ( .A1(N4135), .A2(n27253), .B1(N4102), .B2(n26268), .ZN(
        n3520) );
  OAI21_X1 U23128 ( .B1(n21164), .B2(n10294), .A(n3522), .ZN(n5705) );
  AOI22_X1 U23129 ( .A1(N4133), .A2(n25546), .B1(N4100), .B2(n26285), .ZN(
        n3522) );
  OAI21_X1 U23130 ( .B1(n21175), .B2(n10299), .A(n3523), .ZN(n5706) );
  AOI22_X1 U23131 ( .A1(N4132), .A2(n19186), .B1(N4099), .B2(n23410), .ZN(
        n3523) );
  OAI21_X1 U23132 ( .B1(n21175), .B2(n10304), .A(n3524), .ZN(n5707) );
  AOI22_X1 U23133 ( .A1(N4131), .A2(n24573), .B1(N4098), .B2(n21798), .ZN(
        n3524) );
  OAI21_X1 U23134 ( .B1(n20732), .B2(n10309), .A(n3525), .ZN(n5708) );
  AOI22_X1 U23135 ( .A1(N4130), .A2(n24573), .B1(N4097), .B2(n24291), .ZN(
        n3525) );
  OAI21_X1 U23136 ( .B1(n24952), .B2(n10314), .A(n3526), .ZN(n5709) );
  AOI22_X1 U23137 ( .A1(N4129), .A2(n19187), .B1(N4096), .B2(n24279), .ZN(
        n3526) );
  OAI21_X1 U23138 ( .B1(n24952), .B2(n10822), .A(n3354), .ZN(n55920) );
  AOI22_X1 U23139 ( .A1(N3545), .A2(n21219), .B1(N3512), .B2(n26284), .ZN(
        n3354) );
  OAI21_X1 U23140 ( .B1(n26689), .B2(n10830), .A(n3356), .ZN(n55940) );
  AOI22_X1 U23141 ( .A1(N3543), .A2(n24568), .B1(N3510), .B2(n26262), .ZN(
        n3356) );
  OAI21_X1 U23142 ( .B1(n20739), .B2(n10834), .A(n3357), .ZN(n55950) );
  AOI22_X1 U23143 ( .A1(N3542), .A2(n25543), .B1(N3509), .B2(n26286), .ZN(
        n3357) );
  OAI21_X1 U23144 ( .B1(n21156), .B2(n10838), .A(n3358), .ZN(n55960) );
  AOI22_X1 U23145 ( .A1(N3541), .A2(n25547), .B1(N3508), .B2(n26282), .ZN(
        n3358) );
  OAI21_X1 U23146 ( .B1(n24956), .B2(n10842), .A(n3359), .ZN(n55970) );
  AOI22_X1 U23147 ( .A1(N3540), .A2(n24541), .B1(N3507), .B2(n21793), .ZN(
        n3359) );
  OAI21_X1 U23148 ( .B1(n25534), .B2(n10850), .A(n3361), .ZN(n55990) );
  AOI22_X1 U23149 ( .A1(N3538), .A2(n21212), .B1(N3505), .B2(n24283), .ZN(
        n3361) );
  OAI21_X1 U23150 ( .B1(n17090), .B2(n10854), .A(n3362), .ZN(n56000) );
  AOI22_X1 U23151 ( .A1(N3537), .A2(n19049), .B1(N3504), .B2(n21809), .ZN(
        n3362) );
  OAI21_X1 U23152 ( .B1(n21157), .B2(n10858), .A(n3363), .ZN(n56010) );
  AOI22_X1 U23153 ( .A1(N3536), .A2(n19046), .B1(N3503), .B2(n21796), .ZN(
        n3363) );
  OAI21_X1 U23154 ( .B1(n24958), .B2(n10862), .A(n33640), .ZN(n56020) );
  AOI22_X1 U23155 ( .A1(N3535), .A2(n22937), .B1(N3502), .B2(n23396), .ZN(
        n33640) );
  OAI21_X1 U23156 ( .B1(n22769), .B2(n10866), .A(n33650), .ZN(n56030) );
  AOI22_X1 U23157 ( .A1(N3534), .A2(n25177), .B1(N3501), .B2(n21814), .ZN(
        n33650) );
  OAI21_X1 U23158 ( .B1(n22766), .B2(n10875), .A(n33670), .ZN(n56050) );
  AOI22_X1 U23159 ( .A1(N3532), .A2(n22936), .B1(N3499), .B2(n23395), .ZN(
        n33670) );
  OAI21_X1 U23160 ( .B1(n22770), .B2(n11339), .A(n3187), .ZN(n54860) );
  AOI22_X1 U23161 ( .A1(N2954), .A2(n21195), .B1(N2921), .B2(n267901), .ZN(
        n3187) );
  OAI21_X1 U23162 ( .B1(n22767), .B2(n11349), .A(n3189), .ZN(n54880) );
  AOI22_X1 U23163 ( .A1(N2952), .A2(n25163), .B1(N2919), .B2(n21794), .ZN(
        n3189) );
  OAI21_X1 U23164 ( .B1(n20739), .B2(n11354), .A(n3190), .ZN(n54890) );
  AOI22_X1 U23165 ( .A1(N2951), .A2(n27256), .B1(N2918), .B2(n26281), .ZN(
        n3190) );
  OAI21_X1 U23166 ( .B1(n19037), .B2(n11359), .A(n3191), .ZN(n5490) );
  AOI22_X1 U23167 ( .A1(N2950), .A2(n24582), .B1(N2917), .B2(n21808), .ZN(
        n3191) );
  OAI21_X1 U23168 ( .B1(n20731), .B2(n11364), .A(n3192), .ZN(n5491) );
  AOI22_X1 U23169 ( .A1(N2949), .A2(n24565), .B1(N2916), .B2(n21795), .ZN(
        n3192) );
  OAI21_X1 U23170 ( .B1(n25121), .B2(n11374), .A(n3194), .ZN(n5493) );
  AOI22_X1 U23171 ( .A1(N2947), .A2(n22939), .B1(N2914), .B2(n21813), .ZN(
        n3194) );
  OAI21_X1 U23172 ( .B1(n20735), .B2(n11379), .A(n3195), .ZN(n5494) );
  AOI22_X1 U23173 ( .A1(N2946), .A2(n25545), .B1(N2913), .B2(n24280), .ZN(
        n3195) );
  OAI21_X1 U23174 ( .B1(n19181), .B2(n11384), .A(n31960), .ZN(n5495) );
  AOI22_X1 U23175 ( .A1(N2945), .A2(n19188), .B1(N2912), .B2(n24294), .ZN(
        n31960) );
  OAI21_X1 U23176 ( .B1(n20733), .B2(n11389), .A(n31970), .ZN(n5496) );
  AOI22_X1 U23177 ( .A1(N2944), .A2(n25542), .B1(N2911), .B2(n24292), .ZN(
        n31970) );
  OAI21_X1 U23178 ( .B1(n26692), .B2(n11394), .A(n31980), .ZN(n5497) );
  AOI22_X1 U23179 ( .A1(N2943), .A2(n21192), .B1(N2910), .B2(n24283), .ZN(
        n31980) );
  OAI21_X1 U23180 ( .B1(n26687), .B2(n11404), .A(n32000), .ZN(n5499) );
  AOI22_X1 U23181 ( .A1(N2941), .A2(n24569), .B1(N2908), .B2(n21792), .ZN(
        n32000) );
  OAI21_X1 U23182 ( .B1(n25338), .B2(n11408), .A(n32010), .ZN(n5500) );
  AOI22_X1 U23183 ( .A1(N2940), .A2(n24545), .B1(N2907), .B2(n26269), .ZN(
        n32010) );
  NAND2_X1 U23184 ( .A1(n52250), .A2(n52260), .ZN(mul_outcome[141]) );
  AOI221_X1 U23185 ( .B1(n24400), .B2(n17401), .C1(n17116), .C2(n17377), .A(
        n27738), .ZN(n52250) );
  AOI221_X1 U23186 ( .B1(n19234), .B2(n17461), .C1(n27032), .C2(n17449), .A(
        n27754), .ZN(n52260) );
  INV_X1 U23187 ( .A(n52280), .ZN(n27738) );
  NAND2_X1 U23188 ( .A1(n5126), .A2(n5127), .ZN(mul_outcome[162]) );
  AOI221_X1 U23189 ( .B1(n22430), .B2(n17293), .C1(n19086), .C2(n17281), .A(
        n27732), .ZN(n5126) );
  AOI221_X1 U23190 ( .B1(n25655), .B2(n17365), .C1(n19248), .C2(n17353), .A(
        n27773), .ZN(n5127) );
  INV_X1 U23191 ( .A(n5129), .ZN(n27732) );
  OAI21_X1 U23192 ( .B1(n25531), .B2(n29190), .A(n4451), .ZN(n6311) );
  AOI22_X1 U23193 ( .A1(N7654), .A2(n25563), .B1(N7621), .B2(n26258), .ZN(
        n4451) );
  OAI21_X1 U23194 ( .B1(n25120), .B2(n2931), .A(n4454), .ZN(n6314) );
  AOI22_X1 U23195 ( .A1(N7651), .A2(n25169), .B1(N7618), .B2(n21788), .ZN(
        n4454) );
  OAI21_X1 U23196 ( .B1(n25333), .B2(n2939), .A(n4456), .ZN(n6316) );
  AOI22_X1 U23197 ( .A1(N7649), .A2(n24548), .B1(N7616), .B2(n26805), .ZN(
        n4456) );
  OAI21_X1 U23198 ( .B1(n25336), .B2(n29590), .A(n4461), .ZN(n63210) );
  AOI22_X1 U23199 ( .A1(N7644), .A2(n25555), .B1(N7611), .B2(n19262), .ZN(
        n4461) );
  OAI21_X1 U23200 ( .B1(n21172), .B2(n7679), .A(n4288), .ZN(n6208) );
  AOI22_X1 U23201 ( .A1(N7060), .A2(n24552), .B1(N7027), .B2(n26256), .ZN(
        n4288) );
  OAI21_X1 U23202 ( .B1(n25537), .B2(n7687), .A(n4290), .ZN(n6210) );
  AOI22_X1 U23203 ( .A1(N7058), .A2(n24540), .B1(N7025), .B2(n21777), .ZN(
        n4290) );
  OAI21_X1 U23204 ( .B1(n19183), .B2(n77070), .A(n4295), .ZN(n6215) );
  AOI22_X1 U23205 ( .A1(N7053), .A2(n25180), .B1(N7020), .B2(n26253), .ZN(
        n4295) );
  OAI21_X1 U23206 ( .B1(n19036), .B2(n8196), .A(n4126), .ZN(n61020) );
  AOI22_X1 U23207 ( .A1(N6442), .A2(n24547), .B1(N6409), .B2(n26254), .ZN(
        n4126) );
  OAI21_X1 U23208 ( .B1(n19087), .B2(n8204), .A(n41280), .ZN(n61040) );
  AOI22_X1 U23209 ( .A1(N6440), .A2(n25176), .B1(N6407), .B2(n26804), .ZN(
        n41280) );
  OAI21_X1 U23210 ( .B1(n19088), .B2(n8224), .A(n41330), .ZN(n61090) );
  AOI22_X1 U23211 ( .A1(N6435), .A2(n21205), .B1(N6402), .B2(n23380), .ZN(
        n41330) );
  OAI21_X1 U23212 ( .B1(n25532), .B2(n8249), .A(n41390), .ZN(n6115) );
  AOI22_X1 U23213 ( .A1(N6429), .A2(n21208), .B1(N6396), .B2(n21785), .ZN(
        n41390) );
  OAI21_X1 U23214 ( .B1(n21183), .B2(n8727), .A(n39640), .ZN(n59960) );
  AOI22_X1 U23215 ( .A1(N5857), .A2(n24559), .B1(N5824), .B2(n21790), .ZN(
        n39640) );
  OAI21_X1 U23216 ( .B1(n21167), .B2(n8737), .A(n39660), .ZN(n5998) );
  AOI22_X1 U23217 ( .A1(N5855), .A2(n19194), .B1(N5822), .B2(n26250), .ZN(
        n39660) );
  OAI21_X1 U23218 ( .B1(n25119), .B2(n8762), .A(n39710), .ZN(n6003) );
  AOI22_X1 U23219 ( .A1(N5850), .A2(n25566), .B1(N5817), .B2(n21781), .ZN(
        n39710) );
  OAI21_X1 U23220 ( .B1(n25334), .B2(n8792), .A(n39770), .ZN(n6009) );
  AOI22_X1 U23221 ( .A1(N5844), .A2(n25168), .B1(N5811), .B2(n26801), .ZN(
        n39770) );
  OAI21_X1 U23222 ( .B1(n25526), .B2(n9181), .A(n3829), .ZN(n59060) );
  AOI22_X1 U23223 ( .A1(N5353), .A2(n25560), .B1(N5320), .B2(n26283), .ZN(
        n3829) );
  OAI21_X1 U23224 ( .B1(n25122), .B2(n9196), .A(n3832), .ZN(n5909) );
  AOI22_X1 U23225 ( .A1(N5350), .A2(n25166), .B1(N5317), .B2(n21811), .ZN(
        n3832) );
  OAI21_X1 U23226 ( .B1(n25338), .B2(n9206), .A(n3834), .ZN(n5911) );
  AOI22_X1 U23227 ( .A1(N5348), .A2(n24564), .B1(N5315), .B2(n26799), .ZN(
        n3834) );
  OAI21_X1 U23228 ( .B1(n25342), .B2(n9231), .A(n38390), .ZN(n5916) );
  AOI22_X1 U23229 ( .A1(N5343), .A2(n25542), .B1(N5310), .B2(n19263), .ZN(
        n38390) );
  OAI21_X1 U23230 ( .B1(n25335), .B2(n9266), .A(n38080), .ZN(n58920) );
  AOI22_X1 U23231 ( .A1(N5263), .A2(n25559), .B1(N5230), .B2(n23381), .ZN(
        n38080) );
  OAI21_X1 U23232 ( .B1(n25533), .B2(n9291), .A(n3813), .ZN(n58970) );
  AOI22_X1 U23233 ( .A1(N5258), .A2(n25182), .B1(N5225), .B2(n26248), .ZN(
        n3813) );
  OAI21_X1 U23234 ( .B1(n25538), .B2(n9321), .A(n3819), .ZN(n59030) );
  AOI22_X1 U23235 ( .A1(N5252), .A2(n25557), .B1(N5219), .B2(n20500), .ZN(
        n3819) );
  OAI21_X1 U23236 ( .B1(n21165), .B2(n9725), .A(n36740), .ZN(n5803) );
  AOI22_X1 U23237 ( .A1(N4740), .A2(n24570), .B1(N4707), .B2(n26281), .ZN(
        n36740) );
  OAI21_X1 U23238 ( .B1(n25534), .B2(n9735), .A(n36760), .ZN(n5805) );
  AOI22_X1 U23239 ( .A1(N4738), .A2(n24544), .B1(N4705), .B2(n21793), .ZN(
        n36760) );
  OAI21_X1 U23240 ( .B1(n19181), .B2(n9760), .A(n36810), .ZN(n58100) );
  AOI22_X1 U23241 ( .A1(N4733), .A2(n25178), .B1(N4700), .B2(n26270), .ZN(
        n36810) );
  OAI21_X1 U23242 ( .B1(n19037), .B2(n10254), .A(n35140), .ZN(n5697) );
  AOI22_X1 U23243 ( .A1(N4141), .A2(n24565), .B1(N4108), .B2(n26791), .ZN(
        n35140) );
  OAI21_X1 U23244 ( .B1(n19089), .B2(n10264), .A(n3516), .ZN(n5699) );
  AOI22_X1 U23245 ( .A1(N4139), .A2(n25174), .B1(N4106), .B2(n26262), .ZN(
        n3516) );
  OAI21_X1 U23246 ( .B1(n19090), .B2(n10289), .A(n3521), .ZN(n5704) );
  AOI22_X1 U23247 ( .A1(N4134), .A2(n21196), .B1(N4101), .B2(n23395), .ZN(
        n3521) );
  OAI21_X1 U23248 ( .B1(n25529), .B2(n10318), .A(n3527), .ZN(n5710) );
  AOI22_X1 U23249 ( .A1(N4128), .A2(n21199), .B1(N4095), .B2(n21810), .ZN(
        n3527) );
  OAI21_X1 U23250 ( .B1(n21176), .B2(n10818), .A(n3353), .ZN(n55910) );
  AOI22_X1 U23251 ( .A1(N3546), .A2(n24576), .B1(N3513), .B2(n21813), .ZN(
        n3353) );
  OAI21_X1 U23252 ( .B1(n21156), .B2(n10826), .A(n3355), .ZN(n55930) );
  AOI22_X1 U23253 ( .A1(N3544), .A2(n19193), .B1(N3511), .B2(n26267), .ZN(
        n3355) );
  OAI21_X1 U23254 ( .B1(n25121), .B2(n10846), .A(n3360), .ZN(n55980) );
  AOI22_X1 U23255 ( .A1(N3539), .A2(n25564), .B1(N3506), .B2(n21797), .ZN(
        n3360) );
  OAI21_X1 U23256 ( .B1(n25339), .B2(n10870), .A(n33660), .ZN(n56040) );
  AOI22_X1 U23257 ( .A1(N3533), .A2(n25164), .B1(N3500), .B2(n26279), .ZN(
        n33660) );
  OAI21_X1 U23258 ( .B1(n25341), .B2(n11344), .A(n3188), .ZN(n54870) );
  AOI22_X1 U23259 ( .A1(N2953), .A2(n25546), .B1(N2920), .B2(n23396), .ZN(
        n3188) );
  OAI21_X1 U23260 ( .B1(n25530), .B2(n11369), .A(n3193), .ZN(n5492) );
  AOI22_X1 U23261 ( .A1(N2948), .A2(n25172), .B1(N2915), .B2(n26265), .ZN(
        n3193) );
  OAI21_X1 U23262 ( .B1(n25535), .B2(n11399), .A(n31990), .ZN(n5498) );
  AOI22_X1 U23263 ( .A1(N2942), .A2(n25544), .B1(N2909), .B2(n26279), .ZN(
        n31990) );
  NAND3_X1 U23264 ( .A1(n47940), .A2(n47950), .A3(n47960), .ZN(mul_outcome[81]) );
  AOI22_X1 U23265 ( .A1(n21185), .A2(n17719), .B1(n20694), .B2(n17671), .ZN(
        n47940) );
  AOI22_X1 U23266 ( .A1(n27103), .A2(n17743), .B1(n21189), .B2(n17731), .ZN(
        n47950) );
  AOI221_X1 U23267 ( .B1(n26078), .B2(n17683), .C1(n23975), .C2(n17659), .A(
        n27762), .ZN(n47960) );
  NAND3_X1 U23268 ( .A1(n4806), .A2(n4807), .A3(n4808), .ZN(mul_outcome[79])
         );
  AOI22_X1 U23269 ( .A1(n25755), .A2(n17723), .B1(n23725), .B2(n17675), .ZN(
        n4806) );
  AOI22_X1 U23270 ( .A1(n27101), .A2(n17747), .B1(n25747), .B2(n17735), .ZN(
        n4807) );
  AOI221_X1 U23271 ( .B1(n265201), .B2(n17687), .C1(n23974), .C2(n17663), .A(
        n27764), .ZN(n4808) );
  NAND3_X1 U23272 ( .A1(n47900), .A2(n47910), .A3(n47920), .ZN(mul_outcome[82]) );
  AOI22_X1 U23273 ( .A1(n25759), .A2(n17717), .B1(n20688), .B2(n17669), .ZN(
        n47900) );
  AOI22_X1 U23274 ( .A1(n27104), .A2(n17741), .B1(n21178), .B2(n17729), .ZN(
        n47910) );
  AOI221_X1 U23275 ( .B1(n26305), .B2(n17681), .C1(n22880), .C2(n17657), .A(
        n27761), .ZN(n47920) );
  NAND3_X1 U23276 ( .A1(n54000), .A2(n5401), .A3(n5402), .ZN(mul_outcome[103])
         );
  AOI221_X1 U23277 ( .B1(n23967), .B2(n17573), .C1(n24396), .C2(n17561), .A(
        n27756), .ZN(n5402) );
  AOI22_X1 U23278 ( .A1(n21596), .A2(n17621), .B1(n21602), .B2(n17609), .ZN(
        n54000) );
  AOI22_X1 U23279 ( .A1(n19302), .A2(n17645), .B1(n19300), .B2(n17633), .ZN(
        n5401) );
  NAND3_X1 U23280 ( .A1(n5408), .A2(n5409), .A3(n5410), .ZN(mul_outcome[101])
         );
  AOI221_X1 U23281 ( .B1(n22677), .B2(n17577), .C1(n26402), .C2(n17565), .A(
        n27758), .ZN(n5410) );
  AOI22_X1 U23282 ( .A1(n21947), .A2(n17625), .B1(n21938), .B2(n17613), .ZN(
        n5408) );
  AOI22_X1 U23283 ( .A1(n24167), .A2(n17649), .B1(n24163), .B2(n17637), .ZN(
        n5409) );
  OAI21_X1 U23284 ( .B1(n24013), .B2(n2432), .A(n44760), .ZN(n63260) );
  AOI22_X1 U23285 ( .A1(N7743), .A2(n17081), .B1(N7710), .B2(n20575), .ZN(
        n44760) );
  OAI21_X1 U23286 ( .B1(n24005), .B2(n2556), .A(n44770), .ZN(n63270) );
  AOI22_X1 U23287 ( .A1(N7742), .A2(n25752), .B1(N7709), .B2(n20872), .ZN(
        n44770) );
  OAI21_X1 U23288 ( .B1(n25013), .B2(n265000), .A(n44780), .ZN(n63280) );
  AOI22_X1 U23289 ( .A1(N7741), .A2(n20793), .B1(N7708), .B2(n26387), .ZN(
        n44780) );
  OAI21_X1 U23290 ( .B1(n25013), .B2(n265400), .A(n44790), .ZN(n63290) );
  AOI22_X1 U23291 ( .A1(N7740), .A2(n25751), .B1(N7707), .B2(n21963), .ZN(
        n44790) );
  OAI21_X1 U23292 ( .B1(n24011), .B2(n268800), .A(n44800), .ZN(n63300) );
  AOI22_X1 U23293 ( .A1(N7739), .A2(n25004), .B1(N7706), .B2(n26386), .ZN(
        n44800) );
  OAI21_X1 U23294 ( .B1(n24003), .B2(n278200), .A(n44810), .ZN(n63310) );
  AOI22_X1 U23295 ( .A1(N7738), .A2(n22724), .B1(N7705), .B2(n25216), .ZN(
        n44810) );
  OAI21_X1 U23296 ( .B1(n25362), .B2(n278600), .A(n44820), .ZN(n63320) );
  AOI22_X1 U23297 ( .A1(N7737), .A2(n25753), .B1(N7704), .B2(n21960), .ZN(
        n44820) );
  OAI21_X1 U23298 ( .B1(n25016), .B2(n28200), .A(n44830), .ZN(n6333) );
  AOI22_X1 U23299 ( .A1(N7736), .A2(n20802), .B1(N7703), .B2(n26398), .ZN(
        n44830) );
  OAI21_X1 U23300 ( .B1(n26636), .B2(n2884), .A(n44840), .ZN(n6334) );
  AOI22_X1 U23301 ( .A1(N7735), .A2(n22731), .B1(N7702), .B2(n25220), .ZN(
        n44840) );
  OAI21_X1 U23302 ( .B1(n19277), .B2(n2888), .A(n4485), .ZN(n6335) );
  AOI22_X1 U23303 ( .A1(N7734), .A2(n24735), .B1(N7701), .B2(n25068), .ZN(
        n4485) );
  OAI21_X1 U23304 ( .B1(n21003), .B2(n2892), .A(n4486), .ZN(n6336) );
  AOI22_X1 U23305 ( .A1(N7733), .A2(n20524), .B1(N7700), .B2(n25074), .ZN(
        n4486) );
  OAI21_X1 U23306 ( .B1(n24821), .B2(n2896), .A(n4487), .ZN(n6337) );
  AOI22_X1 U23307 ( .A1(N7732), .A2(n24066), .B1(N7699), .B2(n26396), .ZN(
        n4487) );
  OAI21_X1 U23308 ( .B1(n26636), .B2(n2900), .A(n4488), .ZN(n6338) );
  AOI22_X1 U23309 ( .A1(N7731), .A2(n20797), .B1(N7698), .B2(n25214), .ZN(
        n4488) );
  OAI21_X1 U23310 ( .B1(n19277), .B2(n2904), .A(n4489), .ZN(n6339) );
  AOI22_X1 U23311 ( .A1(N7730), .A2(n20526), .B1(N7697), .B2(n25206), .ZN(
        n4489) );
  OAI21_X1 U23312 ( .B1(n22878), .B2(n29090), .A(n4490), .ZN(n6340) );
  AOI22_X1 U23313 ( .A1(N7729), .A2(n24075), .B1(N7696), .B2(n21959), .ZN(
        n4490) );
  OAI21_X1 U23314 ( .B1(n25363), .B2(n7592), .A(n43080), .ZN(n6221) );
  AOI22_X1 U23315 ( .A1(N7144), .A2(n24737), .B1(N7111), .B2(n21963), .ZN(
        n43080) );
  OAI21_X1 U23316 ( .B1(n24013), .B2(n7597), .A(n43090), .ZN(n6222) );
  AOI22_X1 U23317 ( .A1(N7143), .A2(n24070), .B1(N7110), .B2(n20576), .ZN(
        n43090) );
  OAI21_X1 U23318 ( .B1(n24005), .B2(n7602), .A(n43100), .ZN(n6223) );
  AOI22_X1 U23319 ( .A1(N7142), .A2(n25744), .B1(N7109), .B2(n24771), .ZN(
        n43100) );
  OAI21_X1 U23320 ( .B1(n25014), .B2(n76070), .A(n43110), .ZN(n6224) );
  AOI22_X1 U23321 ( .A1(N7141), .A2(n25112), .B1(N7108), .B2(n21962), .ZN(
        n43110) );
  OAI21_X1 U23322 ( .B1(n25243), .B2(n76120), .A(n43120), .ZN(n6225) );
  AOI22_X1 U23323 ( .A1(N7140), .A2(n24078), .B1(N7107), .B2(n21965), .ZN(
        n43120) );
  OAI21_X1 U23324 ( .B1(n24010), .B2(n76170), .A(n43130), .ZN(n6226) );
  AOI22_X1 U23325 ( .A1(N7139), .A2(n25743), .B1(N7106), .B2(n25215), .ZN(
        n43130) );
  OAI21_X1 U23326 ( .B1(n24002), .B2(n76220), .A(n43140), .ZN(n6227) );
  AOI22_X1 U23327 ( .A1(N7138), .A2(n20525), .B1(N7105), .B2(n26388), .ZN(
        n43140) );
  OAI21_X1 U23328 ( .B1(n24821), .B2(n7627), .A(n43150), .ZN(n62280) );
  AOI22_X1 U23329 ( .A1(N7137), .A2(n20799), .B1(N7104), .B2(n20573), .ZN(
        n43150) );
  OAI21_X1 U23330 ( .B1(n26922), .B2(n7632), .A(n43160), .ZN(n62290) );
  AOI22_X1 U23331 ( .A1(N7136), .A2(n20926), .B1(N7103), .B2(n26398), .ZN(
        n43160) );
  OAI21_X1 U23332 ( .B1(n19278), .B2(n7637), .A(n4317), .ZN(n62300) );
  AOI22_X1 U23333 ( .A1(N7135), .A2(n25114), .B1(N7102), .B2(n24774), .ZN(
        n4317) );
  OAI21_X1 U23334 ( .B1(n26632), .B2(n76420), .A(n4318), .ZN(n62310) );
  AOI22_X1 U23335 ( .A1(N7134), .A2(n24996), .B1(N7101), .B2(n25074), .ZN(
        n4318) );
  OAI21_X1 U23336 ( .B1(n20619), .B2(n76470), .A(n4319), .ZN(n62320) );
  AOI22_X1 U23337 ( .A1(N7133), .A2(n26654), .B1(N7100), .B2(n21961), .ZN(
        n4319) );
  OAI21_X1 U23338 ( .B1(n22877), .B2(n76520), .A(n4320), .ZN(n62330) );
  AOI22_X1 U23339 ( .A1(N7132), .A2(n25745), .B1(N7099), .B2(n25222), .ZN(
        n4320) );
  OAI21_X1 U23340 ( .B1(n19278), .B2(n76570), .A(n4321), .ZN(n62340) );
  AOI22_X1 U23341 ( .A1(N7131), .A2(n22723), .B1(N7098), .B2(n21959), .ZN(
        n4321) );
  OAI21_X1 U23342 ( .B1(n26632), .B2(n7661), .A(n4322), .ZN(n62350) );
  AOI22_X1 U23343 ( .A1(N7130), .A2(n25742), .B1(N7097), .B2(n25204), .ZN(
        n4322) );
  OAI21_X1 U23344 ( .B1(n25014), .B2(n8113), .A(n41470), .ZN(n6116) );
  AOI22_X1 U23345 ( .A1(N6532), .A2(n19289), .B1(N6499), .B2(n26394), .ZN(
        n41470) );
  OAI21_X1 U23346 ( .B1(n26634), .B2(n8118), .A(n41480), .ZN(n6117) );
  AOI22_X1 U23347 ( .A1(N6531), .A2(n24079), .B1(N6498), .B2(n21964), .ZN(
        n41480) );
  OAI21_X1 U23348 ( .B1(n24014), .B2(n8123), .A(n4149), .ZN(n6118) );
  AOI22_X1 U23349 ( .A1(N6530), .A2(n19033), .B1(N6497), .B2(n26387), .ZN(
        n4149) );
  OAI21_X1 U23350 ( .B1(n24006), .B2(n8128), .A(n4150), .ZN(n6119) );
  AOI22_X1 U23351 ( .A1(N6529), .A2(n19287), .B1(N6496), .B2(n20873), .ZN(
        n4150) );
  OAI21_X1 U23352 ( .B1(n25362), .B2(n8133), .A(n4151), .ZN(n6120) );
  AOI22_X1 U23353 ( .A1(N6528), .A2(n25752), .B1(N6495), .B2(n24771), .ZN(
        n4151) );
  OAI21_X1 U23354 ( .B1(n26634), .B2(n8138), .A(n4152), .ZN(n6121) );
  AOI22_X1 U23355 ( .A1(N6527), .A2(n25745), .B1(N6494), .B2(n26397), .ZN(
        n4152) );
  OAI21_X1 U23356 ( .B1(n24010), .B2(n8143), .A(n4153), .ZN(n6122) );
  AOI22_X1 U23357 ( .A1(N6526), .A2(n20801), .B1(N6493), .B2(n20572), .ZN(
        n4153) );
  OAI21_X1 U23358 ( .B1(n24003), .B2(n8148), .A(n4154), .ZN(n6123) );
  AOI22_X1 U23359 ( .A1(N6525), .A2(n20792), .B1(N6492), .B2(n20867), .ZN(
        n4154) );
  OAI21_X1 U23360 ( .B1(n20620), .B2(n8153), .A(n4155), .ZN(n6124) );
  AOI22_X1 U23361 ( .A1(N6524), .A2(n25743), .B1(N6491), .B2(n26394), .ZN(
        n4155) );
  OAI21_X1 U23362 ( .B1(n21058), .B2(n8158), .A(n4156), .ZN(n6125) );
  AOI22_X1 U23363 ( .A1(N6523), .A2(n24069), .B1(N6490), .B2(n25222), .ZN(
        n4156) );
  OAI21_X1 U23364 ( .B1(n24007), .B2(n8163), .A(n4157), .ZN(n6126) );
  AOI22_X1 U23365 ( .A1(N6522), .A2(n20800), .B1(N6489), .B2(n21961), .ZN(
        n4157) );
  OAI21_X1 U23366 ( .B1(n26633), .B2(n8168), .A(n4158), .ZN(n6127) );
  AOI22_X1 U23367 ( .A1(N6521), .A2(n25113), .B1(N6488), .B2(n20572), .ZN(
        n4158) );
  OAI21_X1 U23368 ( .B1(n25017), .B2(n8173), .A(n4159), .ZN(n6128) );
  AOI22_X1 U23369 ( .A1(N6520), .A2(n25006), .B1(N6487), .B2(n25221), .ZN(
        n4159) );
  OAI21_X1 U23370 ( .B1(n25244), .B2(n8178), .A(n4160), .ZN(n6129) );
  AOI22_X1 U23371 ( .A1(N6519), .A2(n22730), .B1(N6486), .B2(n25205), .ZN(
        n4160) );
  OAI21_X1 U23372 ( .B1(n24007), .B2(n8182), .A(n4161), .ZN(n6130) );
  AOI22_X1 U23373 ( .A1(N6518), .A2(n25753), .B1(N6485), .B2(n25221), .ZN(
        n4161) );
  OAI21_X1 U23374 ( .B1(n23999), .B2(n8647), .A(n3989), .ZN(n6011) );
  AOI22_X1 U23375 ( .A1(N5939), .A2(n26650), .B1(N5906), .B2(n20866), .ZN(
        n3989) );
  OAI21_X1 U23376 ( .B1(n25243), .B2(n8652), .A(n3990), .ZN(n6012) );
  AOI22_X1 U23377 ( .A1(N5938), .A2(n20796), .B1(N5905), .B2(n25068), .ZN(
        n3990) );
  OAI21_X1 U23378 ( .B1(n26922), .B2(n8657), .A(n3991), .ZN(n6013) );
  AOI22_X1 U23379 ( .A1(N5937), .A2(n25750), .B1(N5904), .B2(n21965), .ZN(
        n3991) );
  OAI21_X1 U23380 ( .B1(n24014), .B2(n8662), .A(n3992), .ZN(n60140) );
  AOI22_X1 U23381 ( .A1(N5936), .A2(n24075), .B1(N5903), .B2(n20872), .ZN(
        n3992) );
  OAI21_X1 U23382 ( .B1(n24006), .B2(n8667), .A(n3993), .ZN(n60150) );
  AOI22_X1 U23383 ( .A1(N5935), .A2(n24735), .B1(N5902), .B2(n26388), .ZN(
        n3993) );
  OAI21_X1 U23384 ( .B1(n25017), .B2(n8672), .A(n3994), .ZN(n60160) );
  AOI22_X1 U23385 ( .A1(N5934), .A2(n25114), .B1(N5901), .B2(n26392), .ZN(
        n3994) );
  OAI21_X1 U23386 ( .B1(n25016), .B2(n8677), .A(n3995), .ZN(n60170) );
  AOI22_X1 U23387 ( .A1(N5933), .A2(n24066), .B1(N5900), .B2(n20866), .ZN(
        n3995) );
  OAI21_X1 U23388 ( .B1(n24011), .B2(n8682), .A(n3996), .ZN(n60180) );
  AOI22_X1 U23389 ( .A1(N5932), .A2(n19032), .B1(N5899), .B2(n26393), .ZN(
        n3996) );
  OAI21_X1 U23390 ( .B1(n24002), .B2(n8687), .A(n3997), .ZN(n60190) );
  AOI22_X1 U23391 ( .A1(N5931), .A2(n19244), .B1(N5898), .B2(n24774), .ZN(
        n3997) );
  OAI21_X1 U23392 ( .B1(n25363), .B2(n8692), .A(n3998), .ZN(n60200) );
  AOI22_X1 U23393 ( .A1(N5930), .A2(n24079), .B1(N5897), .B2(n20575), .ZN(
        n3998) );
  OAI21_X1 U23394 ( .B1(n24417), .B2(n8697), .A(n3999), .ZN(n60210) );
  AOI22_X1 U23395 ( .A1(N5929), .A2(n25113), .B1(N5896), .B2(n25215), .ZN(
        n3999) );
  OAI21_X1 U23396 ( .B1(n26635), .B2(n8702), .A(n4000), .ZN(n60220) );
  AOI22_X1 U23397 ( .A1(N5928), .A2(n24999), .B1(N5895), .B2(n25216), .ZN(
        n4000) );
  OAI21_X1 U23398 ( .B1(n23999), .B2(n8707), .A(n4001), .ZN(n60230) );
  AOI22_X1 U23399 ( .A1(N5927), .A2(n24070), .B1(N5894), .B2(n21966), .ZN(
        n4001) );
  OAI21_X1 U23400 ( .B1(n25244), .B2(n8712), .A(n4002), .ZN(n60240) );
  AOI22_X1 U23401 ( .A1(N5926), .A2(n20523), .B1(N5893), .B2(n25206), .ZN(
        n4002) );
  OAI21_X1 U23402 ( .B1(n24417), .B2(n8716), .A(n4003), .ZN(n60250) );
  AOI22_X1 U23403 ( .A1(N5925), .A2(n21412), .B1(N5892), .B2(n25205), .ZN(
        n4003) );
  OAI21_X1 U23404 ( .B1(n23989), .B2(n9795), .A(n3648), .ZN(n5786) );
  AOI22_X1 U23405 ( .A1(N4660), .A2(n20518), .B1(N4627), .B2(n25072), .ZN(
        n3648) );
  OAI21_X1 U23406 ( .B1(n23997), .B2(n9800), .A(n3649), .ZN(n5787) );
  AOI22_X1 U23407 ( .A1(N4659), .A2(n22715), .B1(N4626), .B2(n20871), .ZN(
        n3649) );
  OAI21_X1 U23408 ( .B1(n22682), .B2(n9805), .A(n3650), .ZN(n5788) );
  AOI22_X1 U23409 ( .A1(N4658), .A2(n25008), .B1(N4625), .B2(n20876), .ZN(
        n3650) );
  OAI21_X1 U23410 ( .B1(n25246), .B2(n9810), .A(n3651), .ZN(n5789) );
  AOI22_X1 U23411 ( .A1(N4657), .A2(n22714), .B1(N4624), .B2(n26391), .ZN(
        n3651) );
  OAI21_X1 U23412 ( .B1(n23987), .B2(n9815), .A(n3652), .ZN(n5790) );
  AOI22_X1 U23413 ( .A1(N4656), .A2(n20805), .B1(N4623), .B2(n25202), .ZN(
        n3652) );
  OAI21_X1 U23414 ( .B1(n23994), .B2(n9820), .A(n3653), .ZN(n5791) );
  AOI22_X1 U23415 ( .A1(N4655), .A2(n22721), .B1(N4622), .B2(n25078), .ZN(
        n3653) );
  OAI21_X1 U23416 ( .B1(n26625), .B2(n9825), .A(n3654), .ZN(n5792) );
  AOI22_X1 U23417 ( .A1(N4654), .A2(n25111), .B1(N4621), .B2(n26382), .ZN(
        n3654) );
  OAI21_X1 U23418 ( .B1(n19103), .B2(n9830), .A(n3655), .ZN(n5793) );
  AOI22_X1 U23419 ( .A1(N4653), .A2(n27261), .B1(N4620), .B2(n21955), .ZN(
        n3655) );
  OAI21_X1 U23420 ( .B1(n19275), .B2(n9835), .A(n3656), .ZN(n5794) );
  AOI22_X1 U23421 ( .A1(N4652), .A2(n24056), .B1(N4619), .B2(n25212), .ZN(
        n3656) );
  OAI21_X1 U23422 ( .B1(n26630), .B2(n9840), .A(n3657), .ZN(n5795) );
  AOI22_X1 U23423 ( .A1(N4651), .A2(n22946), .B1(N4618), .B2(n20571), .ZN(
        n3657) );
  OAI21_X1 U23424 ( .B1(n24422), .B2(n9845), .A(n3658), .ZN(n5796) );
  AOI22_X1 U23425 ( .A1(N4650), .A2(n25737), .B1(N4617), .B2(n25209), .ZN(
        n3658) );
  OAI21_X1 U23426 ( .B1(n25021), .B2(n9850), .A(n3659), .ZN(n5797) );
  AOI22_X1 U23427 ( .A1(N4649), .A2(n19286), .B1(N4616), .B2(n26391), .ZN(
        n3659) );
  OAI21_X1 U23428 ( .B1(n19275), .B2(n9855), .A(n3660), .ZN(n5798) );
  AOI22_X1 U23429 ( .A1(N4648), .A2(n25012), .B1(N4615), .B2(n25213), .ZN(
        n3660) );
  OAI21_X1 U23430 ( .B1(n26630), .B2(n9860), .A(n3661), .ZN(n5799) );
  AOI22_X1 U23431 ( .A1(N4647), .A2(n25738), .B1(N4614), .B2(n20870), .ZN(
        n3661) );
  OAI21_X1 U23432 ( .B1(n25246), .B2(n9864), .A(n3662), .ZN(n5800) );
  AOI22_X1 U23433 ( .A1(N4646), .A2(n19285), .B1(N4613), .B2(n26383), .ZN(
        n3662) );
  OAI21_X1 U23434 ( .B1(n22682), .B2(n10329), .A(n3491), .ZN(n56810) );
  AOI22_X1 U23435 ( .A1(N4053), .A2(n19027), .B1(N4020), .B2(n21956), .ZN(
        n3491) );
  OAI21_X1 U23436 ( .B1(n23989), .B2(n10334), .A(n3492), .ZN(n56820) );
  AOI22_X1 U23437 ( .A1(N4052), .A2(n24065), .B1(N4019), .B2(n20877), .ZN(
        n3492) );
  OAI21_X1 U23438 ( .B1(n23998), .B2(n10339), .A(n3493), .ZN(n56830) );
  AOI22_X1 U23439 ( .A1(N4051), .A2(n257401), .B1(N4018), .B2(n25213), .ZN(
        n3493) );
  OAI21_X1 U23440 ( .B1(n25367), .B2(n10344), .A(n3494), .ZN(n56840) );
  AOI22_X1 U23441 ( .A1(N4050), .A2(n19031), .B1(N4017), .B2(n21949), .ZN(
        n3494) );
  OAI21_X1 U23442 ( .B1(n26925), .B2(n10349), .A(n3495), .ZN(n56850) );
  AOI22_X1 U23443 ( .A1(N4049), .A2(n24060), .B1(N4016), .B2(n26390), .ZN(
        n3495) );
  OAI21_X1 U23444 ( .B1(n23986), .B2(n10354), .A(n3496), .ZN(n56860) );
  AOI22_X1 U23445 ( .A1(N4048), .A2(n25103), .B1(N4015), .B2(n20570), .ZN(
        n3496) );
  OAI21_X1 U23446 ( .B1(n23995), .B2(n10359), .A(n3497), .ZN(n56870) );
  AOI22_X1 U23447 ( .A1(N4047), .A2(n25111), .B1(N4014), .B2(n20567), .ZN(
        n3497) );
  OAI21_X1 U23448 ( .B1(n24422), .B2(n10364), .A(n3498), .ZN(n56880) );
  AOI22_X1 U23449 ( .A1(N4046), .A2(n25010), .B1(N4013), .B2(n25212), .ZN(
        n3498) );
  OAI21_X1 U23450 ( .B1(n25022), .B2(n10369), .A(n34990), .ZN(n56890) );
  AOI22_X1 U23451 ( .A1(N4045), .A2(n25110), .B1(N4012), .B2(n21955), .ZN(
        n34990) );
  OAI21_X1 U23452 ( .B1(n26628), .B2(n10374), .A(n35000), .ZN(n56900) );
  AOI22_X1 U23453 ( .A1(N4044), .A2(n24733), .B1(N4011), .B2(n20568), .ZN(
        n35000) );
  OAI21_X1 U23454 ( .B1(n19276), .B2(n10379), .A(n35010), .ZN(n56910) );
  AOI22_X1 U23455 ( .A1(N4043), .A2(n20803), .B1(N4010), .B2(n20870), .ZN(
        n35010) );
  OAI21_X1 U23456 ( .B1(n26627), .B2(n10384), .A(n35020), .ZN(n56920) );
  AOI22_X1 U23457 ( .A1(N4042), .A2(n26648), .B1(N4009), .B2(n21950), .ZN(
        n35020) );
  OAI21_X1 U23458 ( .B1(n17123), .B2(n10389), .A(n35030), .ZN(n56930) );
  AOI22_X1 U23459 ( .A1(N4041), .A2(n25104), .B1(N4008), .B2(n24769), .ZN(
        n35030) );
  OAI21_X1 U23460 ( .B1(n26628), .B2(n10394), .A(n35040), .ZN(n56940) );
  AOI22_X1 U23461 ( .A1(N4040), .A2(n26649), .B1(N4007), .B2(n21951), .ZN(
        n35040) );
  OAI21_X1 U23462 ( .B1(n19276), .B2(n10398), .A(n35050), .ZN(n56950) );
  AOI22_X1 U23463 ( .A1(N4039), .A2(n19284), .B1(N4006), .B2(n25209), .ZN(
        n35050) );
  OAI21_X1 U23464 ( .B1(n24421), .B2(n10897), .A(n33310), .ZN(n5576) );
  AOI22_X1 U23465 ( .A1(N3467), .A2(n24056), .B1(N3434), .B2(n21949), .ZN(
        n33310) );
  OAI21_X1 U23466 ( .B1(n21065), .B2(n10901), .A(n33320), .ZN(n5577) );
  AOI22_X1 U23467 ( .A1(N3466), .A2(n24060), .B1(N3433), .B2(n21957), .ZN(
        n33320) );
  OAI21_X1 U23468 ( .B1(n23990), .B2(n10905), .A(n33330), .ZN(n5578) );
  AOI22_X1 U23469 ( .A1(N3465), .A2(n25741), .B1(N3432), .B2(n25208), .ZN(
        n33330) );
  OAI21_X1 U23470 ( .B1(n23997), .B2(n10909), .A(n33340), .ZN(n5579) );
  AOI22_X1 U23471 ( .A1(N3464), .A2(n24061), .B1(N3431), .B2(n25201), .ZN(
        n33340) );
  OAI21_X1 U23472 ( .B1(n26926), .B2(n10913), .A(n33350), .ZN(n5580) );
  AOI22_X1 U23473 ( .A1(N3463), .A2(n25012), .B1(N3430), .B2(n25203), .ZN(
        n33350) );
  OAI21_X1 U23474 ( .B1(n26926), .B2(n10917), .A(n33360), .ZN(n5581) );
  AOI22_X1 U23475 ( .A1(N3462), .A2(n25736), .B1(N3429), .B2(n26389), .ZN(
        n33360) );
  OAI21_X1 U23476 ( .B1(n23987), .B2(n10921), .A(n33370), .ZN(n5582) );
  AOI22_X1 U23477 ( .A1(N3461), .A2(n20921), .B1(N3428), .B2(n25199), .ZN(
        n33370) );
  OAI21_X1 U23478 ( .B1(n23994), .B2(n10925), .A(n33380), .ZN(n5583) );
  AOI22_X1 U23479 ( .A1(N3460), .A2(n20804), .B1(N3427), .B2(n25210), .ZN(
        n33380) );
  OAI21_X1 U23480 ( .B1(n19066), .B2(n10929), .A(n33390), .ZN(n5584) );
  AOI22_X1 U23481 ( .A1(N3459), .A2(n20808), .B1(N3426), .B2(n21951), .ZN(
        n33390) );
  OAI21_X1 U23482 ( .B1(n26627), .B2(n10933), .A(n33400), .ZN(n5585) );
  AOI22_X1 U23483 ( .A1(N3458), .A2(n24065), .B1(N3425), .B2(n25198), .ZN(
        n33400) );
  OAI21_X1 U23484 ( .B1(n26629), .B2(n10937), .A(n33410), .ZN(n55860) );
  AOI22_X1 U23485 ( .A1(N3457), .A2(n20806), .B1(N3424), .B2(n26383), .ZN(
        n33410) );
  OAI21_X1 U23486 ( .B1(n23991), .B2(n10941), .A(n33420), .ZN(n55870) );
  AOI22_X1 U23487 ( .A1(N3456), .A2(n25104), .B1(N3423), .B2(n25078), .ZN(
        n33420) );
  OAI21_X1 U23488 ( .B1(n19103), .B2(n10945), .A(n33430), .ZN(n55880) );
  AOI22_X1 U23489 ( .A1(N3455), .A2(n26647), .B1(N3422), .B2(n20567), .ZN(
        n33430) );
  OAI21_X1 U23490 ( .B1(n25021), .B2(n10949), .A(n33440), .ZN(n55890) );
  AOI22_X1 U23491 ( .A1(N3454), .A2(n22718), .B1(N3421), .B2(n24766), .ZN(
        n33440) );
  OAI21_X1 U23492 ( .B1(n23983), .B2(n10954), .A(n33450), .ZN(n55900) );
  AOI22_X1 U23493 ( .A1(N3453), .A2(n26647), .B1(N3420), .B2(n25200), .ZN(
        n33450) );
  OAI21_X1 U23494 ( .B1(n23991), .B2(n11419), .A(n3162), .ZN(n5471) );
  AOI22_X1 U23495 ( .A1(N2862), .A2(n22720), .B1(N2829), .B2(n25200), .ZN(
        n3162) );
  OAI21_X1 U23496 ( .B1(n25019), .B2(n11424), .A(n31630), .ZN(n5472) );
  AOI22_X1 U23497 ( .A1(N2861), .A2(n21406), .B1(N2828), .B2(n25199), .ZN(
        n31630) );
  OAI21_X1 U23498 ( .B1(n26924), .B2(n11429), .A(n31640), .ZN(n5473) );
  AOI22_X1 U23499 ( .A1(N2860), .A2(n20519), .B1(N2827), .B2(n21957), .ZN(
        n31640) );
  OAI21_X1 U23500 ( .B1(n23990), .B2(n11434), .A(n31650), .ZN(n54740) );
  AOI22_X1 U23501 ( .A1(N2859), .A2(n22717), .B1(N2826), .B2(n25072), .ZN(
        n31650) );
  OAI21_X1 U23502 ( .B1(n23998), .B2(n11439), .A(n31660), .ZN(n54750) );
  AOI22_X1 U23503 ( .A1(N2858), .A2(n20807), .B1(N2825), .B2(n24769), .ZN(
        n31660) );
  OAI21_X1 U23504 ( .B1(n22683), .B2(n11444), .A(n31670), .ZN(n54760) );
  AOI22_X1 U23505 ( .A1(N2857), .A2(n26646), .B1(N2824), .B2(n21952), .ZN(
        n31670) );
  OAI21_X1 U23506 ( .B1(n19066), .B2(n11449), .A(n31680), .ZN(n54770) );
  AOI22_X1 U23507 ( .A1(N2856), .A2(n24061), .B1(N2823), .B2(n24766), .ZN(
        n31680) );
  OAI21_X1 U23508 ( .B1(n23986), .B2(n11454), .A(n31690), .ZN(n54780) );
  AOI22_X1 U23509 ( .A1(N2855), .A2(n25741), .B1(N2822), .B2(n26381), .ZN(
        n31690) );
  OAI21_X1 U23510 ( .B1(n23995), .B2(n11459), .A(n31700), .ZN(n54790) );
  AOI22_X1 U23511 ( .A1(N2854), .A2(n25110), .B1(N2821), .B2(n25210), .ZN(
        n31700) );
  OAI21_X1 U23512 ( .B1(n25018), .B2(n11464), .A(n31710), .ZN(n54800) );
  AOI22_X1 U23513 ( .A1(N2853), .A2(n24059), .B1(N2820), .B2(n20570), .ZN(
        n31710) );
  OAI21_X1 U23514 ( .B1(n25367), .B2(n11469), .A(n31720), .ZN(n54810) );
  AOI22_X1 U23515 ( .A1(N2852), .A2(n25739), .B1(N2819), .B2(n25203), .ZN(
        n31720) );
  OAI21_X1 U23516 ( .B1(n23983), .B2(n11474), .A(n31730), .ZN(n54820) );
  AOI22_X1 U23517 ( .A1(N2851), .A2(n25109), .B1(N2818), .B2(n25211), .ZN(
        n31730) );
  OAI21_X1 U23518 ( .B1(n26631), .B2(n11479), .A(n31740), .ZN(n54830) );
  AOI22_X1 U23519 ( .A1(N2850), .A2(n24064), .B1(N2817), .B2(n21958), .ZN(
        n31740) );
  OAI21_X1 U23520 ( .B1(n25018), .B2(n11484), .A(n31750), .ZN(n54840) );
  AOI22_X1 U23521 ( .A1(N2849), .A2(n22945), .B1(N2816), .B2(n25202), .ZN(
        n31750) );
  OAI21_X1 U23522 ( .B1(n26625), .B2(n11488), .A(n31760), .ZN(n54850) );
  AOI22_X1 U23523 ( .A1(N2848), .A2(n25108), .B1(N2815), .B2(n20876), .ZN(
        n31760) );
  NAND3_X1 U23524 ( .A1(n50930), .A2(n50940), .A3(n50950), .ZN(mul_outcome[18]) );
  AOI22_X1 U23525 ( .A1(n26981), .A2(n17911), .B1(n25328), .B2(n17971), .ZN(
        n50930) );
  AOI22_X1 U23526 ( .A1(n21870), .A2(n17983), .B1(n25320), .B2(n17959), .ZN(
        n50940) );
  AOI221_X1 U23527 ( .B1(n17127), .B2(n17935), .C1(n17947), .C2(n25311), .A(
        n27785), .ZN(n50950) );
  NAND3_X1 U23528 ( .A1(n53110), .A2(n53120), .A3(n53130), .ZN(
        mul_outcome[123]) );
  AOI221_X1 U23529 ( .B1(n21972), .B2(n17479), .C1(n21437), .C2(n17467), .A(
        n27776), .ZN(n53130) );
  AOI22_X1 U23530 ( .A1(n27019), .A2(n17551), .B1(n27027), .B2(n17539), .ZN(
        n53120) );
  AOI22_X1 U23531 ( .A1(n27005), .A2(n17527), .B1(n19247), .B2(n17515), .ZN(
        n53110) );
  NAND3_X1 U23532 ( .A1(n4895), .A2(n4896), .A3(n4897), .ZN(mul_outcome[60])
         );
  AOI22_X1 U23533 ( .A1(n27052), .A2(n17815), .B1(n21340), .B2(n17803), .ZN(
        n4895) );
  AOI22_X1 U23534 ( .A1(n27066), .A2(n17839), .B1(n27079), .B2(n17827), .ZN(
        n4896) );
  AOI221_X1 U23535 ( .B1(n27090), .B2(n17791), .C1(n21358), .C2(n17779), .A(
        n27745), .ZN(n4897) );
  NAND2_X1 U23536 ( .A1(n4980), .A2(n4981), .ZN(mul_outcome[41]) );
  AOI221_X1 U23537 ( .B1(n21895), .B2(n17859), .C1(n26074), .C2(n17847), .A(
        n4988), .ZN(n4980) );
  AOI221_X1 U23538 ( .B1(n21880), .B2(n17883), .C1(n21885), .C2(n17871), .A(
        n4984), .ZN(n4981) );
  OAI22_X1 U23539 ( .A1(n2064), .A2(n19208), .B1(n2043), .B2(n19198), .ZN(
        n4988) );
  NAND3_X1 U23540 ( .A1(n5101), .A2(n5102), .A3(n5103), .ZN(mul_outcome[16])
         );
  AOI22_X1 U23541 ( .A1(n26979), .A2(n17915), .B1(n24155), .B2(n17975), .ZN(
        n5101) );
  AOI22_X1 U23542 ( .A1(n17118), .A2(n17987), .B1(n19084), .B2(n17963), .ZN(
        n5102) );
  AOI221_X1 U23543 ( .B1(n25939), .B2(n17939), .C1(n17951), .C2(n25309), .A(
        n27787), .ZN(n5103) );
  NAND3_X1 U23544 ( .A1(n53190), .A2(n53200), .A3(n53210), .ZN(
        mul_outcome[121]) );
  AOI221_X1 U23545 ( .B1(n24402), .B2(n17483), .C1(n21503), .C2(n17471), .A(
        n27778), .ZN(n53210) );
  AOI22_X1 U23546 ( .A1(n27017), .A2(n17555), .B1(n25184), .B2(n17543), .ZN(
        n53200) );
  AOI22_X1 U23547 ( .A1(n27003), .A2(n17531), .B1(n22827), .B2(n17519), .ZN(
        n53190) );
  NAND3_X1 U23548 ( .A1(n49070), .A2(n49080), .A3(n49090), .ZN(mul_outcome[58]) );
  AOI22_X1 U23549 ( .A1(n27050), .A2(n17819), .B1(n21342), .B2(n17807), .ZN(
        n49070) );
  AOI22_X1 U23550 ( .A1(n27064), .A2(n17843), .B1(n27077), .B2(n17831), .ZN(
        n49080) );
  AOI221_X1 U23551 ( .B1(n27088), .B2(n17795), .C1(n19231), .C2(n17783), .A(
        n27747), .ZN(n49090) );
  NAND3_X1 U23552 ( .A1(n53150), .A2(n53160), .A3(n53170), .ZN(
        mul_outcome[122]) );
  AOI221_X1 U23553 ( .B1(n26401), .B2(n17481), .C1(n22831), .C2(n17469), .A(
        n27777), .ZN(n53170) );
  AOI22_X1 U23554 ( .A1(n27018), .A2(n17553), .B1(n19052), .B2(n17541), .ZN(
        n53160) );
  AOI22_X1 U23555 ( .A1(n27004), .A2(n17529), .B1(n25917), .B2(n17517), .ZN(
        n53150) );
  NAND3_X1 U23556 ( .A1(n49030), .A2(n49040), .A3(n49050), .ZN(mul_outcome[59]) );
  AOI22_X1 U23557 ( .A1(n27051), .A2(n17817), .B1(n21333), .B2(n17805), .ZN(
        n49030) );
  AOI22_X1 U23558 ( .A1(n27065), .A2(n17841), .B1(n27078), .B2(n17829), .ZN(
        n49040) );
  AOI221_X1 U23559 ( .B1(n27089), .B2(n17793), .C1(n21350), .C2(n17781), .A(
        n27746), .ZN(n49050) );
  NAND3_X1 U23560 ( .A1(n53070), .A2(n53080), .A3(n53090), .ZN(
        mul_outcome[124]) );
  AOI221_X1 U23561 ( .B1(n23492), .B2(n17477), .C1(n26076), .C2(n17465), .A(
        n27775), .ZN(n53090) );
  AOI22_X1 U23562 ( .A1(n27020), .A2(n17549), .B1(n25183), .B2(n17537), .ZN(
        n53080) );
  AOI22_X1 U23563 ( .A1(n27006), .A2(n17525), .B1(n24259), .B2(n17513), .ZN(
        n53070) );
  NAND3_X1 U23564 ( .A1(n4891), .A2(n4892), .A3(n4893), .ZN(mul_outcome[61])
         );
  AOI22_X1 U23565 ( .A1(n27053), .A2(n17813), .B1(n21344), .B2(n17801), .ZN(
        n4891) );
  AOI22_X1 U23566 ( .A1(n27067), .A2(n17837), .B1(n27083), .B2(n17825), .ZN(
        n4892) );
  AOI221_X1 U23567 ( .B1(n27091), .B2(n17789), .C1(n21347), .C2(n17777), .A(
        n27744), .ZN(n4893) );
  NAND2_X1 U23568 ( .A1(n5203), .A2(n5204), .ZN(mul_outcome[146]) );
  AOI221_X1 U23569 ( .B1(n26902), .B2(n17391), .C1(n23378), .C2(n17367), .A(
        n27733), .ZN(n5203) );
  AOI221_X1 U23570 ( .B1(n19233), .B2(n17451), .C1(n27037), .C2(n17439), .A(
        n27749), .ZN(n5204) );
  INV_X1 U23571 ( .A(n5208), .ZN(n27733) );
  OAI21_X1 U23572 ( .B1(n22119), .B2(n11657), .A(n4572), .ZN(n6386) );
  NAND2_X1 U23573 ( .A1(n19368), .A2(n19079), .ZN(n4572) );
  OAI21_X1 U23574 ( .B1(n22089), .B2(n11660), .A(n4573), .ZN(n6387) );
  NAND2_X1 U23575 ( .A1(n19371), .A2(n22797), .ZN(n4573) );
  OAI21_X1 U23576 ( .B1(n22083), .B2(n11663), .A(n4574), .ZN(n6388) );
  NAND2_X1 U23577 ( .A1(n19374), .A2(n25283), .ZN(n4574) );
  OAI21_X1 U23578 ( .B1(n22053), .B2(n11666), .A(n4575), .ZN(n6389) );
  NAND2_X1 U23579 ( .A1(n19377), .A2(n25928), .ZN(n4575) );
  OAI21_X1 U23580 ( .B1(n22047), .B2(n11669), .A(n4576), .ZN(n6390) );
  NAND2_X1 U23581 ( .A1(n19380), .A2(n24921), .ZN(n4576) );
  OAI21_X1 U23582 ( .B1(n22017), .B2(n11672), .A(n4577), .ZN(n6391) );
  NAND2_X1 U23583 ( .A1(n19383), .A2(n22806), .ZN(n4577) );
  OAI21_X1 U23584 ( .B1(n22011), .B2(n11675), .A(n4578), .ZN(n6392) );
  NAND2_X1 U23585 ( .A1(n19386), .A2(n25629), .ZN(n4578) );
  OAI21_X1 U23586 ( .B1(n21981), .B2(n11678), .A(n4579), .ZN(n6393) );
  NAND2_X1 U23587 ( .A1(n19390), .A2(n25608), .ZN(n4579) );
  OAI21_X1 U23588 ( .B1(n22101), .B2(n11681), .A(n4580), .ZN(n6394) );
  NAND2_X1 U23589 ( .A1(n19392), .A2(n22792), .ZN(n4580) );
  OAI21_X1 U23590 ( .B1(n22095), .B2(n11684), .A(n4581), .ZN(n6395) );
  NAND2_X1 U23591 ( .A1(n19395), .A2(n25292), .ZN(n4581) );
  OAI21_X1 U23592 ( .B1(n22065), .B2(n11687), .A(n4582), .ZN(n63960) );
  NAND2_X1 U23593 ( .A1(n19398), .A2(n22806), .ZN(n4582) );
  OAI21_X1 U23594 ( .B1(n22059), .B2(n11690), .A(n4583), .ZN(n63970) );
  NAND2_X1 U23595 ( .A1(n19401), .A2(n24219), .ZN(n4583) );
  OAI21_X1 U23596 ( .B1(n22029), .B2(n11693), .A(n4584), .ZN(n63980) );
  NAND2_X1 U23597 ( .A1(n19404), .A2(n25319), .ZN(n4584) );
  OAI21_X1 U23598 ( .B1(n22023), .B2(n11696), .A(n4585), .ZN(n63990) );
  NAND2_X1 U23599 ( .A1(n19407), .A2(n25290), .ZN(n4585) );
  OAI21_X1 U23600 ( .B1(n21993), .B2(n11699), .A(n4586), .ZN(n64000) );
  NAND2_X1 U23601 ( .A1(n19410), .A2(n21014), .ZN(n4586) );
  OAI21_X1 U23602 ( .B1(n21987), .B2(n11702), .A(n4587), .ZN(n64010) );
  NAND2_X1 U23603 ( .A1(n19414), .A2(n19212), .ZN(n4587) );
  OAI21_X1 U23604 ( .B1(n22273), .B2(n11705), .A(n4588), .ZN(n64020) );
  NAND2_X1 U23605 ( .A1(n19416), .A2(n25316), .ZN(n4588) );
  OAI21_X1 U23606 ( .B1(n22256), .B2(n11708), .A(n4589), .ZN(n64030) );
  NAND2_X1 U23607 ( .A1(n19419), .A2(n26726), .ZN(n4589) );
  OAI21_X1 U23608 ( .B1(n22239), .B2(n11711), .A(n4590), .ZN(n64040) );
  NAND2_X1 U23609 ( .A1(n19422), .A2(n25282), .ZN(n4590) );
  OAI21_X1 U23610 ( .B1(n22221), .B2(n11714), .A(n4591), .ZN(n64050) );
  NAND2_X1 U23611 ( .A1(n19425), .A2(n25929), .ZN(n4591) );
  OAI21_X1 U23612 ( .B1(n22209), .B2(n11717), .A(n4592), .ZN(n64060) );
  NAND2_X1 U23613 ( .A1(n19428), .A2(n25287), .ZN(n4592) );
  OAI21_X1 U23614 ( .B1(n22169), .B2(n11720), .A(n4593), .ZN(n64070) );
  NAND2_X1 U23615 ( .A1(n19431), .A2(n19071), .ZN(n4593) );
  OAI21_X1 U23616 ( .B1(n22162), .B2(n11723), .A(n4594), .ZN(n64080) );
  NAND2_X1 U23617 ( .A1(n19434), .A2(n24221), .ZN(n4594) );
  OAI21_X1 U23618 ( .B1(n22125), .B2(n11726), .A(n4595), .ZN(n64090) );
  NAND2_X1 U23619 ( .A1(n19438), .A2(n25608), .ZN(n4595) );
  OAI21_X1 U23620 ( .B1(n23583), .B2(n11753), .A(n4604), .ZN(n6418) );
  NAND2_X1 U23621 ( .A1(n19464), .A2(n24922), .ZN(n4604) );
  OAI21_X1 U23622 ( .B1(n22251), .B2(n11756), .A(n4605), .ZN(n6419) );
  NAND2_X1 U23623 ( .A1(n19467), .A2(n19070), .ZN(n4605) );
  OAI21_X1 U23624 ( .B1(n22233), .B2(n11759), .A(n4606), .ZN(n6420) );
  NAND2_X1 U23625 ( .A1(n19470), .A2(n19225), .ZN(n4606) );
  OAI21_X1 U23626 ( .B1(n22215), .B2(n11762), .A(n4607), .ZN(n6421) );
  NAND2_X1 U23627 ( .A1(n19473), .A2(n25606), .ZN(n4607) );
  OAI21_X1 U23628 ( .B1(n22185), .B2(n11765), .A(n4608), .ZN(n6422) );
  NAND2_X1 U23629 ( .A1(n19476), .A2(n24921), .ZN(n4608) );
  OAI21_X1 U23630 ( .B1(n22176), .B2(n11768), .A(n4609), .ZN(n6423) );
  NAND2_X1 U23631 ( .A1(n19479), .A2(n25319), .ZN(n4609) );
  OAI21_X1 U23632 ( .B1(n22139), .B2(n11771), .A(n4610), .ZN(n6424) );
  NAND2_X1 U23633 ( .A1(n19482), .A2(n21014), .ZN(n4610) );
  OAI21_X1 U23634 ( .B1(n22132), .B2(n11774), .A(n4611), .ZN(n6425) );
  NAND2_X1 U23635 ( .A1(n19486), .A2(n22803), .ZN(n4611) );
  OAI21_X1 U23636 ( .B1(n21685), .B2(n11777), .A(n4612), .ZN(n6426) );
  NAND2_X1 U23637 ( .A1(n19488), .A2(n19080), .ZN(n4612) );
  OAI21_X1 U23638 ( .B1(n21673), .B2(n11780), .A(n46130), .ZN(n6427) );
  NAND2_X1 U23639 ( .A1(n19491), .A2(n25287), .ZN(n46130) );
  OAI21_X1 U23640 ( .B1(n21677), .B2(n11783), .A(n46140), .ZN(n6428) );
  NAND2_X1 U23641 ( .A1(n19494), .A2(n21323), .ZN(n46140) );
  OAI21_X1 U23642 ( .B1(n21665), .B2(n11786), .A(n46150), .ZN(n64290) );
  NAND2_X1 U23643 ( .A1(n19497), .A2(n259301), .ZN(n46150) );
  OAI21_X1 U23644 ( .B1(n21669), .B2(n11789), .A(n46160), .ZN(n64300) );
  NAND2_X1 U23645 ( .A1(n19500), .A2(n25317), .ZN(n46160) );
  OAI21_X1 U23646 ( .B1(n21657), .B2(n11792), .A(n46170), .ZN(n64310) );
  NAND2_X1 U23647 ( .A1(n19503), .A2(n22796), .ZN(n46170) );
  OAI21_X1 U23648 ( .B1(n21661), .B2(n11795), .A(n46180), .ZN(n64320) );
  NAND2_X1 U23649 ( .A1(n19506), .A2(n25284), .ZN(n46180) );
  OAI21_X1 U23650 ( .B1(n21649), .B2(n11798), .A(n46190), .ZN(n64330) );
  NAND2_X1 U23651 ( .A1(n19510), .A2(n24217), .ZN(n46190) );
  OAI21_X1 U23652 ( .B1(n24363), .B2(n11801), .A(n46200), .ZN(n64340) );
  NAND2_X1 U23653 ( .A1(n19512), .A2(n22791), .ZN(n46200) );
  OAI21_X1 U23654 ( .B1(n21705), .B2(n11804), .A(n46210), .ZN(n64350) );
  NAND2_X1 U23655 ( .A1(n19515), .A2(n25291), .ZN(n46210) );
  OAI21_X1 U23656 ( .B1(n21709), .B2(n11807), .A(n46220), .ZN(n64360) );
  NAND2_X1 U23657 ( .A1(n19518), .A2(n25284), .ZN(n46220) );
  OAI21_X1 U23658 ( .B1(n21697), .B2(n11810), .A(n46230), .ZN(n64370) );
  NAND2_X1 U23659 ( .A1(n19521), .A2(n24997), .ZN(n46230) );
  OAI21_X1 U23660 ( .B1(n21701), .B2(n11813), .A(n46240), .ZN(n64380) );
  NAND2_X1 U23661 ( .A1(n19524), .A2(n24923), .ZN(n46240) );
  OAI21_X1 U23662 ( .B1(n21689), .B2(n11816), .A(n46250), .ZN(n64390) );
  NAND2_X1 U23663 ( .A1(n19527), .A2(n20609), .ZN(n46250) );
  OAI21_X1 U23664 ( .B1(n21693), .B2(n11819), .A(n46260), .ZN(n64400) );
  NAND2_X1 U23665 ( .A1(n19530), .A2(n24220), .ZN(n46260) );
  OAI21_X1 U23666 ( .B1(n21681), .B2(n11822), .A(n46270), .ZN(n64410) );
  NAND2_X1 U23667 ( .A1(n19534), .A2(n19069), .ZN(n46270) );
  OAI21_X1 U23668 ( .B1(n22146), .B2(n14537), .A(n46990), .ZN(n7353) );
  NAND2_X1 U23669 ( .A1(n19584), .A2(n20794), .ZN(n46990) );
  OAI21_X1 U23670 ( .B1(n22155), .B2(n14540), .A(n46980), .ZN(n7352) );
  NAND2_X1 U23671 ( .A1(n19587), .A2(n22802), .ZN(n46980) );
  OAI21_X1 U23672 ( .B1(n22192), .B2(n14543), .A(n46970), .ZN(n7351) );
  NAND2_X1 U23673 ( .A1(n19590), .A2(n20610), .ZN(n46970) );
  OAI21_X1 U23674 ( .B1(n22200), .B2(n14546), .A(n46960), .ZN(n7350) );
  NAND2_X1 U23675 ( .A1(n19593), .A2(n25317), .ZN(n46960) );
  OAI21_X1 U23676 ( .B1(n22227), .B2(n14549), .A(n46950), .ZN(n7349) );
  NAND2_X1 U23677 ( .A1(n19596), .A2(n24217), .ZN(n46950) );
  OAI21_X1 U23678 ( .B1(n22245), .B2(n14552), .A(n4694), .ZN(n7348) );
  NAND2_X1 U23679 ( .A1(n19599), .A2(n24087), .ZN(n4694) );
  OAI21_X1 U23680 ( .B1(n22262), .B2(n14555), .A(n4693), .ZN(n7347) );
  NAND2_X1 U23681 ( .A1(n19602), .A2(n25286), .ZN(n4693) );
  OAI21_X1 U23682 ( .B1(n22281), .B2(n14558), .A(n4692), .ZN(n7346) );
  NAND2_X1 U23683 ( .A1(n19605), .A2(n25070), .ZN(n4692) );
  OAI21_X1 U23684 ( .B1(n21999), .B2(n14857), .A(n4691), .ZN(n7289) );
  NAND2_X1 U23685 ( .A1(n19608), .A2(n19069), .ZN(n4691) );
  OAI21_X1 U23686 ( .B1(n22005), .B2(n14860), .A(n4690), .ZN(n7288) );
  NAND2_X1 U23687 ( .A1(n19611), .A2(n21280), .ZN(n4690) );
  OAI21_X1 U23688 ( .B1(n22035), .B2(n14863), .A(n4689), .ZN(n7287) );
  NAND2_X1 U23689 ( .A1(n19614), .A2(n23717), .ZN(n4689) );
  OAI21_X1 U23690 ( .B1(n22041), .B2(n14866), .A(n4688), .ZN(n72860) );
  NAND2_X1 U23691 ( .A1(n19617), .A2(n24922), .ZN(n4688) );
  OAI21_X1 U23692 ( .B1(n22071), .B2(n14869), .A(n4687), .ZN(n72850) );
  NAND2_X1 U23693 ( .A1(n19620), .A2(n24085), .ZN(n4687) );
  OAI21_X1 U23694 ( .B1(n22077), .B2(n14872), .A(n4686), .ZN(n72840) );
  NAND2_X1 U23695 ( .A1(n19623), .A2(n21324), .ZN(n4686) );
  OAI21_X1 U23696 ( .B1(n22107), .B2(n14875), .A(n4685), .ZN(n72830) );
  NAND2_X1 U23697 ( .A1(n19626), .A2(n25288), .ZN(n4685) );
  OAI21_X1 U23698 ( .B1(n22113), .B2(n14878), .A(n4684), .ZN(n72820) );
  NAND2_X1 U23699 ( .A1(n19629), .A2(n24814), .ZN(n4684) );
  OAI21_X1 U23700 ( .B1(n22123), .B2(n15177), .A(n4683), .ZN(n72250) );
  NAND2_X1 U23701 ( .A1(n19632), .A2(n259301), .ZN(n4683) );
  OAI21_X1 U23702 ( .B1(n22160), .B2(n15180), .A(n4682), .ZN(n72240) );
  NAND2_X1 U23703 ( .A1(n19635), .A2(n24086), .ZN(n4682) );
  OAI21_X1 U23704 ( .B1(n22167), .B2(n15183), .A(n4681), .ZN(n72230) );
  NAND2_X1 U23705 ( .A1(n19638), .A2(n25070), .ZN(n4681) );
  OAI21_X1 U23706 ( .B1(n22206), .B2(n15186), .A(n4680), .ZN(n72220) );
  NAND2_X1 U23707 ( .A1(n19641), .A2(n19079), .ZN(n4680) );
  OAI21_X1 U23708 ( .B1(n22219), .B2(n15189), .A(n4679), .ZN(n7221) );
  NAND2_X1 U23709 ( .A1(n19644), .A2(n25283), .ZN(n4679) );
  OAI21_X1 U23710 ( .B1(n22237), .B2(n15192), .A(n4678), .ZN(n7220) );
  NAND2_X1 U23711 ( .A1(n19647), .A2(n24219), .ZN(n4678) );
  OAI21_X1 U23712 ( .B1(n22255), .B2(n15195), .A(n4677), .ZN(n7219) );
  NAND2_X1 U23713 ( .A1(n19650), .A2(n23721), .ZN(n4677) );
  OAI21_X1 U23714 ( .B1(n22270), .B2(n15198), .A(n4676), .ZN(n7218) );
  NAND2_X1 U23715 ( .A1(n19653), .A2(n24809), .ZN(n4676) );
  OAI21_X1 U23716 ( .B1(n22129), .B2(n15817), .A(n4667), .ZN(n70970) );
  NAND2_X1 U23717 ( .A1(n19680), .A2(n24084), .ZN(n4667) );
  OAI21_X1 U23718 ( .B1(n22137), .B2(n15820), .A(n46660), .ZN(n7096) );
  NAND2_X1 U23719 ( .A1(n19683), .A2(n24216), .ZN(n46660) );
  OAI21_X1 U23720 ( .B1(n22173), .B2(n15823), .A(n46650), .ZN(n7095) );
  NAND2_X1 U23721 ( .A1(n19686), .A2(n18853), .ZN(n46650) );
  OAI21_X1 U23722 ( .B1(n22182), .B2(n15826), .A(n46640), .ZN(n7094) );
  NAND2_X1 U23723 ( .A1(n19689), .A2(n23718), .ZN(n46640) );
  OAI21_X1 U23724 ( .B1(n22213), .B2(n15829), .A(n46630), .ZN(n7093) );
  NAND2_X1 U23725 ( .A1(n19692), .A2(n19225), .ZN(n46630) );
  OAI21_X1 U23726 ( .B1(n22231), .B2(n15832), .A(n46620), .ZN(n7092) );
  NAND2_X1 U23727 ( .A1(n19695), .A2(n24082), .ZN(n46620) );
  OAI21_X1 U23728 ( .B1(n22249), .B2(n15835), .A(n46610), .ZN(n7091) );
  NAND2_X1 U23729 ( .A1(n19698), .A2(n20868), .ZN(n46610) );
  OAI21_X1 U23730 ( .B1(n24369), .B2(n15838), .A(n46600), .ZN(n7090) );
  NAND2_X1 U23731 ( .A1(n19701), .A2(n26715), .ZN(n46600) );
  OAI21_X1 U23732 ( .B1(n21979), .B2(n16137), .A(n46590), .ZN(n7033) );
  NAND2_X1 U23733 ( .A1(n19704), .A2(n20795), .ZN(n46590) );
  OAI21_X1 U23734 ( .B1(n22009), .B2(n16140), .A(n46580), .ZN(n7032) );
  NAND2_X1 U23735 ( .A1(n19707), .A2(n24086), .ZN(n46580) );
  OAI21_X1 U23736 ( .B1(n22015), .B2(n16143), .A(n46570), .ZN(n7031) );
  NAND2_X1 U23737 ( .A1(n19710), .A2(n18852), .ZN(n46570) );
  OAI21_X1 U23738 ( .B1(n22045), .B2(n16146), .A(n46560), .ZN(n70300) );
  NAND2_X1 U23739 ( .A1(n19713), .A2(n26585), .ZN(n46560) );
  OAI21_X1 U23740 ( .B1(n22051), .B2(n16149), .A(n46550), .ZN(n70290) );
  NAND2_X1 U23741 ( .A1(n19716), .A2(n24084), .ZN(n46550) );
  OAI21_X1 U23742 ( .B1(n22081), .B2(n16152), .A(n46540), .ZN(n70280) );
  NAND2_X1 U23743 ( .A1(n19719), .A2(n21279), .ZN(n46540) );
  OAI21_X1 U23744 ( .B1(n22087), .B2(n16155), .A(n46530), .ZN(n70270) );
  NAND2_X1 U23745 ( .A1(n19722), .A2(n23720), .ZN(n46530) );
  OAI21_X1 U23746 ( .B1(n22117), .B2(n16158), .A(n46520), .ZN(n70260) );
  NAND2_X1 U23747 ( .A1(n19725), .A2(n19071), .ZN(n46520) );
  OAI21_X1 U23748 ( .B1(n21985), .B2(n16457), .A(n46510), .ZN(n69690) );
  NAND2_X1 U23749 ( .A1(n19728), .A2(n22805), .ZN(n46510) );
  OAI21_X1 U23750 ( .B1(n21991), .B2(n16460), .A(n46500), .ZN(n69680) );
  NAND2_X1 U23751 ( .A1(n19731), .A2(n25929), .ZN(n46500) );
  OAI21_X1 U23752 ( .B1(n22021), .B2(n16463), .A(n46490), .ZN(n69670) );
  NAND2_X1 U23753 ( .A1(n19734), .A2(n22793), .ZN(n46490) );
  OAI21_X1 U23754 ( .B1(n22027), .B2(n16466), .A(n46480), .ZN(n69660) );
  NAND2_X1 U23755 ( .A1(n19737), .A2(n24814), .ZN(n46480) );
  OAI21_X1 U23756 ( .B1(n22057), .B2(n16469), .A(n46470), .ZN(n69650) );
  NAND2_X1 U23757 ( .A1(n19740), .A2(n24083), .ZN(n46470) );
  OAI21_X1 U23758 ( .B1(n22063), .B2(n16472), .A(n46460), .ZN(n69640) );
  NAND2_X1 U23759 ( .A1(n19743), .A2(n21015), .ZN(n46460) );
  OAI21_X1 U23760 ( .B1(n22093), .B2(n16475), .A(n4645), .ZN(n69630) );
  NAND2_X1 U23761 ( .A1(n19746), .A2(n23717), .ZN(n4645) );
  OAI21_X1 U23762 ( .B1(n22099), .B2(n16478), .A(n4644), .ZN(n69620) );
  NAND2_X1 U23763 ( .A1(n19749), .A2(n19070), .ZN(n4644) );
  OAI21_X1 U23764 ( .B1(n21769), .B2(n11729), .A(n4596), .ZN(n64100) );
  NAND2_X1 U23765 ( .A1(n19440), .A2(n19080), .ZN(n4596) );
  OAI21_X1 U23766 ( .B1(n21761), .B2(n11732), .A(n4597), .ZN(n64110) );
  NAND2_X1 U23767 ( .A1(n19443), .A2(n23718), .ZN(n4597) );
  OAI21_X1 U23768 ( .B1(n21753), .B2(n11735), .A(n4598), .ZN(n6412) );
  NAND2_X1 U23769 ( .A1(n19446), .A2(n19212), .ZN(n4598) );
  OAI21_X1 U23770 ( .B1(n21745), .B2(n11738), .A(n4599), .ZN(n6413) );
  NAND2_X1 U23771 ( .A1(n19449), .A2(n24087), .ZN(n4599) );
  OAI21_X1 U23772 ( .B1(n21737), .B2(n11741), .A(n4600), .ZN(n6414) );
  NAND2_X1 U23773 ( .A1(n19452), .A2(n20869), .ZN(n4600) );
  OAI21_X1 U23774 ( .B1(n21729), .B2(n11744), .A(n4601), .ZN(n6415) );
  NAND2_X1 U23775 ( .A1(n19455), .A2(n26585), .ZN(n4601) );
  OAI21_X1 U23776 ( .B1(n21721), .B2(n11747), .A(n4602), .ZN(n6416) );
  NAND2_X1 U23777 ( .A1(n19458), .A2(n25629), .ZN(n4602) );
  OAI21_X1 U23778 ( .B1(n21713), .B2(n11750), .A(n4603), .ZN(n6417) );
  NAND2_X1 U23779 ( .A1(n19462), .A2(n25927), .ZN(n4603) );
  OAI21_X1 U23780 ( .B1(n21773), .B2(n11825), .A(n46280), .ZN(n64420) );
  NAND2_X1 U23781 ( .A1(n19536), .A2(n23720), .ZN(n46280) );
  OAI21_X1 U23782 ( .B1(n21765), .B2(n11828), .A(n4629), .ZN(n64430) );
  NAND2_X1 U23783 ( .A1(n19539), .A2(n24809), .ZN(n4629) );
  OAI21_X1 U23784 ( .B1(n21757), .B2(n11831), .A(n4630), .ZN(n64440) );
  NAND2_X1 U23785 ( .A1(n19542), .A2(n24085), .ZN(n4630) );
  OAI21_X1 U23786 ( .B1(n21749), .B2(n11834), .A(n4631), .ZN(n64450) );
  NAND2_X1 U23787 ( .A1(n19545), .A2(n25607), .ZN(n4631) );
  OAI21_X1 U23788 ( .B1(n21741), .B2(n11837), .A(n4632), .ZN(n64460) );
  NAND2_X1 U23789 ( .A1(n19548), .A2(n22531), .ZN(n4632) );
  OAI21_X1 U23790 ( .B1(n21733), .B2(n11840), .A(n4633), .ZN(n64470) );
  NAND2_X1 U23791 ( .A1(n19551), .A2(n25289), .ZN(n4633) );
  OAI21_X1 U23792 ( .B1(n21725), .B2(n11843), .A(n4634), .ZN(n64480) );
  NAND2_X1 U23793 ( .A1(n19554), .A2(n22801), .ZN(n4634) );
  OAI21_X1 U23794 ( .B1(n21717), .B2(n11846), .A(n4635), .ZN(n64490) );
  NAND2_X1 U23795 ( .A1(n19558), .A2(n24082), .ZN(n4635) );
  OAI21_X1 U23796 ( .B1(n22417), .B2(n14217), .A(n4636), .ZN(n6898) );
  NAND2_X1 U23797 ( .A1(n19560), .A2(n22790), .ZN(n4636) );
  OAI21_X1 U23798 ( .B1(n22405), .B2(n14220), .A(n4637), .ZN(n6899) );
  NAND2_X1 U23799 ( .A1(n19563), .A2(n20606), .ZN(n4637) );
  OAI21_X1 U23800 ( .B1(n22393), .B2(n14223), .A(n4638), .ZN(n6900) );
  NAND2_X1 U23801 ( .A1(n19566), .A2(n25928), .ZN(n4638) );
  OAI21_X1 U23802 ( .B1(n22381), .B2(n14226), .A(n4639), .ZN(n6901) );
  NAND2_X1 U23803 ( .A1(n19569), .A2(n22803), .ZN(n4639) );
  OAI21_X1 U23804 ( .B1(n22369), .B2(n14229), .A(n4640), .ZN(n6902) );
  NAND2_X1 U23805 ( .A1(n19572), .A2(n22530), .ZN(n4640) );
  OAI21_X1 U23806 ( .B1(n22357), .B2(n14232), .A(n4641), .ZN(n6903) );
  NAND2_X1 U23807 ( .A1(n19575), .A2(n25292), .ZN(n4641) );
  OAI21_X1 U23808 ( .B1(n22345), .B2(n14235), .A(n4642), .ZN(n6904) );
  NAND2_X1 U23809 ( .A1(n19578), .A2(n24083), .ZN(n4642) );
  OAI21_X1 U23810 ( .B1(n22333), .B2(n14238), .A(n4643), .ZN(n6905) );
  NAND2_X1 U23811 ( .A1(n19581), .A2(n24221), .ZN(n4643) );
  OAI21_X1 U23812 ( .B1(n22327), .B2(n15497), .A(n4675), .ZN(n7161) );
  NAND2_X1 U23813 ( .A1(n19656), .A2(n22805), .ZN(n4675) );
  OAI21_X1 U23814 ( .B1(n22339), .B2(n15500), .A(n4674), .ZN(n7160) );
  NAND2_X1 U23815 ( .A1(n19659), .A2(n24997), .ZN(n4674) );
  OAI21_X1 U23816 ( .B1(n22351), .B2(n15503), .A(n4673), .ZN(n7159) );
  NAND2_X1 U23817 ( .A1(n19662), .A2(n25318), .ZN(n4673) );
  OAI21_X1 U23818 ( .B1(n22363), .B2(n15506), .A(n4672), .ZN(n7158) );
  NAND2_X1 U23819 ( .A1(n19665), .A2(n25290), .ZN(n4672) );
  OAI21_X1 U23820 ( .B1(n22375), .B2(n15509), .A(n4671), .ZN(n7157) );
  NAND2_X1 U23821 ( .A1(n19668), .A2(n24218), .ZN(n4671) );
  OAI21_X1 U23822 ( .B1(n22387), .B2(n15512), .A(n4670), .ZN(n7156) );
  NAND2_X1 U23823 ( .A1(n19671), .A2(n25606), .ZN(n4670) );
  OAI21_X1 U23824 ( .B1(n22399), .B2(n15515), .A(n4669), .ZN(n7155) );
  NAND2_X1 U23825 ( .A1(n19674), .A2(n23721), .ZN(n4669) );
  OAI21_X1 U23826 ( .B1(n22411), .B2(n15518), .A(n4668), .ZN(n7154) );
  NAND2_X1 U23827 ( .A1(n19677), .A2(n20606), .ZN(n4668) );
  NAND2_X1 U23828 ( .A1(n49990), .A2(n50000), .ZN(mul_outcome[39]) );
  AOI221_X1 U23829 ( .B1(n21547), .B2(n17863), .C1(n26072), .C2(n17851), .A(
        n50020), .ZN(n49990) );
  AOI221_X1 U23830 ( .B1(n21551), .B2(n17887), .C1(n21538), .C2(n17875), .A(
        n50010), .ZN(n50000) );
  OAI22_X1 U23831 ( .A1(n2066), .A2(n21258), .B1(n2045), .B2(n21221), .ZN(
        n50020) );
  OAI21_X1 U23832 ( .B1(n26371), .B2(n32100), .A(n4407), .ZN(n6286) );
  AOI22_X1 U23833 ( .A1(N7481), .A2(n21482), .B1(N7448), .B2(n25900), .ZN(
        n4407) );
  OAI21_X1 U23834 ( .B1(n26360), .B2(n33010), .A(n4408), .ZN(n6287) );
  AOI22_X1 U23835 ( .A1(N7480), .A2(n21468), .B1(N7447), .B2(n25896), .ZN(
        n4408) );
  OAI21_X1 U23836 ( .B1(n26364), .B2(n38460), .A(n4409), .ZN(n6288) );
  AOI22_X1 U23837 ( .A1(N7479), .A2(n24256), .B1(N7446), .B2(n20585), .ZN(
        n4409) );
  OAI21_X1 U23838 ( .B1(n21920), .B2(n4568), .A(n4410), .ZN(n6289) );
  AOI22_X1 U23839 ( .A1(N7478), .A2(n21474), .B1(N7445), .B2(n21270), .ZN(
        n4410) );
  OAI21_X1 U23840 ( .B1(n26357), .B2(n47870), .A(n4411), .ZN(n6290) );
  AOI22_X1 U23841 ( .A1(N7477), .A2(n21837), .B1(N7444), .B2(n25588), .ZN(
        n4411) );
  OAI21_X1 U23842 ( .B1(n21940), .B2(n5107), .A(n4412), .ZN(n6291) );
  AOI22_X1 U23843 ( .A1(N7476), .A2(n26045), .B1(N7443), .B2(n21268), .ZN(
        n4412) );
  OAI21_X1 U23844 ( .B1(n21928), .B2(n5417), .A(n4413), .ZN(n6292) );
  AOI22_X1 U23845 ( .A1(N7475), .A2(n24247), .B1(N7442), .B2(n22887), .ZN(
        n4413) );
  OAI21_X1 U23846 ( .B1(n21932), .B2(n7414), .A(n4414), .ZN(n6293) );
  AOI22_X1 U23847 ( .A1(N7474), .A2(n22867), .B1(N7441), .B2(n25890), .ZN(
        n4414) );
  OAI21_X1 U23848 ( .B1(n21923), .B2(n7423), .A(n4416), .ZN(n6295) );
  AOI22_X1 U23849 ( .A1(N7472), .A2(n21461), .B1(N7439), .B2(n24793), .ZN(
        n4416) );
  OAI21_X1 U23850 ( .B1(n21943), .B2(n7805), .A(n4242), .ZN(n6176) );
  AOI22_X1 U23851 ( .A1(N6888), .A2(n21844), .B1(N6855), .B2(n25595), .ZN(
        n4242) );
  OAI21_X1 U23852 ( .B1(n21930), .B2(n78090), .A(n4243), .ZN(n6177) );
  AOI22_X1 U23853 ( .A1(N6887), .A2(n23168), .B1(N6854), .B2(n22885), .ZN(
        n4243) );
  OAI21_X1 U23854 ( .B1(n21935), .B2(n78130), .A(n4244), .ZN(n6178) );
  AOI22_X1 U23855 ( .A1(N6886), .A2(n19308), .B1(N6853), .B2(n20586), .ZN(
        n4244) );
  OAI21_X1 U23856 ( .B1(n26356), .B2(n78170), .A(n4245), .ZN(n6179) );
  AOI22_X1 U23857 ( .A1(N6885), .A2(n22876), .B1(N6852), .B2(n22884), .ZN(
        n4245) );
  OAI21_X1 U23858 ( .B1(n21925), .B2(n78210), .A(n4246), .ZN(n6180) );
  AOI22_X1 U23859 ( .A1(N6884), .A2(n26766), .B1(N6851), .B2(n20588), .ZN(
        n4246) );
  OAI21_X1 U23860 ( .B1(n26372), .B2(n78250), .A(n4247), .ZN(n6181) );
  AOI22_X1 U23861 ( .A1(N6883), .A2(n26006), .B1(N6850), .B2(n25586), .ZN(
        n4247) );
  OAI21_X1 U23862 ( .B1(n26362), .B2(n7829), .A(n4248), .ZN(n61820) );
  AOI22_X1 U23863 ( .A1(N6882), .A2(n24256), .B1(N6849), .B2(n24788), .ZN(
        n4248) );
  OAI21_X1 U23864 ( .B1(n26365), .B2(n7833), .A(n4249), .ZN(n61830) );
  AOI22_X1 U23865 ( .A1(N6881), .A2(n26314), .B1(N6848), .B2(n24791), .ZN(
        n4249) );
  OAI21_X1 U23866 ( .B1(n26354), .B2(n7837), .A(n4250), .ZN(n61840) );
  AOI22_X1 U23867 ( .A1(N6880), .A2(n24264), .B1(N6847), .B2(n24468), .ZN(
        n4250) );
  OAI21_X1 U23868 ( .B1(n26359), .B2(n7841), .A(n4251), .ZN(n61850) );
  AOI22_X1 U23869 ( .A1(N6879), .A2(n26042), .B1(N6846), .B2(n24465), .ZN(
        n4251) );
  OAI21_X1 U23870 ( .B1(n26348), .B2(n7978), .A(n4199), .ZN(n61510) );
  AOI22_X1 U23871 ( .A1(N6709), .A2(n26063), .B1(N6676), .B2(n25866), .ZN(
        n4199) );
  OAI21_X1 U23872 ( .B1(n26352), .B2(n79830), .A(n4200), .ZN(n61520) );
  AOI22_X1 U23873 ( .A1(N6708), .A2(n21472), .B1(N6675), .B2(n25876), .ZN(
        n4200) );
  OAI21_X1 U23874 ( .B1(n26342), .B2(n79880), .A(n4201), .ZN(n61530) );
  AOI22_X1 U23875 ( .A1(N6707), .A2(n23164), .B1(N6674), .B2(n24492), .ZN(
        n4201) );
  OAI21_X1 U23876 ( .B1(n26347), .B2(n79930), .A(n4202), .ZN(n61540) );
  AOI22_X1 U23877 ( .A1(N6706), .A2(n21479), .B1(N6673), .B2(n24495), .ZN(
        n4202) );
  OAI21_X1 U23878 ( .B1(n26336), .B2(n79980), .A(n4203), .ZN(n61550) );
  AOI22_X1 U23879 ( .A1(N6705), .A2(n21841), .B1(N6672), .B2(n22893), .ZN(
        n4203) );
  OAI21_X1 U23880 ( .B1(n21908), .B2(n8003), .A(n4204), .ZN(n61560) );
  AOI22_X1 U23881 ( .A1(N6704), .A2(n23204), .B1(N6671), .B2(n25576), .ZN(
        n4204) );
  OAI21_X1 U23882 ( .B1(n21912), .B2(n8008), .A(n4205), .ZN(n61570) );
  AOI22_X1 U23883 ( .A1(N6703), .A2(n24240), .B1(N6670), .B2(n20548), .ZN(
        n4205) );
  OAI21_X1 U23884 ( .B1(n21898), .B2(n8013), .A(n4206), .ZN(n61580) );
  AOI22_X1 U23885 ( .A1(N6702), .A2(n26774), .B1(N6669), .B2(n25863), .ZN(
        n4206) );
  OAI21_X1 U23886 ( .B1(n21888), .B2(n8022), .A(n42080), .ZN(n61600) );
  AOI22_X1 U23887 ( .A1(N6700), .A2(n26011), .B1(N6667), .B2(n24487), .ZN(
        n42080) );
  OAI21_X1 U23888 ( .B1(n263701), .B2(n8327), .A(n4081), .ZN(n60710) );
  AOI22_X1 U23889 ( .A1(N6275), .A2(n260201), .B1(N6242), .B2(n25885), .ZN(
        n4081) );
  OAI21_X1 U23890 ( .B1(n26361), .B2(n8332), .A(n4082), .ZN(n60720) );
  AOI22_X1 U23891 ( .A1(N6274), .A2(n26044), .B1(N6241), .B2(n21430), .ZN(
        n4082) );
  OAI21_X1 U23892 ( .B1(n26363), .B2(n8337), .A(n4083), .ZN(n60730) );
  AOI22_X1 U23893 ( .A1(N6273), .A2(n21835), .B1(N6240), .B2(n21431), .ZN(
        n4083) );
  OAI21_X1 U23894 ( .B1(n21918), .B2(n8342), .A(n4084), .ZN(n60740) );
  AOI22_X1 U23895 ( .A1(N6272), .A2(n22842), .B1(N6239), .B2(n24468), .ZN(
        n4084) );
  OAI21_X1 U23896 ( .B1(n26358), .B2(n8347), .A(n4085), .ZN(n60750) );
  AOI22_X1 U23897 ( .A1(N6271), .A2(n19310), .B1(N6238), .B2(n25901), .ZN(
        n4085) );
  OAI21_X1 U23898 ( .B1(n21910), .B2(n8487), .A(n4037), .ZN(n6041) );
  AOI22_X1 U23899 ( .A1(N6107), .A2(n21852), .B1(N6074), .B2(n21253), .ZN(
        n4037) );
  OAI21_X1 U23900 ( .B1(n21915), .B2(n8492), .A(n4038), .ZN(n6042) );
  AOI22_X1 U23901 ( .A1(N6106), .A2(n22844), .B1(N6073), .B2(n24493), .ZN(
        n4038) );
  OAI21_X1 U23902 ( .B1(n21900), .B2(n8497), .A(n40390), .ZN(n6043) );
  AOI22_X1 U23903 ( .A1(N6105), .A2(n22832), .B1(N6072), .B2(n24495), .ZN(
        n40390) );
  OAI21_X1 U23904 ( .B1(n26345), .B2(n8502), .A(n40400), .ZN(n6044) );
  AOI22_X1 U23905 ( .A1(N6104), .A2(n26777), .B1(N6071), .B2(n21255), .ZN(
        n40400) );
  OAI21_X1 U23906 ( .B1(n21890), .B2(n8507), .A(n40410), .ZN(n6045) );
  AOI22_X1 U23907 ( .A1(N6103), .A2(n21498), .B1(N6070), .B2(n25576), .ZN(
        n40410) );
  OAI21_X1 U23908 ( .B1(n26350), .B2(n8512), .A(n40420), .ZN(n6046) );
  AOI22_X1 U23909 ( .A1(N6102), .A2(n26016), .B1(N6069), .B2(n24752), .ZN(
        n40420) );
  OAI21_X1 U23910 ( .B1(n26353), .B2(n8517), .A(n40430), .ZN(n6047) );
  AOI22_X1 U23911 ( .A1(N6101), .A2(n22859), .B1(N6068), .B2(n22890), .ZN(
        n40430) );
  OAI21_X1 U23912 ( .B1(n26344), .B2(n8522), .A(n40440), .ZN(n6048) );
  AOI22_X1 U23913 ( .A1(N6100), .A2(n21856), .B1(N6067), .B2(n24754), .ZN(
        n40440) );
  OAI21_X1 U23914 ( .B1(n21903), .B2(n8527), .A(n40450), .ZN(n6049) );
  AOI22_X1 U23915 ( .A1(N6099), .A2(n22861), .B1(N6066), .B2(n24489), .ZN(
        n40450) );
  OAI21_X1 U23916 ( .B1(n26338), .B2(n8532), .A(n40460), .ZN(n6050) );
  AOI22_X1 U23917 ( .A1(N6098), .A2(n26062), .B1(N6065), .B2(n24491), .ZN(
        n40460) );
  OAI21_X1 U23918 ( .B1(n21941), .B2(n8913), .A(n39300), .ZN(n5976) );
  AOI22_X1 U23919 ( .A1(N5679), .A2(n26772), .B1(N5646), .B2(n24466), .ZN(
        n39300) );
  OAI21_X1 U23920 ( .B1(n21927), .B2(n8917), .A(n39310), .ZN(n5977) );
  AOI22_X1 U23921 ( .A1(N5678), .A2(n25996), .B1(N5645), .B2(n25901), .ZN(
        n39310) );
  OAI21_X1 U23922 ( .B1(n21933), .B2(n8921), .A(n39320), .ZN(n5978) );
  AOI22_X1 U23923 ( .A1(N5677), .A2(n22873), .B1(N5644), .B2(n25898), .ZN(
        n39320) );
  OAI21_X1 U23924 ( .B1(n21921), .B2(n8925), .A(n39330), .ZN(n5979) );
  AOI22_X1 U23925 ( .A1(N5676), .A2(n26036), .B1(N5643), .B2(n21273), .ZN(
        n39330) );
  OAI21_X1 U23926 ( .B1(n21922), .B2(n8930), .A(n39340), .ZN(n5980) );
  AOI22_X1 U23927 ( .A1(N5675), .A2(n26312), .B1(N5642), .B2(n19211), .ZN(
        n39340) );
  OAI21_X1 U23928 ( .B1(n26349), .B2(n9021), .A(n38760), .ZN(n59360) );
  AOI22_X1 U23929 ( .A1(N5521), .A2(n26033), .B1(N5488), .B2(n25859), .ZN(
        n38760) );
  OAI21_X1 U23930 ( .B1(n26351), .B2(n9026), .A(n38770), .ZN(n59370) );
  AOI22_X1 U23931 ( .A1(N5520), .A2(n24232), .B1(N5487), .B2(n24755), .ZN(
        n38770) );
  OAI21_X1 U23932 ( .B1(n26343), .B2(n9031), .A(n38780), .ZN(n59380) );
  AOI22_X1 U23933 ( .A1(N5519), .A2(n21839), .B1(N5486), .B2(n20550), .ZN(
        n38780) );
  OAI21_X1 U23934 ( .B1(n21906), .B2(n9036), .A(n38790), .ZN(n59390) );
  AOI22_X1 U23935 ( .A1(N5518), .A2(n22835), .B1(N5485), .B2(n20551), .ZN(
        n38790) );
  OAI21_X1 U23936 ( .B1(n26337), .B2(n9041), .A(n38800), .ZN(n59400) );
  AOI22_X1 U23937 ( .A1(N5517), .A2(n22860), .B1(N5484), .B2(n25867), .ZN(
        n38800) );
  OAI21_X1 U23938 ( .B1(n21944), .B2(n9446), .A(n37650), .ZN(n5866) );
  AOI22_X1 U23939 ( .A1(N5085), .A2(n19252), .B1(N5052), .B2(n21274), .ZN(
        n37650) );
  OAI21_X1 U23940 ( .B1(n21931), .B2(n9451), .A(n37660), .ZN(n5867) );
  AOI22_X1 U23941 ( .A1(N5084), .A2(n26042), .B1(N5051), .B2(n21277), .ZN(
        n37660) );
  OAI21_X1 U23942 ( .B1(n21936), .B2(n9456), .A(n37670), .ZN(n5868) );
  AOI22_X1 U23943 ( .A1(N5083), .A2(n22851), .B1(N5050), .B2(n25595), .ZN(
        n37670) );
  OAI21_X1 U23944 ( .B1(n26356), .B2(n9461), .A(n37680), .ZN(n5869) );
  AOI22_X1 U23945 ( .A1(N5082), .A2(n26006), .B1(N5049), .B2(n22886), .ZN(
        n37680) );
  OAI21_X1 U23946 ( .B1(n21926), .B2(n9466), .A(n37690), .ZN(n5870) );
  AOI22_X1 U23947 ( .A1(N5081), .A2(n21848), .B1(N5048), .B2(n24786), .ZN(
        n37690) );
  OAI21_X1 U23948 ( .B1(n26372), .B2(n9471), .A(n37700), .ZN(n5871) );
  AOI22_X1 U23949 ( .A1(N5080), .A2(n26308), .B1(N5047), .B2(n24785), .ZN(
        n37700) );
  OAI21_X1 U23950 ( .B1(n26362), .B2(n9476), .A(n37710), .ZN(n5872) );
  AOI22_X1 U23951 ( .A1(N5079), .A2(n25997), .B1(N5046), .B2(n22888), .ZN(
        n37710) );
  OAI21_X1 U23952 ( .B1(n26365), .B2(n9481), .A(n3772), .ZN(n5873) );
  AOI22_X1 U23953 ( .A1(N5078), .A2(n26043), .B1(N5045), .B2(n25589), .ZN(
        n3772) );
  OAI21_X1 U23954 ( .B1(n26359), .B2(n9490), .A(n3774), .ZN(n5875) );
  AOI22_X1 U23955 ( .A1(N5076), .A2(n26019), .B1(N5043), .B2(n25891), .ZN(
        n3774) );
  OAI21_X1 U23956 ( .B1(n21907), .B2(n9607), .A(n3726), .ZN(n5841) );
  AOI22_X1 U23957 ( .A1(N4906), .A2(n24241), .B1(N4873), .B2(n19245), .ZN(
        n3726) );
  OAI21_X1 U23958 ( .B1(n21913), .B2(n9611), .A(n3727), .ZN(n5842) );
  AOI22_X1 U23959 ( .A1(N4905), .A2(n260101), .B1(N4872), .B2(n25868), .ZN(
        n3727) );
  OAI21_X1 U23960 ( .B1(n21897), .B2(n9615), .A(n3728), .ZN(n58430) );
  AOI22_X1 U23961 ( .A1(N4904), .A2(n22865), .B1(N4871), .B2(n25879), .ZN(
        n3728) );
  OAI21_X1 U23962 ( .B1(n21887), .B2(n9624), .A(n3730), .ZN(n58450) );
  AOI22_X1 U23963 ( .A1(N4902), .A2(n26316), .B1(N4869), .B2(n19205), .ZN(
        n3730) );
  OAI21_X1 U23964 ( .B1(n26371), .B2(n9941), .A(n36010), .ZN(n57560) );
  AOI22_X1 U23965 ( .A1(N4478), .A2(n26039), .B1(N4445), .B2(n27201), .ZN(
        n36010) );
  OAI21_X1 U23966 ( .B1(n26361), .B2(n9945), .A(n36020), .ZN(n57570) );
  AOI22_X1 U23967 ( .A1(N4477), .A2(n22870), .B1(N4444), .B2(n255901), .ZN(
        n36020) );
  OAI21_X1 U23968 ( .B1(n26364), .B2(n9949), .A(n36030), .ZN(n57580) );
  AOI22_X1 U23969 ( .A1(N4476), .A2(n23153), .B1(N4443), .B2(n21268), .ZN(
        n36030) );
  OAI21_X1 U23970 ( .B1(n26355), .B2(n9953), .A(n3604), .ZN(n57590) );
  AOI22_X1 U23971 ( .A1(N4475), .A2(n24247), .B1(N4442), .B2(n25589), .ZN(
        n3604) );
  OAI21_X1 U23972 ( .B1(n26358), .B2(n9957), .A(n3605), .ZN(n57600) );
  AOI22_X1 U23973 ( .A1(N4474), .A2(n26781), .B1(N4441), .B2(n27199), .ZN(
        n3605) );
  OAI21_X1 U23974 ( .B1(n21940), .B2(n9961), .A(n3606), .ZN(n57610) );
  AOI22_X1 U23975 ( .A1(N4473), .A2(n26035), .B1(N4440), .B2(n25890), .ZN(
        n3606) );
  OAI21_X1 U23976 ( .B1(n21927), .B2(n9965), .A(n3607), .ZN(n57620) );
  AOI22_X1 U23977 ( .A1(N4472), .A2(n26021), .B1(N4439), .B2(n25885), .ZN(
        n3607) );
  OAI21_X1 U23978 ( .B1(n21932), .B2(n9969), .A(n3608), .ZN(n57630) );
  AOI22_X1 U23979 ( .A1(N4471), .A2(n26311), .B1(N4438), .B2(n25891), .ZN(
        n3608) );
  OAI21_X1 U23980 ( .B1(n21917), .B2(n9973), .A(n3609), .ZN(n57640) );
  AOI22_X1 U23981 ( .A1(N4470), .A2(n26313), .B1(N4437), .B2(n25886), .ZN(
        n3609) );
  OAI21_X1 U23982 ( .B1(n21922), .B2(n9977), .A(n3610), .ZN(n57650) );
  AOI22_X1 U23983 ( .A1(N4469), .A2(n23146), .B1(N4436), .B2(n19246), .ZN(
        n3610) );
  OAI21_X1 U23984 ( .B1(n21911), .B2(n10114), .A(n3562), .ZN(n57310) );
  AOI22_X1 U23985 ( .A1(N4305), .A2(n19253), .B1(N4272), .B2(n25583), .ZN(
        n3562) );
  OAI21_X1 U23986 ( .B1(n21916), .B2(n10119), .A(n3563), .ZN(n57320) );
  AOI22_X1 U23987 ( .A1(N4304), .A2(n26071), .B1(N4271), .B2(n19205), .ZN(
        n3563) );
  OAI21_X1 U23988 ( .B1(n21901), .B2(n10124), .A(n3564), .ZN(n57330) );
  AOI22_X1 U23989 ( .A1(N4303), .A2(n22847), .B1(N4270), .B2(n25580), .ZN(
        n3564) );
  OAI21_X1 U23990 ( .B1(n26347), .B2(n10129), .A(n3565), .ZN(n57340) );
  AOI22_X1 U23991 ( .A1(N4302), .A2(n26015), .B1(N4269), .B2(n24494), .ZN(
        n3565) );
  OAI21_X1 U23992 ( .B1(n21891), .B2(n10134), .A(n3566), .ZN(n57350) );
  AOI22_X1 U23993 ( .A1(N4301), .A2(n26318), .B1(N4268), .B2(n25581), .ZN(
        n3566) );
  OAI21_X1 U23994 ( .B1(n26350), .B2(n10139), .A(n3567), .ZN(n57360) );
  AOI22_X1 U23995 ( .A1(N4300), .A2(n26310), .B1(N4267), .B2(n24749), .ZN(
        n3567) );
  OAI21_X1 U23996 ( .B1(n26353), .B2(n10144), .A(n3568), .ZN(n5737) );
  AOI22_X1 U23997 ( .A1(N4299), .A2(n260101), .B1(N4266), .B2(n25578), .ZN(
        n3568) );
  OAI21_X1 U23998 ( .B1(n26344), .B2(n10149), .A(n3569), .ZN(n5738) );
  AOI22_X1 U23999 ( .A1(N4298), .A2(n26061), .B1(N4265), .B2(n21250), .ZN(
        n3569) );
  OAI21_X1 U24000 ( .B1(n26338), .B2(n10158), .A(n3571), .ZN(n5740) );
  AOI22_X1 U24001 ( .A1(N4296), .A2(n26032), .B1(N4263), .B2(n25864), .ZN(
        n3571) );
  OAI21_X1 U24002 ( .B1(n21943), .B2(n10489), .A(n3444), .ZN(n56510) );
  AOI22_X1 U24003 ( .A1(N3885), .A2(n26005), .B1(N3852), .B2(n24466), .ZN(
        n3444) );
  OAI21_X1 U24004 ( .B1(n21930), .B2(n10494), .A(n3445), .ZN(n56520) );
  AOI22_X1 U24005 ( .A1(N3884), .A2(n22866), .B1(N3851), .B2(n19246), .ZN(
        n3445) );
  OAI21_X1 U24006 ( .B1(n21935), .B2(n10499), .A(n3446), .ZN(n56530) );
  AOI22_X1 U24007 ( .A1(N3883), .A2(n26018), .B1(N3850), .B2(n25902), .ZN(
        n3446) );
  OAI21_X1 U24008 ( .B1(n21920), .B2(n10504), .A(n3447), .ZN(n56540) );
  AOI22_X1 U24009 ( .A1(N3882), .A2(n26307), .B1(N3849), .B2(n25897), .ZN(
        n3447) );
  OAI21_X1 U24010 ( .B1(n21925), .B2(n10509), .A(n3448), .ZN(n56550) );
  AOI22_X1 U24011 ( .A1(N3881), .A2(n26041), .B1(N3848), .B2(n25594), .ZN(
        n3448) );
  OAI21_X1 U24012 ( .B1(n26349), .B2(n10660), .A(n3397), .ZN(n5621) );
  AOI22_X1 U24013 ( .A1(N3714), .A2(n22833), .B1(N3681), .B2(n24749), .ZN(
        n3397) );
  OAI21_X1 U24014 ( .B1(n26352), .B2(n10664), .A(n3398), .ZN(n5622) );
  AOI22_X1 U24015 ( .A1(N3713), .A2(n23164), .B1(N3680), .B2(n20544), .ZN(
        n3398) );
  OAI21_X1 U24016 ( .B1(n26343), .B2(n10668), .A(n3399), .ZN(n5623) );
  AOI22_X1 U24017 ( .A1(N3712), .A2(n24249), .B1(N3679), .B2(n20549), .ZN(
        n3399) );
  OAI21_X1 U24018 ( .B1(n26346), .B2(n10672), .A(n3400), .ZN(n5624) );
  AOI22_X1 U24019 ( .A1(N3711), .A2(n22848), .B1(N3678), .B2(n21250), .ZN(
        n3400) );
  OAI21_X1 U24020 ( .B1(n26337), .B2(n10676), .A(n3401), .ZN(n5625) );
  AOI22_X1 U24021 ( .A1(N3710), .A2(n22862), .B1(N3677), .B2(n24752), .ZN(
        n3401) );
  OAI21_X1 U24022 ( .B1(n21907), .B2(n10680), .A(n3402), .ZN(n5626) );
  AOI22_X1 U24023 ( .A1(N3709), .A2(n23203), .B1(N3676), .B2(n25863), .ZN(
        n3402) );
  OAI21_X1 U24024 ( .B1(n21912), .B2(n10684), .A(n3403), .ZN(n5627) );
  AOI22_X1 U24025 ( .A1(N3708), .A2(n26034), .B1(N3675), .B2(n25859), .ZN(
        n3403) );
  OAI21_X1 U24026 ( .B1(n21897), .B2(n10688), .A(n3404), .ZN(n5628) );
  AOI22_X1 U24027 ( .A1(N3707), .A2(n26315), .B1(N3674), .B2(n25864), .ZN(
        n3404) );
  OAI21_X1 U24028 ( .B1(n21902), .B2(n10692), .A(n3405), .ZN(n5629) );
  AOI22_X1 U24029 ( .A1(N3706), .A2(n26317), .B1(N3673), .B2(n25860), .ZN(
        n3405) );
  OAI21_X1 U24030 ( .B1(n21887), .B2(n10696), .A(n3406), .ZN(n5630) );
  AOI22_X1 U24031 ( .A1(N3705), .A2(n24252), .B1(N3672), .B2(n24754), .ZN(
        n3406) );
  OAI21_X1 U24032 ( .B1(n21910), .B2(n11192), .A(n3237), .ZN(n55160) );
  AOI22_X1 U24033 ( .A1(N3128), .A2(n26014), .B1(N3095), .B2(n24486), .ZN(
        n3237) );
  OAI21_X1 U24034 ( .B1(n21915), .B2(n11197), .A(n3238), .ZN(n55170) );
  AOI22_X1 U24035 ( .A1(N3127), .A2(n26775), .B1(N3094), .B2(n24490), .ZN(
        n3238) );
  OAI21_X1 U24036 ( .B1(n21900), .B2(n11202), .A(n3239), .ZN(n55180) );
  AOI22_X1 U24037 ( .A1(N3126), .A2(n26031), .B1(N3093), .B2(n25868), .ZN(
        n3239) );
  OAI21_X1 U24038 ( .B1(n21905), .B2(n11207), .A(n3240), .ZN(n55190) );
  AOI22_X1 U24039 ( .A1(N3125), .A2(n26309), .B1(N3092), .B2(n25877), .ZN(
        n3240) );
  OAI21_X1 U24040 ( .B1(n21890), .B2(n11212), .A(n3241), .ZN(n55200) );
  AOI22_X1 U24041 ( .A1(N3124), .A2(n260701), .B1(N3091), .B2(n21262), .ZN(
        n3241) );
  OAI21_X1 U24042 ( .B1(n21543), .B2(n16922), .A(n45240), .ZN(n63560) );
  AOI22_X1 U24043 ( .A1(N7911), .A2(n17100), .B1(N7878), .B2(n27138), .ZN(
        n45240) );
  OAI21_X1 U24044 ( .B1(n21530), .B2(n16991), .A(n45250), .ZN(n63570) );
  AOI22_X1 U24045 ( .A1(N7910), .A2(n25959), .B1(N7877), .B2(n27137), .ZN(
        n45250) );
  OAI21_X1 U24046 ( .B1(n21534), .B2(n17006), .A(n45260), .ZN(n63580) );
  AOI22_X1 U24047 ( .A1(N7909), .A2(n25966), .B1(N7876), .B2(n19321), .ZN(
        n45260) );
  OAI21_X1 U24048 ( .B1(n21545), .B2(n16996), .A(n45270), .ZN(n63590) );
  AOI22_X1 U24049 ( .A1(N7908), .A2(n259601), .B1(N7875), .B2(n27139), .ZN(
        n45270) );
  OAI21_X1 U24050 ( .B1(n21532), .B2(n16986), .A(n45280), .ZN(n63600) );
  AOI22_X1 U24051 ( .A1(N7907), .A2(n21444), .B1(N7874), .B2(n27138), .ZN(
        n45280) );
  OAI21_X1 U24052 ( .B1(n21536), .B2(n16897), .A(n4529), .ZN(n63610) );
  AOI22_X1 U24053 ( .A1(N7906), .A2(n25674), .B1(N7873), .B2(n27137), .ZN(
        n4529) );
  OAI21_X1 U24054 ( .B1(n26103), .B2(n16947), .A(n4530), .ZN(n63620) );
  AOI22_X1 U24055 ( .A1(N7905), .A2(n20514), .B1(N7872), .B2(n19321), .ZN(
        n4530) );
  OAI21_X1 U24056 ( .B1(n26095), .B2(n16878), .A(n4531), .ZN(n63630) );
  AOI22_X1 U24057 ( .A1(N7904), .A2(n25675), .B1(N7871), .B2(n27144), .ZN(
        n4531) );
  OAI21_X1 U24058 ( .B1(n26098), .B2(n16854), .A(n4532), .ZN(n63640) );
  AOI22_X1 U24059 ( .A1(N7903), .A2(n20534), .B1(N7870), .B2(n27136), .ZN(
        n4532) );
  OAI21_X1 U24060 ( .B1(n26104), .B2(n16902), .A(n4533), .ZN(n63650) );
  AOI22_X1 U24061 ( .A1(N7902), .A2(n25675), .B1(N7869), .B2(n27135), .ZN(
        n4533) );
  OAI21_X1 U24062 ( .B1(n26096), .B2(n16961), .A(n4534), .ZN(n63660) );
  AOI22_X1 U24063 ( .A1(N7901), .A2(n21440), .B1(N7868), .B2(n27134), .ZN(
        n4534) );
  OAI21_X1 U24064 ( .B1(n26099), .B2(n16942), .A(n4535), .ZN(n63670) );
  AOI22_X1 U24065 ( .A1(N7900), .A2(n25964), .B1(N7867), .B2(n27133), .ZN(
        n4535) );
  OAI21_X1 U24066 ( .B1(n21544), .B2(n16887), .A(n4536), .ZN(n63680) );
  AOI22_X1 U24067 ( .A1(N7899), .A2(n20529), .B1(N7866), .B2(n27132), .ZN(
        n4536) );
  OAI21_X1 U24068 ( .B1(n21529), .B2(n16932), .A(n4537), .ZN(n63690) );
  AOI22_X1 U24069 ( .A1(N7898), .A2(n24741), .B1(N7865), .B2(n27131), .ZN(
        n4537) );
  OAI21_X1 U24070 ( .B1(n21533), .B2(n16956), .A(n4538), .ZN(n63700) );
  AOI22_X1 U24071 ( .A1(N7897), .A2(n25958), .B1(N7864), .B2(n19320), .ZN(
        n4538) );
  OAI21_X1 U24072 ( .B1(n21546), .B2(n16971), .A(n43550), .ZN(n6251) );
  AOI22_X1 U24073 ( .A1(N7318), .A2(n25959), .B1(N7285), .B2(n27135), .ZN(
        n43550) );
  OAI21_X1 U24074 ( .B1(n21531), .B2(n7514), .A(n43560), .ZN(n6252) );
  AOI22_X1 U24075 ( .A1(N7317), .A2(n25965), .B1(N7284), .B2(n27134), .ZN(
        n43560) );
  OAI21_X1 U24076 ( .B1(n21537), .B2(n16937), .A(n43570), .ZN(n6253) );
  AOI22_X1 U24077 ( .A1(N7316), .A2(n20521), .B1(N7283), .B2(n27133), .ZN(
        n43570) );
  OAI21_X1 U24078 ( .B1(n26103), .B2(n16912), .A(n4358), .ZN(n6254) );
  AOI22_X1 U24079 ( .A1(N7315), .A2(n24738), .B1(N7282), .B2(n27132), .ZN(
        n4358) );
  OAI21_X1 U24080 ( .B1(n26095), .B2(n17001), .A(n4359), .ZN(n6255) );
  AOI22_X1 U24081 ( .A1(N7314), .A2(n259601), .B1(N7281), .B2(n27131), .ZN(
        n4359) );
  OAI21_X1 U24082 ( .B1(n26098), .B2(n16952), .A(n4360), .ZN(n6256) );
  AOI22_X1 U24083 ( .A1(N7313), .A2(n20535), .B1(N7280), .B2(n19320), .ZN(
        n4360) );
  OAI21_X1 U24084 ( .B1(n26104), .B2(n16917), .A(n4361), .ZN(n6257) );
  AOI22_X1 U24085 ( .A1(N7312), .A2(n20522), .B1(N7279), .B2(n27144), .ZN(
        n4361) );
  OAI21_X1 U24086 ( .B1(n26096), .B2(n16966), .A(n4362), .ZN(n6258) );
  AOI22_X1 U24087 ( .A1(N7311), .A2(n21439), .B1(N7278), .B2(n27143), .ZN(
        n4362) );
  OAI21_X1 U24088 ( .B1(n26099), .B2(n16976), .A(n4363), .ZN(n6259) );
  AOI22_X1 U24089 ( .A1(N7310), .A2(n25966), .B1(N7277), .B2(n27142), .ZN(
        n4363) );
  OAI21_X1 U24090 ( .B1(n21543), .B2(n16892), .A(n4364), .ZN(n6260) );
  AOI22_X1 U24091 ( .A1(N7309), .A2(n17100), .B1(N7276), .B2(n27141), .ZN(
        n4364) );
  OAI21_X1 U24092 ( .B1(n21529), .B2(n16981), .A(n4365), .ZN(n62610) );
  AOI22_X1 U24093 ( .A1(N7308), .A2(n21443), .B1(N7275), .B2(n27143), .ZN(
        n4365) );
  OAI21_X1 U24094 ( .B1(n21533), .B2(n16869), .A(n4366), .ZN(n62620) );
  AOI22_X1 U24095 ( .A1(N7307), .A2(n19242), .B1(N7274), .B2(n27140), .ZN(
        n4366) );
  OAI21_X1 U24096 ( .B1(n21545), .B2(n16907), .A(n4367), .ZN(n62630) );
  AOI22_X1 U24097 ( .A1(N7306), .A2(n20528), .B1(N7273), .B2(n27142), .ZN(
        n4367) );
  OAI21_X1 U24098 ( .B1(n21531), .B2(n16927), .A(n4368), .ZN(n62640) );
  AOI22_X1 U24099 ( .A1(N7305), .A2(n17098), .B1(N7272), .B2(n27136), .ZN(
        n4368) );
  OAI21_X1 U24100 ( .B1(n21536), .B2(n16882), .A(n4369), .ZN(n62650) );
  AOI22_X1 U24101 ( .A1(N7304), .A2(n20513), .B1(N7271), .B2(n27139), .ZN(
        n4369) );
  OAI21_X1 U24102 ( .B1(n21521), .B2(n11045), .A(n3284), .ZN(n5546) );
  AOI22_X1 U24103 ( .A1(N3299), .A2(n17099), .B1(N3266), .B2(n27286), .ZN(
        n3284) );
  OAI21_X1 U24104 ( .B1(n21526), .B2(n11050), .A(n32850), .ZN(n5547) );
  AOI22_X1 U24105 ( .A1(N3298), .A2(n25962), .B1(N3265), .B2(n27285), .ZN(
        n32850) );
  OAI21_X1 U24106 ( .B1(n21513), .B2(n11055), .A(n32860), .ZN(n5548) );
  AOI22_X1 U24107 ( .A1(N3297), .A2(n25969), .B1(N3264), .B2(n19324), .ZN(
        n32860) );
  OAI21_X1 U24108 ( .B1(n21523), .B2(n11060), .A(n32870), .ZN(n5549) );
  AOI22_X1 U24109 ( .A1(N3296), .A2(n25963), .B1(N3263), .B2(n27287), .ZN(
        n32870) );
  OAI21_X1 U24110 ( .B1(n21527), .B2(n11065), .A(n32880), .ZN(n5550) );
  AOI22_X1 U24111 ( .A1(N3295), .A2(n21446), .B1(N3262), .B2(n27286), .ZN(
        n32880) );
  OAI21_X1 U24112 ( .B1(n21516), .B2(n11070), .A(n32890), .ZN(n5551) );
  AOI22_X1 U24113 ( .A1(N3294), .A2(n25676), .B1(N3261), .B2(n27285), .ZN(
        n32890) );
  OAI21_X1 U24114 ( .B1(n26092), .B2(n11075), .A(n32900), .ZN(n5552) );
  AOI22_X1 U24115 ( .A1(N3293), .A2(n20510), .B1(N3260), .B2(n19324), .ZN(
        n32900) );
  OAI21_X1 U24116 ( .B1(n17076), .B2(n11080), .A(n32910), .ZN(n55530) );
  AOI22_X1 U24117 ( .A1(N3292), .A2(n25677), .B1(N3259), .B2(n27292), .ZN(
        n32910) );
  OAI21_X1 U24118 ( .B1(n26087), .B2(n11085), .A(n32920), .ZN(n55540) );
  AOI22_X1 U24119 ( .A1(N3291), .A2(n20537), .B1(N3258), .B2(n27284), .ZN(
        n32920) );
  OAI21_X1 U24120 ( .B1(n26093), .B2(n11090), .A(n32930), .ZN(n55550) );
  AOI22_X1 U24121 ( .A1(N3290), .A2(n25677), .B1(N3257), .B2(n27283), .ZN(
        n32930) );
  OAI21_X1 U24122 ( .B1(n26094), .B2(n11095), .A(n32940), .ZN(n55560) );
  AOI22_X1 U24123 ( .A1(N3289), .A2(n21442), .B1(N3256), .B2(n27282), .ZN(
        n32940) );
  OAI21_X1 U24124 ( .B1(n26088), .B2(n11100), .A(n32950), .ZN(n55570) );
  AOI22_X1 U24125 ( .A1(N3288), .A2(n25967), .B1(N3255), .B2(n27281), .ZN(
        n32950) );
  OAI21_X1 U24126 ( .B1(n21520), .B2(n11105), .A(n32960), .ZN(n55580) );
  AOI22_X1 U24127 ( .A1(N3287), .A2(n20532), .B1(N3254), .B2(n27280), .ZN(
        n32960) );
  OAI21_X1 U24128 ( .B1(n21525), .B2(n11110), .A(n32970), .ZN(n55590) );
  AOI22_X1 U24129 ( .A1(N3286), .A2(n24743), .B1(N3253), .B2(n27279), .ZN(
        n32970) );
  OAI21_X1 U24130 ( .B1(n21512), .B2(n11114), .A(n32980), .ZN(n55600) );
  AOI22_X1 U24131 ( .A1(N3285), .A2(n25961), .B1(N3252), .B2(n19323), .ZN(
        n32980) );
  OAI21_X1 U24132 ( .B1(n21522), .B2(n11579), .A(n3112), .ZN(n5441) );
  AOI22_X1 U24133 ( .A1(N2688), .A2(n25962), .B1(N2655), .B2(n27283), .ZN(
        n3112) );
  OAI21_X1 U24134 ( .B1(n21528), .B2(n11584), .A(n3113), .ZN(n5442) );
  AOI22_X1 U24135 ( .A1(N2687), .A2(n25968), .B1(N2654), .B2(n27282), .ZN(
        n3113) );
  OAI21_X1 U24136 ( .B1(n21515), .B2(n11589), .A(n31140), .ZN(n5443) );
  AOI22_X1 U24137 ( .A1(N2686), .A2(n20516), .B1(N2653), .B2(n27281), .ZN(
        n31140) );
  OAI21_X1 U24138 ( .B1(n26092), .B2(n11594), .A(n31150), .ZN(n5444) );
  AOI22_X1 U24139 ( .A1(N2685), .A2(n24739), .B1(N2652), .B2(n27280), .ZN(
        n31150) );
  OAI21_X1 U24140 ( .B1(n17076), .B2(n11599), .A(n31160), .ZN(n5445) );
  AOI22_X1 U24141 ( .A1(N2684), .A2(n25963), .B1(N2651), .B2(n27279), .ZN(
        n31160) );
  OAI21_X1 U24142 ( .B1(n26087), .B2(n11604), .A(n31170), .ZN(n5446) );
  AOI22_X1 U24143 ( .A1(N2683), .A2(n20538), .B1(N2650), .B2(n19323), .ZN(
        n31170) );
  OAI21_X1 U24144 ( .B1(n26093), .B2(n11609), .A(n31180), .ZN(n5447) );
  AOI22_X1 U24145 ( .A1(N2682), .A2(n20517), .B1(N2649), .B2(n27292), .ZN(
        n31180) );
  OAI21_X1 U24146 ( .B1(n26094), .B2(n11614), .A(n31190), .ZN(n5448) );
  AOI22_X1 U24147 ( .A1(N2681), .A2(n21441), .B1(N2648), .B2(n27291), .ZN(
        n31190) );
  OAI21_X1 U24148 ( .B1(n26088), .B2(n11619), .A(n31200), .ZN(n5449) );
  AOI22_X1 U24149 ( .A1(N2680), .A2(n25969), .B1(N2647), .B2(n272901), .ZN(
        n31200) );
  OAI21_X1 U24150 ( .B1(n21520), .B2(n11624), .A(n31210), .ZN(n5450) );
  AOI22_X1 U24151 ( .A1(N2679), .A2(n17099), .B1(N2646), .B2(n27289), .ZN(
        n31210) );
  OAI21_X1 U24152 ( .B1(n21525), .B2(n11629), .A(n31220), .ZN(n5451) );
  AOI22_X1 U24153 ( .A1(N2678), .A2(n21445), .B1(N2645), .B2(n27291), .ZN(
        n31220) );
  OAI21_X1 U24154 ( .B1(n21512), .B2(n11634), .A(n31230), .ZN(n5452) );
  AOI22_X1 U24155 ( .A1(N2677), .A2(n19243), .B1(N2644), .B2(n27288), .ZN(
        n31230) );
  OAI21_X1 U24156 ( .B1(n21522), .B2(n11639), .A(n31240), .ZN(n5453) );
  AOI22_X1 U24157 ( .A1(N2676), .A2(n20531), .B1(N2643), .B2(n272901), .ZN(
        n31240) );
  OAI21_X1 U24158 ( .B1(n21527), .B2(n11644), .A(n31250), .ZN(n5454) );
  AOI22_X1 U24159 ( .A1(N2675), .A2(n17101), .B1(N2642), .B2(n27284), .ZN(
        n31250) );
  OAI21_X1 U24160 ( .B1(n21515), .B2(n11648), .A(n31260), .ZN(n5455) );
  AOI22_X1 U24161 ( .A1(N2674), .A2(n20509), .B1(N2641), .B2(n27287), .ZN(
        n31260) );
  NAND2_X1 U24162 ( .A1(n50070), .A2(n50080), .ZN(mul_outcome[37]) );
  AOI221_X1 U24163 ( .B1(n21892), .B2(n17867), .C1(n22839), .C2(n17855), .A(
        n50100), .ZN(n50070) );
  AOI221_X1 U24164 ( .B1(n21877), .B2(n17891), .C1(n21882), .C2(n17879), .A(
        n50090), .ZN(n50080) );
  OAI22_X1 U24165 ( .A1(n2068), .A2(n19209), .B1(n2047), .B2(n19199), .ZN(
        n50100) );
  NAND2_X1 U24166 ( .A1(n50030), .A2(n50040), .ZN(mul_outcome[38]) );
  AOI221_X1 U24167 ( .B1(n26339), .B2(n17865), .C1(n26002), .C2(n17853), .A(
        n50060), .ZN(n50030) );
  AOI221_X1 U24168 ( .B1(n26330), .B2(n17889), .C1(n26333), .C2(n17877), .A(
        n50050), .ZN(n50040) );
  OAI22_X1 U24169 ( .A1(n2067), .A2(n21264), .B1(n2046), .B2(n21227), .ZN(
        n50060) );
  OAI21_X1 U24170 ( .B1(n21588), .B2(n3054), .A(n4402), .ZN(n62810) );
  AOI22_X1 U24171 ( .A1(N7486), .A2(n23185), .B1(N7453), .B2(n25889), .ZN(
        n4402) );
  OAI21_X1 U24172 ( .B1(n21591), .B2(n3059), .A(n4403), .ZN(n6282) );
  AOI22_X1 U24173 ( .A1(N7485), .A2(n22869), .B1(N7452), .B2(n25886), .ZN(
        n4403) );
  OAI21_X1 U24174 ( .B1(n21580), .B2(n3064), .A(n4404), .ZN(n6283) );
  AOI22_X1 U24175 ( .A1(N7484), .A2(n19255), .B1(N7451), .B2(n24794), .ZN(
        n4404) );
  OAI21_X1 U24176 ( .B1(n21584), .B2(n3069), .A(n4405), .ZN(n6284) );
  AOI22_X1 U24177 ( .A1(N7483), .A2(n24238), .B1(N7450), .B2(n25893), .ZN(
        n4405) );
  OAI21_X1 U24178 ( .B1(n21572), .B2(n3110), .A(n4406), .ZN(n6285) );
  AOI22_X1 U24179 ( .A1(N7482), .A2(n22875), .B1(N7449), .B2(n24794), .ZN(
        n4406) );
  OAI21_X1 U24180 ( .B1(n21590), .B2(n7845), .A(n4252), .ZN(n61860) );
  AOI22_X1 U24181 ( .A1(N6878), .A2(n21850), .B1(N6845), .B2(n25902), .ZN(
        n4252) );
  OAI21_X1 U24182 ( .B1(n21593), .B2(n7849), .A(n4253), .ZN(n61870) );
  AOI22_X1 U24183 ( .A1(N6877), .A2(n21843), .B1(N6844), .B2(n25899), .ZN(
        n4253) );
  OAI21_X1 U24184 ( .B1(n21582), .B2(n7853), .A(n4254), .ZN(n61880) );
  AOI22_X1 U24185 ( .A1(N6876), .A2(n260201), .B1(N6843), .B2(n25594), .ZN(
        n4254) );
  OAI21_X1 U24186 ( .B1(n21574), .B2(n7862), .A(n4256), .ZN(n61900) );
  AOI22_X1 U24187 ( .A1(N6874), .A2(n21838), .B1(N6841), .B2(n255901), .ZN(
        n4256) );
  OAI21_X1 U24188 ( .B1(n21575), .B2(n79530), .A(n4194), .ZN(n6146) );
  AOI22_X1 U24189 ( .A1(N6714), .A2(n26761), .B1(N6681), .B2(n25865), .ZN(
        n4194) );
  OAI21_X1 U24190 ( .B1(n21564), .B2(n79580), .A(n4195), .ZN(n6147) );
  AOI22_X1 U24191 ( .A1(N6713), .A2(n22856), .B1(N6680), .B2(n25860), .ZN(
        n4195) );
  OAI21_X1 U24192 ( .B1(n21567), .B2(n7963), .A(n4196), .ZN(n6148) );
  AOI22_X1 U24193 ( .A1(N6712), .A2(n19256), .B1(N6679), .B2(n24491), .ZN(
        n4196) );
  OAI21_X1 U24194 ( .B1(n21556), .B2(n7968), .A(n4197), .ZN(n61490) );
  AOI22_X1 U24195 ( .A1(N6711), .A2(n19257), .B1(N6678), .B2(n24489), .ZN(
        n4197) );
  OAI21_X1 U24196 ( .B1(n21560), .B2(n7973), .A(n4198), .ZN(n61500) );
  AOI22_X1 U24197 ( .A1(N6710), .A2(n22864), .B1(N6677), .B2(n24488), .ZN(
        n4198) );
  OAI21_X1 U24198 ( .B1(n26125), .B2(n8352), .A(n4086), .ZN(n6076) );
  AOI22_X1 U24199 ( .A1(N6270), .A2(n26004), .B1(N6237), .B2(n25898), .ZN(
        n4086) );
  OAI21_X1 U24200 ( .B1(n26127), .B2(n8357), .A(n4087), .ZN(n6077) );
  AOI22_X1 U24201 ( .A1(N6269), .A2(n26773), .B1(N6236), .B2(n19210), .ZN(
        n4087) );
  OAI21_X1 U24202 ( .B1(n26121), .B2(n8362), .A(n4088), .ZN(n6078) );
  AOI22_X1 U24203 ( .A1(N6268), .A2(n25996), .B1(N6235), .B2(n25592), .ZN(
        n4088) );
  OAI21_X1 U24204 ( .B1(n21586), .B2(n8367), .A(n4089), .ZN(n6079) );
  AOI22_X1 U24205 ( .A1(N6267), .A2(n260401), .B1(N6234), .B2(n25593), .ZN(
        n4089) );
  OAI21_X1 U24206 ( .B1(n26117), .B2(n8372), .A(n4090), .ZN(n6080) );
  AOI22_X1 U24207 ( .A1(N6266), .A2(n22854), .B1(N6233), .B2(n22883), .ZN(
        n4090) );
  OAI21_X1 U24208 ( .B1(n26126), .B2(n8377), .A(n4091), .ZN(n6081) );
  AOI22_X1 U24209 ( .A1(N6265), .A2(n26778), .B1(N6232), .B2(n20587), .ZN(
        n4091) );
  OAI21_X1 U24210 ( .B1(n26128), .B2(n8382), .A(n4092), .ZN(n6082) );
  AOI22_X1 U24211 ( .A1(N6264), .A2(n21847), .B1(N6231), .B2(n22881), .ZN(
        n4092) );
  OAI21_X1 U24212 ( .B1(n26122), .B2(n8387), .A(n4093), .ZN(n6083) );
  AOI22_X1 U24213 ( .A1(N6263), .A2(n23147), .B1(N6230), .B2(n25588), .ZN(
        n4093) );
  OAI21_X1 U24214 ( .B1(n26118), .B2(n8396), .A(n40950), .ZN(n6085) );
  AOI22_X1 U24215 ( .A1(N6261), .A2(n21484), .B1(N6228), .B2(n25887), .ZN(
        n40950) );
  OAI21_X1 U24216 ( .B1(n21577), .B2(n8537), .A(n40470), .ZN(n6051) );
  AOI22_X1 U24217 ( .A1(N6097), .A2(n21857), .B1(N6064), .B2(n25869), .ZN(
        n40470) );
  OAI21_X1 U24218 ( .B1(n21566), .B2(n8542), .A(n40480), .ZN(n6052) );
  AOI22_X1 U24219 ( .A1(N6096), .A2(n21851), .B1(N6063), .B2(n25878), .ZN(
        n40480) );
  OAI21_X1 U24220 ( .B1(n21569), .B2(n8547), .A(n40490), .ZN(n6053) );
  AOI22_X1 U24221 ( .A1(N6095), .A2(n21480), .B1(N6062), .B2(n19207), .ZN(
        n40490) );
  OAI21_X1 U24222 ( .B1(n21562), .B2(n8556), .A(n40510), .ZN(n6055) );
  AOI22_X1 U24223 ( .A1(N6093), .A2(n21842), .B1(N6060), .B2(n21256), .ZN(
        n40510) );
  OAI21_X1 U24224 ( .B1(n21587), .B2(n8873), .A(n3920), .ZN(n5966) );
  AOI22_X1 U24225 ( .A1(N5689), .A2(n23184), .B1(N5656), .B2(n25592), .ZN(
        n3920) );
  OAI21_X1 U24226 ( .B1(n21592), .B2(n8877), .A(n3921), .ZN(n5967) );
  AOI22_X1 U24227 ( .A1(N5688), .A2(n25998), .B1(N5655), .B2(n25593), .ZN(
        n3921) );
  OAI21_X1 U24228 ( .B1(n21579), .B2(n8881), .A(n3922), .ZN(n5968) );
  AOI22_X1 U24229 ( .A1(N5687), .A2(n22843), .B1(N5654), .B2(n24785), .ZN(
        n3922) );
  OAI21_X1 U24230 ( .B1(n26123), .B2(n8885), .A(n3923), .ZN(n5969) );
  AOI22_X1 U24231 ( .A1(N5686), .A2(n26008), .B1(N5653), .B2(n24789), .ZN(
        n3923) );
  OAI21_X1 U24232 ( .B1(n21571), .B2(n8889), .A(n3924), .ZN(n5970) );
  AOI22_X1 U24233 ( .A1(N5685), .A2(n26312), .B1(N5652), .B2(n24789), .ZN(
        n3924) );
  OAI21_X1 U24234 ( .B1(n21589), .B2(n8893), .A(n3925), .ZN(n5971) );
  AOI22_X1 U24235 ( .A1(N5684), .A2(n26019), .B1(N5651), .B2(n21269), .ZN(
        n3925) );
  OAI21_X1 U24236 ( .B1(n21594), .B2(n8897), .A(n3926), .ZN(n5972) );
  AOI22_X1 U24237 ( .A1(N5683), .A2(n21836), .B1(N5650), .B2(n25888), .ZN(
        n3926) );
  OAI21_X1 U24238 ( .B1(n21581), .B2(n8901), .A(n39270), .ZN(n5973) );
  AOI22_X1 U24239 ( .A1(N5682), .A2(n26041), .B1(N5649), .B2(n25887), .ZN(
        n39270) );
  OAI21_X1 U24240 ( .B1(n26124), .B2(n8905), .A(n39280), .ZN(n5974) );
  AOI22_X1 U24241 ( .A1(N5681), .A2(n22855), .B1(N5648), .B2(n25895), .ZN(
        n39280) );
  OAI21_X1 U24242 ( .B1(n21573), .B2(n8909), .A(n39290), .ZN(n5975) );
  AOI22_X1 U24243 ( .A1(N5680), .A2(n26005), .B1(N5647), .B2(n25892), .ZN(
        n39290) );
  OAI21_X1 U24244 ( .B1(n26119), .B2(n9046), .A(n38810), .ZN(n59410) );
  AOI22_X1 U24245 ( .A1(N5516), .A2(n21471), .B1(N5483), .B2(n25879), .ZN(
        n38810) );
  OAI21_X1 U24246 ( .B1(n26113), .B2(n9051), .A(n38820), .ZN(n59420) );
  AOI22_X1 U24247 ( .A1(N5515), .A2(n26769), .B1(N5482), .B2(n25583), .ZN(
        n38820) );
  OAI21_X1 U24248 ( .B1(n26115), .B2(n9056), .A(n38830), .ZN(n59430) );
  AOI22_X1 U24249 ( .A1(N5514), .A2(n26009), .B1(N5481), .B2(n20547), .ZN(
        n38830) );
  OAI21_X1 U24250 ( .B1(n21558), .B2(n9061), .A(n38840), .ZN(n59440) );
  AOI22_X1 U24251 ( .A1(N5513), .A2(n26069), .B1(N5480), .B2(n20546), .ZN(
        n38840) );
  OAI21_X1 U24252 ( .B1(n26111), .B2(n9066), .A(n38850), .ZN(n59450) );
  AOI22_X1 U24253 ( .A1(N5512), .A2(n24241), .B1(N5479), .B2(n20545), .ZN(
        n38850) );
  OAI21_X1 U24254 ( .B1(n261201), .B2(n9071), .A(n38860), .ZN(n5946) );
  AOI22_X1 U24255 ( .A1(N5511), .A2(n22857), .B1(N5478), .B2(n22892), .ZN(
        n38860) );
  OAI21_X1 U24256 ( .B1(n26114), .B2(n9076), .A(n38870), .ZN(n5947) );
  AOI22_X1 U24257 ( .A1(N5510), .A2(n21855), .B1(N5477), .B2(n25579), .ZN(
        n38870) );
  OAI21_X1 U24258 ( .B1(n26116), .B2(n9081), .A(n38880), .ZN(n5948) );
  AOI22_X1 U24259 ( .A1(N5509), .A2(n23159), .B1(N5476), .B2(n25578), .ZN(
        n38880) );
  OAI21_X1 U24260 ( .B1(n26112), .B2(n9090), .A(n38900), .ZN(n5950) );
  AOI22_X1 U24261 ( .A1(N5507), .A2(n21494), .B1(N5474), .B2(n25861), .ZN(
        n38900) );
  OAI21_X1 U24262 ( .B1(n26125), .B2(n9421), .A(n37600), .ZN(n58610) );
  AOI22_X1 U24263 ( .A1(N5090), .A2(n25995), .B1(N5057), .B2(n25893), .ZN(
        n37600) );
  OAI21_X1 U24264 ( .B1(n26127), .B2(n9426), .A(n37610), .ZN(n58620) );
  AOI22_X1 U24265 ( .A1(N5089), .A2(n26045), .B1(N5056), .B2(n24467), .ZN(
        n37610) );
  OAI21_X1 U24266 ( .B1(n26121), .B2(n9431), .A(n37620), .ZN(n58630) );
  AOI22_X1 U24267 ( .A1(N5088), .A2(n26007), .B1(N5055), .B2(n24792), .ZN(
        n37620) );
  OAI21_X1 U24268 ( .B1(n21583), .B2(n9436), .A(n37630), .ZN(n5864) );
  AOI22_X1 U24269 ( .A1(N5087), .A2(n24255), .B1(N5054), .B2(n25903), .ZN(
        n37630) );
  OAI21_X1 U24270 ( .B1(n26117), .B2(n9441), .A(n37640), .ZN(n5865) );
  AOI22_X1 U24271 ( .A1(N5086), .A2(n24246), .B1(N5053), .B2(n25899), .ZN(
        n37640) );
  OAI21_X1 U24272 ( .B1(n21576), .B2(n9567), .A(n37160), .ZN(n5831) );
  AOI22_X1 U24273 ( .A1(N4916), .A2(n267601), .B1(N4883), .B2(n24494), .ZN(
        n37160) );
  OAI21_X1 U24274 ( .B1(n21563), .B2(n9571), .A(n37170), .ZN(n5832) );
  AOI22_X1 U24275 ( .A1(N4915), .A2(n26012), .B1(N4882), .B2(n24748), .ZN(
        n37170) );
  OAI21_X1 U24276 ( .B1(n21568), .B2(n9575), .A(n37180), .ZN(n5833) );
  AOI22_X1 U24277 ( .A1(N4914), .A2(n24231), .B1(N4881), .B2(n25581), .ZN(
        n37180) );
  OAI21_X1 U24278 ( .B1(n26109), .B2(n9579), .A(n37190), .ZN(n5834) );
  AOI22_X1 U24279 ( .A1(N4913), .A2(n26017), .B1(N4880), .B2(n27222), .ZN(
        n37190) );
  OAI21_X1 U24280 ( .B1(n21559), .B2(n9583), .A(n37200), .ZN(n5835) );
  AOI22_X1 U24281 ( .A1(N4912), .A2(n26316), .B1(N4879), .B2(n25579), .ZN(
        n37200) );
  OAI21_X1 U24282 ( .B1(n21578), .B2(n9587), .A(n3721), .ZN(n5836) );
  AOI22_X1 U24283 ( .A1(N4911), .A2(n26032), .B1(N4878), .B2(n24751), .ZN(
        n3721) );
  OAI21_X1 U24284 ( .B1(n21565), .B2(n9591), .A(n3722), .ZN(n5837) );
  AOI22_X1 U24285 ( .A1(N4910), .A2(n21840), .B1(N4877), .B2(n25865), .ZN(
        n3722) );
  OAI21_X1 U24286 ( .B1(n21570), .B2(n9595), .A(n3723), .ZN(n5838) );
  AOI22_X1 U24287 ( .A1(N4909), .A2(n260701), .B1(N4876), .B2(n25861), .ZN(
        n3723) );
  OAI21_X1 U24288 ( .B1(n261101), .B2(n9599), .A(n3724), .ZN(n5839) );
  AOI22_X1 U24289 ( .A1(N4908), .A2(n26768), .B1(N4875), .B2(n24487), .ZN(
        n3724) );
  OAI21_X1 U24290 ( .B1(n21561), .B2(n9603), .A(n3725), .ZN(n5840) );
  AOI22_X1 U24291 ( .A1(N4907), .A2(n26015), .B1(N4874), .B2(n24756), .ZN(
        n3725) );
  OAI21_X1 U24292 ( .B1(n26126), .B2(n9981), .A(n3611), .ZN(n57660) );
  AOI22_X1 U24293 ( .A1(N4468), .A2(n267801), .B1(N4435), .B2(n24792), .ZN(
        n3611) );
  OAI21_X1 U24294 ( .B1(n26128), .B2(n9985), .A(n3612), .ZN(n57670) );
  AOI22_X1 U24295 ( .A1(N4467), .A2(n24237), .B1(N4434), .B2(n25895), .ZN(
        n3612) );
  OAI21_X1 U24296 ( .B1(n26122), .B2(n9989), .A(n3613), .ZN(n57680) );
  AOI22_X1 U24297 ( .A1(N4466), .A2(n21846), .B1(N4433), .B2(n25903), .ZN(
        n3613) );
  OAI21_X1 U24298 ( .B1(n26118), .B2(n9998), .A(n3615), .ZN(n57700) );
  AOI22_X1 U24299 ( .A1(N4464), .A2(n26038), .B1(N4431), .B2(n19210), .ZN(
        n3615) );
  OAI21_X1 U24300 ( .B1(n26119), .B2(n10089), .A(n3557), .ZN(n57260) );
  AOI22_X1 U24301 ( .A1(N4310), .A2(n21470), .B1(N4277), .B2(n25871), .ZN(
        n3557) );
  OAI21_X1 U24302 ( .B1(n26113), .B2(n10094), .A(n3558), .ZN(n57270) );
  AOI22_X1 U24303 ( .A1(N4309), .A2(n26063), .B1(N4276), .B2(n25870), .ZN(
        n3558) );
  OAI21_X1 U24304 ( .B1(n26115), .B2(n10099), .A(n3559), .ZN(n57280) );
  AOI22_X1 U24305 ( .A1(N4308), .A2(n24250), .B1(N4275), .B2(n25871), .ZN(
        n3559) );
  OAI21_X1 U24306 ( .B1(n21555), .B2(n10104), .A(n3560), .ZN(n57290) );
  AOI22_X1 U24307 ( .A1(N4307), .A2(n23163), .B1(N4274), .B2(n25867), .ZN(
        n3560) );
  OAI21_X1 U24308 ( .B1(n26111), .B2(n10109), .A(n3561), .ZN(n57300) );
  AOI22_X1 U24309 ( .A1(N4306), .A2(n23181), .B1(N4273), .B2(n25877), .ZN(
        n3561) );
  OAI21_X1 U24310 ( .B1(n21587), .B2(n10514), .A(n3449), .ZN(n56560) );
  AOI22_X1 U24311 ( .A1(N3880), .A2(n26314), .B1(N3847), .B2(n19211), .ZN(
        n3449) );
  OAI21_X1 U24312 ( .B1(n21591), .B2(n10519), .A(n3450), .ZN(n56570) );
  AOI22_X1 U24313 ( .A1(N3879), .A2(n21467), .B1(N3846), .B2(n24786), .ZN(
        n3450) );
  OAI21_X1 U24314 ( .B1(n21579), .B2(n10524), .A(n3451), .ZN(n5658) );
  AOI22_X1 U24315 ( .A1(N3878), .A2(n21473), .B1(N3845), .B2(n21273), .ZN(
        n3451) );
  OAI21_X1 U24316 ( .B1(n21585), .B2(n10529), .A(n3452), .ZN(n5659) );
  AOI22_X1 U24317 ( .A1(N3877), .A2(n22872), .B1(N3844), .B2(n21276), .ZN(
        n3452) );
  OAI21_X1 U24318 ( .B1(n21571), .B2(n10534), .A(n34530), .ZN(n5660) );
  AOI22_X1 U24319 ( .A1(N3876), .A2(n26308), .B1(N3843), .B2(n21271), .ZN(
        n34530) );
  OAI21_X1 U24320 ( .B1(n21589), .B2(n10539), .A(n34540), .ZN(n5661) );
  AOI22_X1 U24321 ( .A1(N3875), .A2(n21481), .B1(N3842), .B2(n22885), .ZN(
        n34540) );
  OAI21_X1 U24322 ( .B1(n21593), .B2(n10544), .A(n34550), .ZN(n5662) );
  AOI22_X1 U24323 ( .A1(N3874), .A2(n23154), .B1(N3841), .B2(n27201), .ZN(
        n34550) );
  OAI21_X1 U24324 ( .B1(n21581), .B2(n10549), .A(n34560), .ZN(n5663) );
  AOI22_X1 U24325 ( .A1(N3873), .A2(n23169), .B1(N3840), .B2(n27199), .ZN(
        n34560) );
  OAI21_X1 U24326 ( .B1(n21573), .B2(n10558), .A(n34580), .ZN(n5665) );
  AOI22_X1 U24327 ( .A1(N3871), .A2(n21460), .B1(N3838), .B2(n25586), .ZN(
        n34580) );
  OAI21_X1 U24328 ( .B1(n261201), .B2(n10700), .A(n3407), .ZN(n5631) );
  AOI22_X1 U24329 ( .A1(N3704), .A2(n26776), .B1(N3671), .B2(n19245), .ZN(
        n3407) );
  OAI21_X1 U24330 ( .B1(n26114), .B2(n10704), .A(n3408), .ZN(n5632) );
  AOI22_X1 U24331 ( .A1(N3703), .A2(n22836), .B1(N3670), .B2(n24756), .ZN(
        n3408) );
  OAI21_X1 U24332 ( .B1(n26116), .B2(n10708), .A(n3409), .ZN(n5633) );
  AOI22_X1 U24333 ( .A1(N3702), .A2(n21854), .B1(N3669), .B2(n25869), .ZN(
        n3409) );
  OAI21_X1 U24334 ( .B1(n26112), .B2(n10717), .A(n3411), .ZN(n5635) );
  AOI22_X1 U24335 ( .A1(N3700), .A2(n26064), .B1(N3667), .B2(n19207), .ZN(
        n3411) );
  OAI21_X1 U24336 ( .B1(n21575), .B2(n11217), .A(n3242), .ZN(n55210) );
  AOI22_X1 U24337 ( .A1(N3123), .A2(n26318), .B1(N3090), .B2(n21254), .ZN(
        n3242) );
  OAI21_X1 U24338 ( .B1(n21563), .B2(n11222), .A(n3243), .ZN(n55220) );
  AOI22_X1 U24339 ( .A1(N3122), .A2(n26016), .B1(N3089), .B2(n20544), .ZN(
        n3243) );
  OAI21_X1 U24340 ( .B1(n21567), .B2(n11227), .A(n3244), .ZN(n55230) );
  AOI22_X1 U24341 ( .A1(N3121), .A2(n26033), .B1(N3088), .B2(n21261), .ZN(
        n3244) );
  OAI21_X1 U24342 ( .B1(n21557), .B2(n11232), .A(n3245), .ZN(n55240) );
  AOI22_X1 U24343 ( .A1(N3120), .A2(n23158), .B1(N3087), .B2(n21253), .ZN(
        n3245) );
  OAI21_X1 U24344 ( .B1(n21559), .B2(n11237), .A(n3246), .ZN(n55250) );
  AOI22_X1 U24345 ( .A1(N3119), .A2(n26310), .B1(N3086), .B2(n24493), .ZN(
        n3246) );
  OAI21_X1 U24346 ( .B1(n21577), .B2(n11242), .A(n3247), .ZN(n55260) );
  AOI22_X1 U24347 ( .A1(N3118), .A2(n21497), .B1(N3085), .B2(n24748), .ZN(
        n3247) );
  OAI21_X1 U24348 ( .B1(n21565), .B2(n11247), .A(n3248), .ZN(n55270) );
  AOI22_X1 U24349 ( .A1(N3117), .A2(n19254), .B1(N3084), .B2(n24492), .ZN(
        n3248) );
  OAI21_X1 U24350 ( .B1(n21569), .B2(n11252), .A(n3249), .ZN(n5528) );
  AOI22_X1 U24351 ( .A1(N3116), .A2(n23182), .B1(N3083), .B2(n27222), .ZN(
        n3249) );
  OAI21_X1 U24352 ( .B1(n21561), .B2(n11261), .A(n3251), .ZN(n5530) );
  AOI22_X1 U24353 ( .A1(N3114), .A2(n26011), .B1(N3081), .B2(n21251), .ZN(
        n3251) );
  NAND2_X1 U24354 ( .A1(n4991), .A2(n4992), .ZN(mul_outcome[40]) );
  AOI221_X1 U24355 ( .B1(n21549), .B2(n17861), .C1(n25916), .C2(n17849), .A(
        n49940), .ZN(n4991) );
  AOI221_X1 U24356 ( .B1(n21553), .B2(n17885), .C1(n21540), .C2(n17873), .A(
        n4993), .ZN(n4992) );
  OAI22_X1 U24357 ( .A1(n2065), .A2(n20480), .B1(n2044), .B2(n20484), .ZN(
        n49940) );
  OAI21_X1 U24358 ( .B1(n21453), .B2(n905), .A(n4500), .ZN(n6341) );
  AOI22_X1 U24359 ( .A1(N7822), .A2(n257101), .B1(N7789), .B2(n24480), .ZN(
        n4500) );
  OAI21_X1 U24360 ( .B1(n21454), .B2(n909), .A(n4501), .ZN(n6342) );
  AOI22_X1 U24361 ( .A1(N7821), .A2(n25706), .B1(N7788), .B2(n26140), .ZN(
        n4501) );
  OAI21_X1 U24362 ( .B1(n259801), .B2(n913), .A(n4502), .ZN(n6343) );
  AOI22_X1 U24363 ( .A1(N7820), .A2(n25696), .B1(N7787), .B2(n24474), .ZN(
        n4502) );
  OAI21_X1 U24364 ( .B1(n20878), .B2(n917), .A(n4503), .ZN(n6344) );
  AOI22_X1 U24365 ( .A1(N7819), .A2(n25714), .B1(N7786), .B2(n21611), .ZN(
        n4503) );
  OAI21_X1 U24366 ( .B1(n24516), .B2(n921), .A(n4504), .ZN(n6345) );
  AOI22_X1 U24367 ( .A1(N7818), .A2(n25728), .B1(N7785), .B2(n23276), .ZN(
        n4504) );
  OAI21_X1 U24368 ( .B1(n25981), .B2(n925), .A(n4505), .ZN(n6346) );
  AOI22_X1 U24369 ( .A1(N7817), .A2(n25735), .B1(N7784), .B2(n27148), .ZN(
        n4505) );
  OAI21_X1 U24370 ( .B1(n25984), .B2(n929), .A(n4506), .ZN(n6347) );
  AOI22_X1 U24371 ( .A1(N7816), .A2(n25527), .B1(N7783), .B2(n21616), .ZN(
        n4506) );
  OAI21_X1 U24372 ( .B1(n25979), .B2(n933), .A(n4507), .ZN(n6348) );
  AOI22_X1 U24373 ( .A1(N7815), .A2(n25715), .B1(N7782), .B2(n17095), .ZN(
        n4507) );
  OAI21_X1 U24374 ( .B1(n24514), .B2(n937), .A(n4508), .ZN(n6349) );
  AOI22_X1 U24375 ( .A1(N7814), .A2(n25718), .B1(N7781), .B2(n27149), .ZN(
        n4508) );
  OAI21_X1 U24376 ( .B1(n24517), .B2(n941), .A(n45090), .ZN(n63500) );
  AOI22_X1 U24377 ( .A1(N7813), .A2(n25711), .B1(N7780), .B2(n21619), .ZN(
        n45090) );
  OAI21_X1 U24378 ( .B1(n25982), .B2(n945), .A(n4510), .ZN(n63510) );
  AOI22_X1 U24379 ( .A1(N7812), .A2(n25707), .B1(N7779), .B2(n21613), .ZN(
        n4510) );
  OAI21_X1 U24380 ( .B1(n25985), .B2(n1920), .A(n4511), .ZN(n63520) );
  AOI22_X1 U24381 ( .A1(N7811), .A2(n25697), .B1(N7778), .B2(n27149), .ZN(
        n4511) );
  OAI21_X1 U24382 ( .B1(n23117), .B2(n1924), .A(n4512), .ZN(n63530) );
  AOI22_X1 U24383 ( .A1(N7810), .A2(n25712), .B1(N7777), .B2(n24479), .ZN(
        n4512) );
  OAI21_X1 U24384 ( .B1(n24513), .B2(n2207), .A(n45130), .ZN(n63540) );
  AOI22_X1 U24385 ( .A1(N7809), .A2(n25729), .B1(N7776), .B2(n27150), .ZN(
        n45130) );
  OAI21_X1 U24386 ( .B1(n25979), .B2(n2287), .A(n45140), .ZN(n63550) );
  AOI22_X1 U24387 ( .A1(N7808), .A2(n25732), .B1(N7775), .B2(n21614), .ZN(
        n45140) );
  OAI21_X1 U24388 ( .B1(n25983), .B2(n7524), .A(n4330), .ZN(n62360) );
  AOI22_X1 U24389 ( .A1(N7236), .A2(n25713), .B1(N7203), .B2(n26139), .ZN(
        n4330) );
  OAI21_X1 U24390 ( .B1(n25986), .B2(n75280), .A(n4331), .ZN(n62370) );
  AOI22_X1 U24391 ( .A1(N7235), .A2(n257301), .B1(N7202), .B2(n20564), .ZN(
        n4331) );
  OAI21_X1 U24392 ( .B1(n23118), .B2(n75320), .A(n4332), .ZN(n62380) );
  AOI22_X1 U24393 ( .A1(N7234), .A2(n25733), .B1(N7201), .B2(n24480), .ZN(
        n4332) );
  OAI21_X1 U24394 ( .B1(n24516), .B2(n75360), .A(n4333), .ZN(n62390) );
  AOI22_X1 U24395 ( .A1(N7233), .A2(n21160), .B1(N7200), .B2(n17095), .ZN(
        n4333) );
  OAI21_X1 U24396 ( .B1(n23118), .B2(n75400), .A(n4334), .ZN(n62400) );
  AOI22_X1 U24397 ( .A1(N7232), .A2(n25719), .B1(N7199), .B2(n26140), .ZN(
        n4334) );
  OAI21_X1 U24398 ( .B1(n21452), .B2(n7544), .A(n4335), .ZN(n62410) );
  AOI22_X1 U24399 ( .A1(N7231), .A2(n25708), .B1(N7198), .B2(n17075), .ZN(
        n4335) );
  OAI21_X1 U24400 ( .B1(n21455), .B2(n7548), .A(n4336), .ZN(n62420) );
  AOI22_X1 U24401 ( .A1(N7230), .A2(n25704), .B1(N7197), .B2(n20566), .ZN(
        n4336) );
  OAI21_X1 U24402 ( .B1(n23117), .B2(n7552), .A(n4337), .ZN(n62430) );
  AOI22_X1 U24403 ( .A1(N7229), .A2(n25705), .B1(N7196), .B2(n21612), .ZN(
        n4337) );
  OAI21_X1 U24404 ( .B1(n25080), .B2(n7556), .A(n4338), .ZN(n6244) );
  AOI22_X1 U24405 ( .A1(N7228), .A2(n25698), .B1(N7195), .B2(n24479), .ZN(
        n4338) );
  OAI21_X1 U24406 ( .B1(n23120), .B2(n7560), .A(n4339), .ZN(n6245) );
  AOI22_X1 U24407 ( .A1(N7227), .A2(n25714), .B1(N7194), .B2(n23274), .ZN(
        n4339) );
  OAI21_X1 U24408 ( .B1(n25981), .B2(n75640), .A(n4340), .ZN(n6246) );
  AOI22_X1 U24409 ( .A1(N7226), .A2(n25731), .B1(N7193), .B2(n24764), .ZN(
        n4340) );
  OAI21_X1 U24410 ( .B1(n25984), .B2(n75680), .A(n4341), .ZN(n6247) );
  AOI22_X1 U24411 ( .A1(N7225), .A2(n25734), .B1(N7192), .B2(n23273), .ZN(
        n4341) );
  OAI21_X1 U24412 ( .B1(n23119), .B2(n75720), .A(n43420), .ZN(n6248) );
  AOI22_X1 U24413 ( .A1(N7224), .A2(n19182), .B1(N7191), .B2(n21618), .ZN(
        n43420) );
  OAI21_X1 U24414 ( .B1(n24515), .B2(n75760), .A(n43430), .ZN(n6249) );
  AOI22_X1 U24415 ( .A1(N7223), .A2(n25716), .B1(N7190), .B2(n26143), .ZN(
        n43430) );
  OAI21_X1 U24416 ( .B1(n20878), .B2(n75810), .A(n43440), .ZN(n6250) );
  AOI22_X1 U24417 ( .A1(N7222), .A2(n25699), .B1(N7189), .B2(n24764), .ZN(
        n43440) );
  OAI21_X1 U24418 ( .B1(n25982), .B2(n8033), .A(n4172), .ZN(n6131) );
  AOI22_X1 U24419 ( .A1(N6614), .A2(n25527), .B1(N6581), .B2(n23273), .ZN(
        n4172) );
  OAI21_X1 U24420 ( .B1(n25985), .B2(n8038), .A(n4173), .ZN(n6132) );
  AOI22_X1 U24421 ( .A1(N6613), .A2(n25717), .B1(N6580), .B2(n23276), .ZN(
        n4173) );
  OAI21_X1 U24422 ( .B1(n23120), .B2(n8043), .A(n41740), .ZN(n6133) );
  AOI22_X1 U24423 ( .A1(N6612), .A2(n25709), .B1(N6579), .B2(n21615), .ZN(
        n41740) );
  OAI21_X1 U24424 ( .B1(n24518), .B2(n8048), .A(n41750), .ZN(n6134) );
  AOI22_X1 U24425 ( .A1(N6611), .A2(n25706), .B1(N6578), .B2(n21618), .ZN(
        n41750) );
  OAI21_X1 U24426 ( .B1(n24514), .B2(n8053), .A(n41760), .ZN(n6135) );
  AOI22_X1 U24427 ( .A1(N6610), .A2(n25698), .B1(N6577), .B2(n23274), .ZN(
        n41760) );
  OAI21_X1 U24428 ( .B1(n25983), .B2(n8058), .A(n41770), .ZN(n6136) );
  AOI22_X1 U24429 ( .A1(N6609), .A2(n25718), .B1(N6576), .B2(n23277), .ZN(
        n41770) );
  OAI21_X1 U24430 ( .B1(n25986), .B2(n8063), .A(n41780), .ZN(n6137) );
  AOI22_X1 U24431 ( .A1(N6608), .A2(n25715), .B1(N6575), .B2(n21613), .ZN(
        n41780) );
  OAI21_X1 U24432 ( .B1(n25080), .B2(n8068), .A(n41790), .ZN(n6138) );
  AOI22_X1 U24433 ( .A1(N6607), .A2(n25731), .B1(N6574), .B2(n24474), .ZN(
        n41790) );
  OAI21_X1 U24434 ( .B1(n24517), .B2(n8073), .A(n41800), .ZN(n6139) );
  AOI22_X1 U24435 ( .A1(N6606), .A2(n25735), .B1(N6573), .B2(n26139), .ZN(
        n41800) );
  OAI21_X1 U24436 ( .B1(n24515), .B2(n8078), .A(n41810), .ZN(n6140) );
  AOI22_X1 U24437 ( .A1(N6605), .A2(n21159), .B1(N6572), .B2(n23277), .ZN(
        n41810) );
  OAI21_X1 U24438 ( .B1(n21452), .B2(n8083), .A(n41820), .ZN(n6141) );
  AOI22_X1 U24439 ( .A1(N6604), .A2(n25719), .B1(N6571), .B2(n20563), .ZN(
        n41820) );
  OAI21_X1 U24440 ( .B1(n21454), .B2(n8088), .A(n41830), .ZN(n6142) );
  AOI22_X1 U24441 ( .A1(N6603), .A2(n257101), .B1(N6570), .B2(n17075), .ZN(
        n41830) );
  OAI21_X1 U24442 ( .B1(n23119), .B2(n8093), .A(n41840), .ZN(n6143) );
  AOI22_X1 U24443 ( .A1(N6602), .A2(n25707), .B1(N6569), .B2(n24473), .ZN(
        n41840) );
  OAI21_X1 U24444 ( .B1(n259801), .B2(n8098), .A(n41850), .ZN(n6144) );
  AOI22_X1 U24445 ( .A1(N6601), .A2(n25711), .B1(N6568), .B2(n20565), .ZN(
        n41850) );
  OAI21_X1 U24446 ( .B1(n24518), .B2(n8102), .A(n41860), .ZN(n6145) );
  AOI22_X1 U24447 ( .A1(N6600), .A2(n25699), .B1(N6567), .B2(n26143), .ZN(
        n41860) );
  OAI21_X1 U24448 ( .B1(n21449), .B2(n10409), .A(n34660), .ZN(n5666) );
  AOI22_X1 U24449 ( .A1(N3974), .A2(n256801), .B1(N3941), .B2(n24483), .ZN(
        n34660) );
  OAI21_X1 U24450 ( .B1(n21450), .B2(n10414), .A(n34670), .ZN(n5667) );
  AOI22_X1 U24451 ( .A1(N3973), .A2(n25693), .B1(N3940), .B2(n26136), .ZN(
        n34670) );
  OAI21_X1 U24452 ( .B1(n25972), .B2(n10419), .A(n34680), .ZN(n5668) );
  AOI22_X1 U24453 ( .A1(N3972), .A2(n25683), .B1(N3939), .B2(n24477), .ZN(
        n34680) );
  OAI21_X1 U24454 ( .B1(n20883), .B2(n10424), .A(n34690), .ZN(n5669) );
  AOI22_X1 U24455 ( .A1(N3971), .A2(n25702), .B1(N3938), .B2(n21607), .ZN(
        n34690) );
  OAI21_X1 U24456 ( .B1(n24523), .B2(n10429), .A(n34700), .ZN(n5670) );
  AOI22_X1 U24457 ( .A1(N3970), .A2(n257201), .B1(N3937), .B2(n23268), .ZN(
        n34700) );
  OAI21_X1 U24458 ( .B1(n25973), .B2(n10434), .A(n34710), .ZN(n5671) );
  AOI22_X1 U24459 ( .A1(N3969), .A2(n25727), .B1(N3936), .B2(n27270), .ZN(
        n34710) );
  OAI21_X1 U24460 ( .B1(n25975), .B2(n10439), .A(n34720), .ZN(n5672) );
  AOI22_X1 U24461 ( .A1(N3968), .A2(n25523), .B1(N3935), .B2(n21620), .ZN(
        n34720) );
  OAI21_X1 U24462 ( .B1(n25971), .B2(n10444), .A(n34730), .ZN(n5673) );
  AOI22_X1 U24463 ( .A1(N3967), .A2(n25703), .B1(N3934), .B2(n17096), .ZN(
        n34730) );
  OAI21_X1 U24464 ( .B1(n24521), .B2(n10449), .A(n3474), .ZN(n5674) );
  AOI22_X1 U24465 ( .A1(N3966), .A2(n25689), .B1(N3933), .B2(n27271), .ZN(
        n3474) );
  OAI21_X1 U24466 ( .B1(n24524), .B2(n10454), .A(n3475), .ZN(n56750) );
  AOI22_X1 U24467 ( .A1(N3965), .A2(n25681), .B1(N3932), .B2(n21623), .ZN(
        n3475) );
  OAI21_X1 U24468 ( .B1(n17079), .B2(n10459), .A(n3476), .ZN(n56760) );
  AOI22_X1 U24469 ( .A1(N3964), .A2(n25694), .B1(N3931), .B2(n21609), .ZN(
        n3476) );
  OAI21_X1 U24470 ( .B1(n25976), .B2(n10464), .A(n3477), .ZN(n56770) );
  AOI22_X1 U24471 ( .A1(N3963), .A2(n25684), .B1(N3930), .B2(n27271), .ZN(
        n3477) );
  OAI21_X1 U24472 ( .B1(n23109), .B2(n10469), .A(n3478), .ZN(n56780) );
  AOI22_X1 U24473 ( .A1(N3962), .A2(n257001), .B1(N3929), .B2(n24482), .ZN(
        n3478) );
  OAI21_X1 U24474 ( .B1(n24520), .B2(n10474), .A(n3479), .ZN(n56790) );
  AOI22_X1 U24475 ( .A1(N3961), .A2(n25721), .B1(N3928), .B2(n27272), .ZN(
        n3479) );
  OAI21_X1 U24476 ( .B1(n25971), .B2(n10478), .A(n3480), .ZN(n56800) );
  AOI22_X1 U24477 ( .A1(N3960), .A2(n25724), .B1(N3927), .B2(n21610), .ZN(
        n3480) );
  OAI21_X1 U24478 ( .B1(n25974), .B2(n10965), .A(n3309), .ZN(n55610) );
  AOI22_X1 U24479 ( .A1(N3378), .A2(n25701), .B1(N3345), .B2(n26135), .ZN(
        n3309) );
  OAI21_X1 U24480 ( .B1(n25977), .B2(n10970), .A(n3310), .ZN(n55620) );
  AOI22_X1 U24481 ( .A1(N3377), .A2(n25722), .B1(N3344), .B2(n17096), .ZN(
        n3310) );
  OAI21_X1 U24482 ( .B1(n23110), .B2(n10975), .A(n3311), .ZN(n55630) );
  AOI22_X1 U24483 ( .A1(N3376), .A2(n25725), .B1(N3343), .B2(n24483), .ZN(
        n3311) );
  OAI21_X1 U24484 ( .B1(n24523), .B2(n10980), .A(n3312), .ZN(n55640) );
  AOI22_X1 U24485 ( .A1(N3375), .A2(n21154), .B1(N3342), .B2(n20558), .ZN(
        n3312) );
  OAI21_X1 U24486 ( .B1(n23110), .B2(n10985), .A(n3313), .ZN(n55650) );
  AOI22_X1 U24487 ( .A1(N3374), .A2(n256901), .B1(N3341), .B2(n26136), .ZN(
        n3313) );
  OAI21_X1 U24488 ( .B1(n21448), .B2(n10990), .A(n3314), .ZN(n55660) );
  AOI22_X1 U24489 ( .A1(N3373), .A2(n25678), .B1(N3340), .B2(n17074), .ZN(
        n3314) );
  OAI21_X1 U24490 ( .B1(n21451), .B2(n10995), .A(n3315), .ZN(n55670) );
  AOI22_X1 U24491 ( .A1(N3372), .A2(n25691), .B1(N3339), .B2(n24762), .ZN(
        n3315) );
  OAI21_X1 U24492 ( .B1(n23109), .B2(n11000), .A(n3316), .ZN(n55680) );
  AOI22_X1 U24493 ( .A1(N3371), .A2(n25692), .B1(N3338), .B2(n21608), .ZN(
        n3316) );
  OAI21_X1 U24494 ( .B1(n25084), .B2(n11005), .A(n3317), .ZN(n5569) );
  AOI22_X1 U24495 ( .A1(N3370), .A2(n25685), .B1(N3337), .B2(n24482), .ZN(
        n3317) );
  OAI21_X1 U24496 ( .B1(n23112), .B2(n11010), .A(n3318), .ZN(n5570) );
  AOI22_X1 U24497 ( .A1(N3369), .A2(n25702), .B1(N3336), .B2(n23265), .ZN(
        n3318) );
  OAI21_X1 U24498 ( .B1(n25973), .B2(n11015), .A(n3319), .ZN(n5571) );
  AOI22_X1 U24499 ( .A1(N3368), .A2(n25723), .B1(N3335), .B2(n20561), .ZN(
        n3319) );
  OAI21_X1 U24500 ( .B1(n25975), .B2(n11020), .A(n3320), .ZN(n5572) );
  AOI22_X1 U24501 ( .A1(N3367), .A2(n25726), .B1(N3334), .B2(n23266), .ZN(
        n3320) );
  OAI21_X1 U24502 ( .B1(n23111), .B2(n11025), .A(n3321), .ZN(n5573) );
  AOI22_X1 U24503 ( .A1(N3366), .A2(n19180), .B1(N3333), .B2(n21623), .ZN(
        n3321) );
  OAI21_X1 U24504 ( .B1(n24522), .B2(n11030), .A(n3322), .ZN(n5574) );
  AOI22_X1 U24505 ( .A1(N3365), .A2(n25687), .B1(N3332), .B2(n26144), .ZN(
        n3322) );
  OAI21_X1 U24506 ( .B1(n20882), .B2(n11034), .A(n3323), .ZN(n5575) );
  AOI22_X1 U24507 ( .A1(N3364), .A2(n25686), .B1(N3331), .B2(n20560), .ZN(
        n3323) );
  OAI21_X1 U24508 ( .B1(n17079), .B2(n11499), .A(n3137), .ZN(n5456) );
  AOI22_X1 U24509 ( .A1(N2780), .A2(n25523), .B1(N2747), .B2(n23265), .ZN(
        n3137) );
  OAI21_X1 U24510 ( .B1(n25976), .B2(n11504), .A(n3138), .ZN(n5457) );
  AOI22_X1 U24511 ( .A1(N2779), .A2(n25688), .B1(N2746), .B2(n23269), .ZN(
        n3138) );
  OAI21_X1 U24512 ( .B1(n23112), .B2(n11509), .A(n3139), .ZN(n5458) );
  AOI22_X1 U24513 ( .A1(N2778), .A2(n25679), .B1(N2745), .B2(n21621), .ZN(
        n3139) );
  OAI21_X1 U24514 ( .B1(n24525), .B2(n11514), .A(n3140), .ZN(n5459) );
  AOI22_X1 U24515 ( .A1(N2777), .A2(n25693), .B1(N2744), .B2(n21624), .ZN(
        n3140) );
  OAI21_X1 U24516 ( .B1(n24521), .B2(n11519), .A(n3141), .ZN(n5460) );
  AOI22_X1 U24517 ( .A1(N2776), .A2(n25685), .B1(N2743), .B2(n23266), .ZN(
        n3141) );
  OAI21_X1 U24518 ( .B1(n25974), .B2(n11524), .A(n3142), .ZN(n5461) );
  AOI22_X1 U24519 ( .A1(N2775), .A2(n25689), .B1(N2742), .B2(n23269), .ZN(
        n3142) );
  OAI21_X1 U24520 ( .B1(n25977), .B2(n11529), .A(n3143), .ZN(n5462) );
  AOI22_X1 U24521 ( .A1(N2774), .A2(n25703), .B1(N2741), .B2(n21609), .ZN(
        n3143) );
  OAI21_X1 U24522 ( .B1(n25084), .B2(n11534), .A(n3144), .ZN(n5463) );
  AOI22_X1 U24523 ( .A1(N2773), .A2(n25723), .B1(N2740), .B2(n24476), .ZN(
        n3144) );
  OAI21_X1 U24524 ( .B1(n24524), .B2(n11539), .A(n3145), .ZN(n5464) );
  AOI22_X1 U24525 ( .A1(N2772), .A2(n25727), .B1(N2739), .B2(n26135), .ZN(
        n3145) );
  OAI21_X1 U24526 ( .B1(n24522), .B2(n11544), .A(n3146), .ZN(n5465) );
  AOI22_X1 U24527 ( .A1(N2771), .A2(n21153), .B1(N2738), .B2(n23268), .ZN(
        n3146) );
  OAI21_X1 U24528 ( .B1(n21448), .B2(n11549), .A(n3147), .ZN(n5466) );
  AOI22_X1 U24529 ( .A1(N2770), .A2(n256901), .B1(N2737), .B2(n20559), .ZN(
        n3147) );
  OAI21_X1 U24530 ( .B1(n21450), .B2(n11554), .A(n3148), .ZN(n5467) );
  AOI22_X1 U24531 ( .A1(N2769), .A2(n256801), .B1(N2736), .B2(n17074), .ZN(
        n3148) );
  OAI21_X1 U24532 ( .B1(n23111), .B2(n11559), .A(n3149), .ZN(n5468) );
  AOI22_X1 U24533 ( .A1(N2768), .A2(n25694), .B1(N2735), .B2(n24477), .ZN(
        n3149) );
  OAI21_X1 U24534 ( .B1(n25972), .B2(n11564), .A(n3150), .ZN(n5469) );
  AOI22_X1 U24535 ( .A1(N2767), .A2(n25681), .B1(N2734), .B2(n24762), .ZN(
        n3150) );
  OAI21_X1 U24536 ( .B1(n24525), .B2(n11568), .A(n3151), .ZN(n5470) );
  AOI22_X1 U24537 ( .A1(N2766), .A2(n25686), .B1(N2733), .B2(n26144), .ZN(
        n3151) );
  OR2_X1 U24538 ( .A1(n26970), .A2(upper_bound[3]), .ZN(n53950) );
  OR2_X1 U24539 ( .A1(n26972), .A2(n26971), .ZN(n26970) );
  NAND2_X1 U24540 ( .A1(n52130), .A2(n5214), .ZN(mul_outcome[144]) );
  AOI221_X1 U24541 ( .B1(n26402), .B2(n17395), .C1(n26496), .C2(n17371), .A(
        n27735), .ZN(n52130) );
  AOI221_X1 U24542 ( .B1(n21361), .B2(n17455), .C1(n27035), .C2(n17443), .A(
        n27751), .ZN(n5214) );
  INV_X1 U24543 ( .A(n5216), .ZN(n27735) );
  NAND2_X1 U24544 ( .A1(n5114), .A2(n5115), .ZN(mul_outcome[165]) );
  AOI221_X1 U24545 ( .B1(n26502), .B2(n17287), .C1(n25330), .C2(n17275), .A(
        n27729), .ZN(n5114) );
  AOI221_X1 U24546 ( .B1(n21389), .B2(n17359), .C1(n26058), .C2(n17347), .A(
        n277701), .ZN(n5115) );
  INV_X1 U24547 ( .A(n5117), .ZN(n27729) );
  NAND2_X1 U24548 ( .A1(n52210), .A2(n52220), .ZN(mul_outcome[142]) );
  AOI221_X1 U24549 ( .B1(n21975), .B2(n17399), .C1(n26240), .C2(n17375), .A(
        n27737), .ZN(n52210) );
  AOI221_X1 U24550 ( .B1(n21363), .B2(n17459), .C1(n27033), .C2(n17447), .A(
        n27753), .ZN(n52220) );
  INV_X1 U24551 ( .A(n52240), .ZN(n27737) );
  NAND2_X1 U24552 ( .A1(n5122), .A2(n5123), .ZN(mul_outcome[163]) );
  AOI221_X1 U24553 ( .B1(n26241), .B2(n17291), .C1(n24159), .C2(n17279), .A(
        n27731), .ZN(n5122) );
  AOI221_X1 U24554 ( .B1(n21375), .B2(n17363), .C1(n26059), .C2(n17351), .A(
        n27772), .ZN(n5123) );
  INV_X1 U24555 ( .A(n5125), .ZN(n27731) );
  NAND2_X1 U24556 ( .A1(n52170), .A2(n52180), .ZN(mul_outcome[143]) );
  AOI221_X1 U24557 ( .B1(n26395), .B2(n17397), .C1(n22419), .C2(n17373), .A(
        n27736), .ZN(n52170) );
  AOI221_X1 U24558 ( .B1(n21354), .B2(n17457), .C1(n27034), .C2(n17445), .A(
        n27752), .ZN(n52180) );
  INV_X1 U24559 ( .A(n52200), .ZN(n27736) );
  NAND2_X1 U24560 ( .A1(n5209), .A2(n5210), .ZN(mul_outcome[145]) );
  AOI221_X1 U24561 ( .B1(n24397), .B2(n17393), .C1(n24312), .C2(n17369), .A(
        n27734), .ZN(n5209) );
  AOI221_X1 U24562 ( .B1(n21365), .B2(n17453), .C1(n27036), .C2(n17441), .A(
        n277501), .ZN(n5210) );
  INV_X1 U24563 ( .A(n5212), .ZN(n27734) );
  NAND2_X1 U24564 ( .A1(n5110), .A2(n5111), .ZN(mul_outcome[166]) );
  AOI221_X1 U24565 ( .B1(n26243), .B2(n17285), .C1(n26707), .C2(n17273), .A(
        n27728), .ZN(n5110) );
  AOI221_X1 U24566 ( .B1(n21377), .B2(n17357), .C1(n24262), .C2(n17345), .A(
        n27769), .ZN(n5111) );
  INV_X1 U24567 ( .A(n5113), .ZN(n27728) );
  OR2_X1 U24568 ( .A1(n546), .A2(sub_127_aco_carry[4]), .ZN(
        sub_127_aco_carry[5]) );
  XOR2_X1 U24569 ( .A(n458), .B(n26969), .Z(n26971) );
  AOI221_X1 U24570 ( .B1(n27095), .B2(matrix_mul_2D_2__4__12_), .C1(n21359), 
        .C2(matrix_mul_2D_2__5__12_), .A(n4926), .ZN(n4925) );
  OAI22_X1 U24571 ( .A1(n2228), .A2(n24966), .B1(n2213), .B2(n22457), .ZN(
        n4926) );
  AOI221_X1 U24572 ( .B1(n27096), .B2(matrix_mul_2D_2__4__13_), .C1(n19231), 
        .C2(matrix_mul_2D_2__5__13_), .A(n49220), .ZN(n49210) );
  OAI22_X1 U24573 ( .A1(n2227), .A2(n25093), .B1(n2212), .B2(n23679), .ZN(
        n49220) );
  AOI221_X1 U24574 ( .B1(n27097), .B2(matrix_mul_2D_2__4__14_), .C1(n21351), 
        .C2(matrix_mul_2D_2__5__14_), .A(n49180), .ZN(n49170) );
  OAI22_X1 U24575 ( .A1(n2226), .A2(n25347), .B1(n2211), .B2(n22504), .ZN(
        n49180) );
  INV_X1 U24576 ( .A(n53140), .ZN(n27776) );
  AOI22_X1 U24577 ( .A1(n17491), .A2(n23970), .B1(n17503), .B2(n25519), .ZN(
        n53140) );
  INV_X1 U24578 ( .A(n53100), .ZN(n27775) );
  AOI22_X1 U24579 ( .A1(n17489), .A2(n23978), .B1(n17501), .B2(n22535), .ZN(
        n53100) );
  INV_X1 U24580 ( .A(n5116), .ZN(n277701) );
  AOI22_X1 U24581 ( .A1(n17323), .A2(n19312), .B1(n17335), .B2(n24856), .ZN(
        n5116) );
  INV_X1 U24582 ( .A(n5112), .ZN(n27769) );
  AOI22_X1 U24583 ( .A1(n17321), .A2(n22678), .B1(n17333), .B2(n26588), .ZN(
        n5112) );
  INV_X1 U24584 ( .A(n5303), .ZN(n27774) );
  AOI22_X1 U24585 ( .A1(n17487), .A2(n25366), .B1(n17499), .B2(n26586), .ZN(
        n5303) );
  INV_X1 U24586 ( .A(n53180), .ZN(n27777) );
  AOI22_X1 U24587 ( .A1(n17493), .A2(n19064), .B1(n17505), .B2(n23729), .ZN(
        n53180) );
  INV_X1 U24588 ( .A(n5322), .ZN(n27778) );
  AOI22_X1 U24589 ( .A1(n17495), .A2(n26624), .B1(n17507), .B2(n26587), .ZN(
        n5322) );
  INV_X1 U24590 ( .A(n5326), .ZN(n27779) );
  AOI22_X1 U24591 ( .A1(n17497), .A2(n25025), .B1(n17509), .B2(n20862), .ZN(
        n5326) );
  INV_X1 U24592 ( .A(n5108), .ZN(n27768) );
  AOI22_X1 U24593 ( .A1(n17319), .A2(n23979), .B1(n17331), .B2(n22539), .ZN(
        n5108) );
  INV_X1 U24594 ( .A(n5120), .ZN(n27771) );
  AOI22_X1 U24595 ( .A1(n17325), .A2(n23981), .B1(n17337), .B2(n22538), .ZN(
        n5120) );
  INV_X1 U24596 ( .A(n5124), .ZN(n27772) );
  AOI22_X1 U24597 ( .A1(n17327), .A2(n19102), .B1(n17339), .B2(n23733), .ZN(
        n5124) );
  INV_X1 U24598 ( .A(n5128), .ZN(n27773) );
  AOI22_X1 U24599 ( .A1(n17329), .A2(n26622), .B1(n17341), .B2(n26591), .ZN(
        n5128) );
  AOI22_X1 U24600 ( .A1(n27011), .A2(matrix_mul_2D_5__2__12_), .B1(n26003), 
        .B2(matrix_mul_2D_5__3__12_), .ZN(n53390) );
  AOI22_X1 U24601 ( .A1(n27012), .A2(matrix_mul_2D_5__2__13_), .B1(n26057), 
        .B2(matrix_mul_2D_5__3__13_), .ZN(n5335) );
  AOI22_X1 U24602 ( .A1(n27013), .A2(matrix_mul_2D_5__2__14_), .B1(n25906), 
        .B2(matrix_mul_2D_5__3__14_), .ZN(n5331) );
  AOI221_X1 U24603 ( .B1(n19234), .B2(matrix_mul_2D_6__0__12_), .C1(n27040), 
        .C2(matrix_mul_2D_6__1__12_), .A(n5243), .ZN(n5242) );
  OAI22_X1 U24604 ( .A1(n2672), .A2(n25520), .B1(n2657), .B2(n23680), .ZN(
        n5243) );
  AOI221_X1 U24605 ( .B1(n21366), .B2(matrix_mul_2D_6__0__13_), .C1(n27041), 
        .C2(matrix_mul_2D_6__1__13_), .A(n5239), .ZN(n5238) );
  OAI22_X1 U24606 ( .A1(n2671), .A2(n19091), .B1(n265600), .B2(n265501), .ZN(
        n5239) );
  AOI221_X1 U24607 ( .B1(n21355), .B2(matrix_mul_2D_6__0__14_), .C1(n27042), 
        .C2(matrix_mul_2D_6__1__14_), .A(n52310), .ZN(n52300) );
  OAI22_X1 U24608 ( .A1(n2670), .A2(n26685), .B1(n265500), .B2(n22509), .ZN(
        n52310) );
  AOI22_X1 U24609 ( .A1(n22960), .A2(matrix_mul_2D_2__0__12_), .B1(n27082), 
        .B2(matrix_mul_2D_2__1__12_), .ZN(n4924) );
  AOI22_X1 U24610 ( .A1(n22961), .A2(matrix_mul_2D_2__0__13_), .B1(n27083), 
        .B2(matrix_mul_2D_2__1__13_), .ZN(n49200) );
  AOI22_X1 U24611 ( .A1(n22960), .A2(matrix_mul_2D_2__0__14_), .B1(n27084), 
        .B2(matrix_mul_2D_2__1__14_), .ZN(n49160) );
  INV_X1 U24612 ( .A(n5403), .ZN(n27756) );
  AOI22_X1 U24613 ( .A1(n17585), .A2(n25065), .B1(n17597), .B2(n21499), .ZN(
        n5403) );
  INV_X1 U24614 ( .A(n5215), .ZN(n27751) );
  AOI22_X1 U24615 ( .A1(n17419), .A2(n23725), .B1(n17431), .B2(n21489), .ZN(
        n5215) );
  INV_X1 U24616 ( .A(n5211), .ZN(n277501) );
  AOI22_X1 U24617 ( .A1(n17417), .A2(n20693), .B1(n17429), .B2(n21831), .ZN(
        n5211) );
  INV_X1 U24618 ( .A(n4898), .ZN(n27745) );
  AOI22_X1 U24619 ( .A1(n17755), .A2(n26591), .B1(n17767), .B2(n21462), .ZN(
        n4898) );
  INV_X1 U24620 ( .A(n4894), .ZN(n27744) );
  AOI22_X1 U24621 ( .A1(n17753), .A2(n23728), .B1(n17765), .B2(n23683), .ZN(
        n4894) );
  INV_X1 U24622 ( .A(n4712), .ZN(n27742) );
  AOI22_X1 U24623 ( .A1(n17593), .A2(n22533), .B1(n17605), .B2(n21833), .ZN(
        n4712) );
  INV_X1 U24624 ( .A(n5407), .ZN(n27757) );
  AOI22_X1 U24625 ( .A1(n17587), .A2(n20692), .B1(n17599), .B2(n17078), .ZN(
        n5407) );
  INV_X1 U24626 ( .A(n5411), .ZN(n27758) );
  AOI22_X1 U24627 ( .A1(n17589), .A2(n22536), .B1(n17601), .B2(n26055), .ZN(
        n5411) );
  INV_X1 U24628 ( .A(n5415), .ZN(n27759) );
  AOI22_X1 U24629 ( .A1(n17591), .A2(n22534), .B1(n17603), .B2(n26001), .ZN(
        n5415) );
  INV_X1 U24630 ( .A(n5207), .ZN(n27749) );
  AOI22_X1 U24631 ( .A1(n17415), .A2(n23732), .B1(n17427), .B2(n26073), .ZN(
        n5207) );
  INV_X1 U24632 ( .A(n52190), .ZN(n27752) );
  AOI22_X1 U24633 ( .A1(n17421), .A2(n24858), .B1(n17433), .B2(n260001), .ZN(
        n52190) );
  INV_X1 U24634 ( .A(n52230), .ZN(n27753) );
  AOI22_X1 U24635 ( .A1(n17423), .A2(n26589), .B1(n17435), .B2(n21433), .ZN(
        n52230) );
  INV_X1 U24636 ( .A(n52270), .ZN(n27754) );
  AOI22_X1 U24637 ( .A1(n17425), .A2(n20687), .B1(n17437), .B2(n26003), .ZN(
        n52270) );
  INV_X1 U24638 ( .A(n49060), .ZN(n27746) );
  AOI22_X1 U24639 ( .A1(n17757), .A2(n24859), .B1(n17769), .B2(n18496), .ZN(
        n49060) );
  INV_X1 U24640 ( .A(n49100), .ZN(n27747) );
  AOI22_X1 U24641 ( .A1(n17759), .A2(n23726), .B1(n17771), .B2(n25906), .ZN(
        n49100) );
  INV_X1 U24642 ( .A(n49140), .ZN(n27748) );
  AOI22_X1 U24643 ( .A1(n17761), .A2(n26904), .B1(n17773), .B2(n26947), .ZN(
        n49140) );
  XNOR2_X1 U24644 ( .A(n463), .B(n26974), .ZN(n26972) );
  NAND2_X1 U24645 ( .A1(n26969), .A2(n546), .ZN(n26974) );
  NOR2_X1 U24646 ( .A1(n27793), .A2(n549), .ZN(n54240) );
  INV_X1 U24647 ( .A(n54250), .ZN(n27793) );
  INV_X1 U24648 ( .A(n4370), .ZN(n27678) );
  AOI221_X1 U24649 ( .B1(n19843), .B2(n22498), .C1(N7413), .C2(n26202), .A(
        n25494), .ZN(n4370) );
  INV_X1 U24650 ( .A(n4372), .ZN(n27679) );
  AOI221_X1 U24651 ( .B1(n19845), .B2(n26548), .C1(N7412), .C2(n24354), .A(
        n25495), .ZN(n4372) );
  INV_X1 U24652 ( .A(n4373), .ZN(n276801) );
  AOI221_X1 U24653 ( .B1(n19847), .B2(n24857), .C1(N7411), .C2(n24357), .A(
        n19167), .ZN(n4373) );
  INV_X1 U24654 ( .A(n4374), .ZN(n27681) );
  AOI221_X1 U24655 ( .B1(n19849), .B2(n20690), .C1(N7410), .C2(n24342), .A(
        n25494), .ZN(n4374) );
  INV_X1 U24656 ( .A(n43750), .ZN(n27682) );
  AOI221_X1 U24657 ( .B1(n19851), .B2(n22496), .C1(N7409), .C2(n23340), .A(
        n25495), .ZN(n43750) );
  INV_X1 U24658 ( .A(n43760), .ZN(n27683) );
  AOI221_X1 U24659 ( .B1(n19853), .B2(n26547), .C1(N7408), .C2(n23337), .A(
        n19167), .ZN(n43760) );
  INV_X1 U24660 ( .A(n42130), .ZN(n27636) );
  AOI221_X1 U24661 ( .B1(n19927), .B2(n24406), .C1(N6802), .C2(n24361), .A(
        n25476), .ZN(n42130) );
  INV_X1 U24662 ( .A(n42150), .ZN(n27637) );
  AOI221_X1 U24663 ( .B1(n19929), .B2(n24405), .C1(N6801), .C2(n23343), .A(
        n19158), .ZN(n42150) );
  INV_X1 U24664 ( .A(n42160), .ZN(n27638) );
  AOI221_X1 U24665 ( .B1(n19931), .B2(n26545), .C1(N6800), .C2(n22306), .A(
        n25477), .ZN(n42160) );
  INV_X1 U24666 ( .A(n42170), .ZN(n27639) );
  AOI221_X1 U24667 ( .B1(n19933), .B2(n26546), .C1(N6799), .C2(n22296), .A(
        n25476), .ZN(n42170) );
  INV_X1 U24668 ( .A(n42180), .ZN(n27640) );
  AOI221_X1 U24669 ( .B1(n19935), .B2(n20689), .C1(N6798), .C2(n22286), .A(
        n19158), .ZN(n42180) );
  INV_X1 U24670 ( .A(n42190), .ZN(n27641) );
  AOI221_X1 U24671 ( .B1(n19937), .B2(n24857), .C1(N6797), .C2(n22316), .A(
        n25477), .ZN(n42190) );
  INV_X1 U24672 ( .A(n40520), .ZN(n27594) );
  AOI221_X1 U24673 ( .B1(n20011), .B2(n26544), .C1(N6202), .C2(n22311), .A(
        n25466), .ZN(n40520) );
  INV_X1 U24674 ( .A(n40540), .ZN(n27595) );
  AOI221_X1 U24675 ( .B1(n20013), .B2(n22500), .C1(N6201), .C2(n22301), .A(
        n19153), .ZN(n40540) );
  INV_X1 U24676 ( .A(n40550), .ZN(n27596) );
  AOI221_X1 U24677 ( .B1(n20015), .B2(n24405), .C1(N6200), .C2(n22291), .A(
        n25467), .ZN(n40550) );
  INV_X1 U24678 ( .A(n40560), .ZN(n27597) );
  AOI221_X1 U24679 ( .B1(n20017), .B2(n24406), .C1(N6199), .C2(n22321), .A(
        n25466), .ZN(n40560) );
  INV_X1 U24680 ( .A(n40570), .ZN(n27598) );
  AOI221_X1 U24681 ( .B1(n20019), .B2(n22499), .C1(N6198), .C2(n26848), .A(
        n19153), .ZN(n40570) );
  INV_X1 U24682 ( .A(n40580), .ZN(n27599) );
  AOI221_X1 U24683 ( .B1(n20021), .B2(n26793), .C1(N6197), .C2(n26851), .A(
        n25467), .ZN(n40580) );
  INV_X1 U24684 ( .A(n38910), .ZN(n27552) );
  AOI221_X1 U24685 ( .B1(n20095), .B2(n23669), .C1(N5606), .C2(n26854), .A(
        n25447), .ZN(n38910) );
  INV_X1 U24686 ( .A(n3893), .ZN(n27553) );
  AOI221_X1 U24687 ( .B1(n20097), .B2(n23670), .C1(N5605), .C2(n26844), .A(
        n19144), .ZN(n3893) );
  INV_X1 U24688 ( .A(n3894), .ZN(n27554) );
  AOI221_X1 U24689 ( .B1(n20099), .B2(n22495), .C1(N5604), .C2(n24346), .A(
        n25448), .ZN(n3894) );
  INV_X1 U24690 ( .A(n3895), .ZN(n27555) );
  AOI221_X1 U24691 ( .B1(n20101), .B2(n26782), .C1(N5603), .C2(n24352), .A(
        n25447), .ZN(n3895) );
  INV_X1 U24692 ( .A(n3896), .ZN(n27556) );
  AOI221_X1 U24693 ( .B1(n20103), .B2(n23667), .C1(N5602), .C2(n23334), .A(
        n19144), .ZN(n3896) );
  INV_X1 U24694 ( .A(n3897), .ZN(n27557) );
  AOI221_X1 U24695 ( .B1(n20105), .B2(n23668), .C1(N5601), .C2(n24340), .A(
        n25448), .ZN(n3897) );
  INV_X1 U24696 ( .A(n3731), .ZN(n27510) );
  AOI221_X1 U24697 ( .B1(n20179), .B2(n26545), .C1(N5014), .C2(n22303), .A(
        n25437), .ZN(n3731) );
  INV_X1 U24698 ( .A(n3733), .ZN(n27511) );
  AOI221_X1 U24699 ( .B1(n20181), .B2(n26786), .C1(N5013), .C2(n22293), .A(
        n19139), .ZN(n3733) );
  INV_X1 U24700 ( .A(n3734), .ZN(n27512) );
  AOI221_X1 U24701 ( .B1(n20183), .B2(n23670), .C1(N5012), .C2(n22283), .A(
        n25438), .ZN(n3734) );
  INV_X1 U24702 ( .A(n3735), .ZN(n27513) );
  AOI221_X1 U24703 ( .B1(n20185), .B2(n23669), .C1(N5011), .C2(n22313), .A(
        n25437), .ZN(n3735) );
  INV_X1 U24704 ( .A(n3736), .ZN(n27514) );
  AOI221_X1 U24705 ( .B1(n20187), .B2(n26544), .C1(N5010), .C2(n22308), .A(
        n19139), .ZN(n3736) );
  INV_X1 U24706 ( .A(n3737), .ZN(n27515) );
  AOI221_X1 U24707 ( .B1(n20189), .B2(n22501), .C1(N5009), .C2(n22298), .A(
        n25438), .ZN(n3737) );
  INV_X1 U24708 ( .A(n3572), .ZN(n27468) );
  AOI221_X1 U24709 ( .B1(n20263), .B2(n23668), .C1(N4395), .C2(n22288), .A(
        n25419), .ZN(n3572) );
  INV_X1 U24710 ( .A(n3574), .ZN(n27469) );
  AOI221_X1 U24711 ( .B1(n20265), .B2(n23667), .C1(N4394), .C2(n22318), .A(
        n19130), .ZN(n3574) );
  INV_X1 U24712 ( .A(n3575), .ZN(n274701) );
  AOI221_X1 U24713 ( .B1(n20267), .B2(n22498), .C1(N4393), .C2(n26847), .A(
        n25420), .ZN(n3575) );
  INV_X1 U24714 ( .A(n3576), .ZN(n27471) );
  AOI221_X1 U24715 ( .B1(n20269), .B2(n26548), .C1(N4392), .C2(n268501), .A(
        n25419), .ZN(n3576) );
  INV_X1 U24716 ( .A(n3577), .ZN(n27472) );
  AOI221_X1 U24717 ( .B1(n20271), .B2(n24403), .C1(N4391), .C2(n26852), .A(
        n19130), .ZN(n3577) );
  INV_X1 U24718 ( .A(n3578), .ZN(n27473) );
  AOI221_X1 U24719 ( .B1(n20273), .B2(n24404), .C1(N4390), .C2(n26843), .A(
        n25420), .ZN(n3578) );
  INV_X1 U24720 ( .A(n3412), .ZN(n27426) );
  AOI221_X1 U24721 ( .B1(n20347), .B2(n22495), .C1(N3809), .C2(n24348), .A(
        n25409), .ZN(n3412) );
  INV_X1 U24722 ( .A(n3414), .ZN(n27427) );
  AOI221_X1 U24723 ( .B1(n20349), .B2(n26547), .C1(N3808), .C2(n26198), .A(
        n19125), .ZN(n3414) );
  INV_X1 U24724 ( .A(n3415), .ZN(n27428) );
  AOI221_X1 U24725 ( .B1(n20351), .B2(n26541), .C1(N3807), .C2(n26194), .A(
        n25410), .ZN(n3415) );
  INV_X1 U24726 ( .A(n3416), .ZN(n27429) );
  AOI221_X1 U24727 ( .B1(n20353), .B2(n26541), .C1(N3806), .C2(n26206), .A(
        n25409), .ZN(n3416) );
  INV_X1 U24728 ( .A(n3417), .ZN(n274301) );
  AOI221_X1 U24729 ( .B1(n20355), .B2(n26543), .C1(N3805), .C2(n26469), .A(
        n19125), .ZN(n3417) );
  INV_X1 U24730 ( .A(n3418), .ZN(n27431) );
  AOI221_X1 U24731 ( .B1(n20357), .B2(n26546), .C1(N3804), .C2(n26463), .A(
        n25410), .ZN(n3418) );
  INV_X1 U24732 ( .A(n32520), .ZN(n27384) );
  AOI221_X1 U24733 ( .B1(n20383), .B2(n24404), .C1(N3216), .C2(n26457), .A(
        n25391), .ZN(n32520) );
  INV_X1 U24734 ( .A(n32550), .ZN(n27385) );
  AOI221_X1 U24735 ( .B1(n20385), .B2(n24403), .C1(N3215), .C2(n26475), .A(
        n19116), .ZN(n32550) );
  INV_X1 U24736 ( .A(n32560), .ZN(n27386) );
  AOI221_X1 U24737 ( .B1(n20387), .B2(n26542), .C1(N3214), .C2(n26471), .A(
        n25392), .ZN(n32560) );
  INV_X1 U24738 ( .A(n32570), .ZN(n27387) );
  AOI221_X1 U24739 ( .B1(n20389), .B2(n22500), .C1(N3213), .C2(n26466), .A(
        n25391), .ZN(n32570) );
  INV_X1 U24740 ( .A(n32580), .ZN(n27388) );
  AOI221_X1 U24741 ( .B1(n20391), .B2(n265401), .C1(N3212), .C2(n264601), .A(
        n19116), .ZN(n32580) );
  INV_X1 U24742 ( .A(n32590), .ZN(n27389) );
  AOI221_X1 U24743 ( .B1(n20393), .B2(n265401), .C1(N3211), .C2(n26478), .A(
        n25392), .ZN(n32590) );
  INV_X1 U24744 ( .A(n43950), .ZN(n27684) );
  AOI221_X1 U24745 ( .B1(n19831), .B2(n21314), .C1(N7492), .C2(n24265), .A(
        n25492), .ZN(n43950) );
  INV_X1 U24746 ( .A(n4397), .ZN(n27685) );
  AOI221_X1 U24747 ( .B1(n19833), .B2(n21296), .C1(N7491), .C2(n26044), .A(
        n19166), .ZN(n4397) );
  INV_X1 U24748 ( .A(n4398), .ZN(n27686) );
  AOI221_X1 U24749 ( .B1(n19835), .B2(n25619), .C1(N7490), .C2(n26007), .A(
        n25493), .ZN(n4398) );
  INV_X1 U24750 ( .A(n4399), .ZN(n27687) );
  AOI221_X1 U24751 ( .B1(n19837), .B2(n25625), .C1(N7489), .C2(n24238), .A(
        n25492), .ZN(n4399) );
  INV_X1 U24752 ( .A(n4400), .ZN(n27688) );
  AOI221_X1 U24753 ( .B1(n19839), .B2(n24198), .C1(N7488), .C2(n19255), .A(
        n19166), .ZN(n4400) );
  INV_X1 U24754 ( .A(n4401), .ZN(n27689) );
  AOI221_X1 U24755 ( .B1(n19841), .B2(n24210), .C1(N7487), .C2(n19252), .A(
        n25493), .ZN(n4401) );
  INV_X1 U24756 ( .A(n4235), .ZN(n27642) );
  AOI221_X1 U24757 ( .B1(n19915), .B2(n25274), .C1(N6894), .C2(n26307), .A(
        n25482), .ZN(n4235) );
  INV_X1 U24758 ( .A(n4237), .ZN(n27643) );
  AOI221_X1 U24759 ( .B1(n19917), .B2(n25261), .C1(N6893), .C2(n26313), .A(
        n25483), .ZN(n4237) );
  INV_X1 U24760 ( .A(n4238), .ZN(n27644) );
  AOI221_X1 U24761 ( .B1(n19919), .B2(n256201), .C1(N6892), .C2(n26036), .A(
        n19161), .ZN(n4238) );
  INV_X1 U24762 ( .A(n4239), .ZN(n27645) );
  AOI221_X1 U24763 ( .B1(n19921), .B2(n25626), .C1(N6891), .C2(n26311), .A(
        n25482), .ZN(n4239) );
  INV_X1 U24764 ( .A(n4240), .ZN(n27646) );
  AOI221_X1 U24765 ( .B1(n19923), .B2(n21294), .C1(N6890), .C2(n26018), .A(
        n25483), .ZN(n4240) );
  INV_X1 U24766 ( .A(n4241), .ZN(n27647) );
  AOI221_X1 U24767 ( .B1(n19925), .B2(n267401), .C1(N6889), .C2(n25995), .A(
        n19161), .ZN(n4241) );
  INV_X1 U24768 ( .A(n41870), .ZN(n27630) );
  AOI221_X1 U24769 ( .B1(n19939), .B2(n21320), .C1(N6720), .C2(n23159), .A(
        n25478), .ZN(n41870) );
  INV_X1 U24770 ( .A(n41890), .ZN(n27631) );
  AOI221_X1 U24771 ( .B1(n19941), .B2(n21308), .C1(N6719), .C2(n26062), .A(
        n19159), .ZN(n41890) );
  INV_X1 U24772 ( .A(n4190), .ZN(n27632) );
  AOI221_X1 U24773 ( .B1(n19943), .B2(n25623), .C1(N6718), .C2(n19254), .A(
        n25479), .ZN(n4190) );
  INV_X1 U24774 ( .A(n4191), .ZN(n27633) );
  AOI221_X1 U24775 ( .B1(n19945), .B2(n25627), .C1(N6717), .C2(n23204), .A(
        n25478), .ZN(n4191) );
  INV_X1 U24776 ( .A(n4192), .ZN(n27634) );
  AOI221_X1 U24777 ( .B1(n19947), .B2(n24195), .C1(N6716), .C2(n19256), .A(
        n19159), .ZN(n4192) );
  INV_X1 U24778 ( .A(n4193), .ZN(n27635) );
  AOI221_X1 U24779 ( .B1(n19949), .B2(n24204), .C1(N6715), .C2(n19253), .A(
        n25479), .ZN(n4193) );
  INV_X1 U24780 ( .A(n4074), .ZN(n27600) );
  AOI221_X1 U24781 ( .B1(n19999), .B2(n21312), .C1(N6281), .C2(n26773), .A(
        n25463), .ZN(n4074) );
  INV_X1 U24782 ( .A(n4076), .ZN(n27601) );
  AOI221_X1 U24783 ( .B1(n20001), .B2(n26731), .C1(N6280), .C2(n23147), .A(
        n25464), .ZN(n4076) );
  INV_X1 U24784 ( .A(n4077), .ZN(n27602) );
  AOI221_X1 U24785 ( .B1(n20003), .B2(n24199), .C1(N6279), .C2(n260401), .A(
        n19152), .ZN(n4077) );
  INV_X1 U24786 ( .A(n4078), .ZN(n27603) );
  AOI221_X1 U24787 ( .B1(n20005), .B2(n24211), .C1(N6278), .C2(n26004), .A(
        n25463), .ZN(n4078) );
  INV_X1 U24788 ( .A(n4079), .ZN(n27604) );
  AOI221_X1 U24789 ( .B1(n20007), .B2(n19222), .C1(N6277), .C2(n26778), .A(
        n25464), .ZN(n4079) );
  INV_X1 U24790 ( .A(n4080), .ZN(n27605) );
  AOI221_X1 U24791 ( .B1(n20009), .B2(n19216), .C1(N6276), .C2(n26772), .A(
        n19152), .ZN(n4080) );
  INV_X1 U24792 ( .A(n4030), .ZN(n27588) );
  AOI221_X1 U24793 ( .B1(n20023), .B2(n25278), .C1(N6113), .C2(n26309), .A(
        n25459), .ZN(n4030) );
  INV_X1 U24794 ( .A(n4032), .ZN(n27589) );
  AOI221_X1 U24795 ( .B1(n20025), .B2(n25270), .C1(N6112), .C2(n26317), .A(
        n25460), .ZN(n4032) );
  INV_X1 U24796 ( .A(n4033), .ZN(n27590) );
  AOI221_X1 U24797 ( .B1(n20027), .B2(n25624), .C1(N6111), .C2(n19257), .A(
        n19150), .ZN(n4033) );
  INV_X1 U24798 ( .A(n4034), .ZN(n27591) );
  AOI221_X1 U24799 ( .B1(n20029), .B2(n25628), .C1(N6110), .C2(n26315), .A(
        n25459), .ZN(n4034) );
  INV_X1 U24800 ( .A(n4035), .ZN(n27592) );
  AOI221_X1 U24801 ( .B1(n20031), .B2(n21306), .C1(N6109), .C2(n26031), .A(
        n25460), .ZN(n4035) );
  INV_X1 U24802 ( .A(n4036), .ZN(n27593) );
  AOI221_X1 U24803 ( .B1(n20033), .B2(n26733), .C1(N6108), .C2(n26009), .A(
        n19150), .ZN(n4036) );
  INV_X1 U24804 ( .A(n3913), .ZN(n27558) );
  AOI221_X1 U24805 ( .B1(n20083), .B2(n19221), .C1(N5695), .C2(n21849), .A(
        n25453), .ZN(n3913) );
  INV_X1 U24806 ( .A(n3915), .ZN(n27559) );
  AOI221_X1 U24807 ( .B1(n20085), .B2(n19215), .C1(N5694), .C2(n22875), .A(
        n25454), .ZN(n3915) );
  INV_X1 U24808 ( .A(n3916), .ZN(n27560) );
  AOI221_X1 U24809 ( .B1(n20087), .B2(n25276), .C1(N5693), .C2(n21837), .A(
        n19147), .ZN(n3916) );
  INV_X1 U24810 ( .A(n3917), .ZN(n27561) );
  AOI221_X1 U24811 ( .B1(n20089), .B2(n25263), .C1(N5692), .C2(n26043), .A(
        n25453), .ZN(n3917) );
  INV_X1 U24812 ( .A(n3918), .ZN(n27562) );
  AOI221_X1 U24813 ( .B1(n20091), .B2(n26739), .C1(N5691), .C2(n19310), .A(
        n25454), .ZN(n3918) );
  INV_X1 U24814 ( .A(n3919), .ZN(n27563) );
  AOI221_X1 U24815 ( .B1(n20093), .B2(n19305), .C1(N5690), .C2(n19308), .A(
        n19147), .ZN(n3919) );
  INV_X1 U24816 ( .A(n3869), .ZN(n27546) );
  AOI221_X1 U24817 ( .B1(n20107), .B2(n21318), .C1(N5527), .C2(n26769), .A(
        n25449), .ZN(n3869) );
  INV_X1 U24818 ( .A(n38710), .ZN(n27547) );
  AOI221_X1 U24819 ( .B1(n20109), .B2(n26730), .C1(N5526), .C2(n24253), .A(
        n25450), .ZN(n38710) );
  INV_X1 U24820 ( .A(n38720), .ZN(n27548) );
  AOI221_X1 U24821 ( .B1(n20111), .B2(n24196), .C1(N5525), .C2(n26069), .A(
        n19145), .ZN(n38720) );
  INV_X1 U24822 ( .A(n38730), .ZN(n27549) );
  AOI221_X1 U24823 ( .B1(n20113), .B2(n24205), .C1(N5524), .C2(n26014), .A(
        n25449), .ZN(n38730) );
  INV_X1 U24824 ( .A(n38740), .ZN(n27550) );
  AOI221_X1 U24825 ( .B1(n20115), .B2(n19224), .C1(N5523), .C2(n26775), .A(
        n25450), .ZN(n38740) );
  INV_X1 U24826 ( .A(n38750), .ZN(n27551) );
  AOI221_X1 U24827 ( .B1(n20117), .B2(n19220), .C1(N5522), .C2(n22847), .A(
        n19145), .ZN(n38750) );
  INV_X1 U24828 ( .A(n3753), .ZN(n27516) );
  AOI221_X1 U24829 ( .B1(n20167), .B2(n21315), .C1(N5096), .C2(n21845), .A(
        n25435), .ZN(n3753) );
  INV_X1 U24830 ( .A(n3755), .ZN(n27517) );
  AOI221_X1 U24831 ( .B1(n20169), .B2(n21297), .C1(N5095), .C2(n21473), .A(
        n19138), .ZN(n3755) );
  INV_X1 U24832 ( .A(n37560), .ZN(n27518) );
  AOI221_X1 U24833 ( .B1(n20171), .B2(n25619), .C1(N5094), .C2(n21460), .A(
        n25436), .ZN(n37560) );
  INV_X1 U24834 ( .A(n37570), .ZN(n27519) );
  AOI221_X1 U24835 ( .B1(n20173), .B2(n25625), .C1(N5093), .C2(n23169), .A(
        n25435), .ZN(n37570) );
  INV_X1 U24836 ( .A(n37580), .ZN(n27520) );
  AOI221_X1 U24837 ( .B1(n20175), .B2(n25261), .C1(N5092), .C2(n26766), .A(
        n19138), .ZN(n37580) );
  INV_X1 U24838 ( .A(n37590), .ZN(n27521) );
  AOI221_X1 U24839 ( .B1(n20177), .B2(n25264), .C1(N5091), .C2(n21467), .A(
        n25436), .ZN(n37590) );
  INV_X1 U24840 ( .A(n37090), .ZN(n27504) );
  AOI221_X1 U24841 ( .B1(n20191), .B2(n19223), .C1(N4922), .C2(n21857), .A(
        n25431), .ZN(n37090) );
  INV_X1 U24842 ( .A(n37110), .ZN(n27505) );
  AOI221_X1 U24843 ( .B1(n20193), .B2(n19219), .C1(N4921), .C2(n26776), .A(
        n25432), .ZN(n37110) );
  INV_X1 U24844 ( .A(n37120), .ZN(n27506) );
  AOI221_X1 U24845 ( .B1(n20195), .B2(n25280), .C1(N4920), .C2(n21841), .A(
        n19136), .ZN(n37120) );
  INV_X1 U24846 ( .A(n37130), .ZN(n27507) );
  AOI221_X1 U24847 ( .B1(n20197), .B2(n25272), .C1(N4919), .C2(n26061), .A(
        n25431), .ZN(n37130) );
  INV_X1 U24848 ( .A(n37140), .ZN(n27508) );
  AOI221_X1 U24849 ( .B1(n20199), .B2(n26732), .C1(N4918), .C2(n22859), .A(
        n25432), .ZN(n37140) );
  INV_X1 U24850 ( .A(n37150), .ZN(n27509) );
  AOI221_X1 U24851 ( .B1(n20201), .B2(n19304), .C1(N4917), .C2(n24232), .A(
        n19136), .ZN(n37150) );
  INV_X1 U24852 ( .A(n35940), .ZN(n27474) );
  AOI221_X1 U24853 ( .B1(n20251), .B2(n25276), .C1(N4484), .C2(n23154), .A(
        n25425), .ZN(n35940) );
  INV_X1 U24854 ( .A(n35960), .ZN(n27475) );
  AOI221_X1 U24855 ( .B1(n20253), .B2(n25277), .C1(N4483), .C2(n21481), .A(
        n25426), .ZN(n35960) );
  INV_X1 U24856 ( .A(n35970), .ZN(n27476) );
  AOI221_X1 U24857 ( .B1(n20255), .B2(n256201), .C1(N4482), .C2(n22854), .A(
        n19133), .ZN(n35970) );
  INV_X1 U24858 ( .A(n35980), .ZN(n27477) );
  AOI221_X1 U24859 ( .B1(n20257), .B2(n25626), .C1(N4481), .C2(n26781), .A(
        n25425), .ZN(n35980) );
  INV_X1 U24860 ( .A(n35990), .ZN(n27478) );
  AOI221_X1 U24861 ( .B1(n20259), .B2(n21293), .C1(N4480), .C2(n21483), .A(
        n25426), .ZN(n35990) );
  INV_X1 U24862 ( .A(n36000), .ZN(n27479) );
  AOI221_X1 U24863 ( .B1(n20261), .B2(n21311), .C1(N4479), .C2(n22869), .A(
        n19133), .ZN(n36000) );
  INV_X1 U24864 ( .A(n35500), .ZN(n27462) );
  AOI221_X1 U24865 ( .B1(n20275), .B2(n21321), .C1(N4316), .C2(n21853), .A(
        n25421), .ZN(n35500) );
  INV_X1 U24866 ( .A(n35520), .ZN(n27463) );
  AOI221_X1 U24867 ( .B1(n20277), .B2(n21309), .C1(N4315), .C2(n21479), .A(
        n19131), .ZN(n35520) );
  INV_X1 U24868 ( .A(n3553), .ZN(n27464) );
  AOI221_X1 U24869 ( .B1(n20279), .B2(n25623), .C1(N4314), .C2(n21469), .A(
        n25422), .ZN(n3553) );
  INV_X1 U24870 ( .A(n3554), .ZN(n27465) );
  AOI221_X1 U24871 ( .B1(n20281), .B2(n25627), .C1(N4313), .C2(n23182), .A(
        n25421), .ZN(n3554) );
  INV_X1 U24872 ( .A(n3555), .ZN(n27466) );
  AOI221_X1 U24873 ( .B1(n20283), .B2(n25270), .C1(N4312), .C2(n22835), .A(
        n19131), .ZN(n3555) );
  INV_X1 U24874 ( .A(n3556), .ZN(n27467) );
  AOI221_X1 U24875 ( .B1(n20285), .B2(n25273), .C1(N4311), .C2(n21471), .A(
        n25422), .ZN(n3556) );
  INV_X1 U24876 ( .A(n34340), .ZN(n27432) );
  AOI221_X1 U24877 ( .B1(n20335), .B2(n24199), .C1(N3891), .C2(n26038), .A(
        n25407), .ZN(n34340) );
  INV_X1 U24878 ( .A(n3437), .ZN(n27433) );
  AOI221_X1 U24879 ( .B1(n20337), .B2(n24211), .C1(N3890), .C2(n21843), .A(
        n19124), .ZN(n3437) );
  INV_X1 U24880 ( .A(n3438), .ZN(n27434) );
  AOI221_X1 U24881 ( .B1(n20339), .B2(n25277), .C1(N3889), .C2(n21847), .A(
        n25408), .ZN(n3438) );
  INV_X1 U24882 ( .A(n3439), .ZN(n27435) );
  AOI221_X1 U24883 ( .B1(n20341), .B2(n25260), .C1(N3888), .C2(n267801), .A(
        n25407), .ZN(n3439) );
  INV_X1 U24884 ( .A(n3440), .ZN(n27436) );
  AOI221_X1 U24885 ( .B1(n20343), .B2(n19222), .C1(N3887), .C2(n21835), .A(
        n19124), .ZN(n3440) );
  INV_X1 U24886 ( .A(n3441), .ZN(n27437) );
  AOI221_X1 U24887 ( .B1(n20345), .B2(n19216), .C1(N3886), .C2(n23185), .A(
        n25408), .ZN(n3441) );
  INV_X1 U24888 ( .A(n3390), .ZN(n274201) );
  AOI221_X1 U24889 ( .B1(matrix_mul_2D_1__5__20_), .B2(n25280), .C1(N3720), 
        .C2(n24250), .A(n25403), .ZN(n3390) );
  INV_X1 U24890 ( .A(n3392), .ZN(n27421) );
  AOI221_X1 U24891 ( .B1(matrix_mul_2D_1__5__19_), .B2(n25281), .C1(N3719), 
        .C2(n21497), .A(n25404), .ZN(n3392) );
  INV_X1 U24892 ( .A(n3393), .ZN(n27422) );
  AOI221_X1 U24893 ( .B1(matrix_mul_2D_1__5__18_), .B2(n25624), .C1(N3718), 
        .C2(n26768), .A(n19122), .ZN(n3393) );
  INV_X1 U24894 ( .A(n3394), .ZN(n27423) );
  AOI221_X1 U24895 ( .B1(matrix_mul_2D_1__5__17_), .B2(n25628), .C1(N3717), 
        .C2(n26777), .A(n25403), .ZN(n3394) );
  INV_X1 U24896 ( .A(n3395), .ZN(n27424) );
  AOI221_X1 U24897 ( .B1(matrix_mul_2D_1__5__16_), .B2(n21305), .C1(N3716), 
        .C2(n21493), .A(n25404), .ZN(n3395) );
  INV_X1 U24898 ( .A(n3396), .ZN(n27425) );
  AOI221_X1 U24899 ( .B1(matrix_mul_2D_1__5__15_), .B2(n21317), .C1(N3715), 
        .C2(n26774), .A(n19122), .ZN(n3396) );
  INV_X1 U24900 ( .A(n3227), .ZN(n27378) );
  AOI221_X1 U24901 ( .B1(n20395), .B2(n24196), .C1(N3134), .C2(n26761), .A(
        n25393), .ZN(n3227) );
  INV_X1 U24902 ( .A(n3230), .ZN(n27379) );
  AOI221_X1 U24903 ( .B1(n20397), .B2(n24205), .C1(N3133), .C2(n21851), .A(
        n19117), .ZN(n3230) );
  INV_X1 U24904 ( .A(n3231), .ZN(n273801) );
  AOI221_X1 U24905 ( .B1(n20399), .B2(n25281), .C1(N3132), .C2(n21855), .A(
        n25394), .ZN(n3231) );
  INV_X1 U24906 ( .A(n3232), .ZN(n27381) );
  AOI221_X1 U24907 ( .B1(n20401), .B2(n25269), .C1(N3131), .C2(n22864), .A(
        n25393), .ZN(n3232) );
  INV_X1 U24908 ( .A(n3233), .ZN(n27382) );
  AOI221_X1 U24909 ( .B1(n20403), .B2(n19224), .C1(N3130), .C2(n21839), .A(
        n19117), .ZN(n3233) );
  INV_X1 U24910 ( .A(n3234), .ZN(n27383) );
  AOI221_X1 U24911 ( .B1(n20405), .B2(n19220), .C1(N3129), .C2(n267601), .A(
        n25394), .ZN(n3234) );
  INV_X1 U24912 ( .A(n4420), .ZN(n276901) );
  AOI221_X1 U24913 ( .B1(n19819), .B2(n21475), .C1(N7581), .C2(n25854), .A(
        n25499), .ZN(n4420) );
  INV_X1 U24914 ( .A(n4422), .ZN(n27691) );
  AOI221_X1 U24915 ( .B1(n19821), .B2(n21477), .C1(N7580), .C2(n27178), .A(
        n19169), .ZN(n4422) );
  INV_X1 U24916 ( .A(n4423), .ZN(n27692) );
  AOI221_X1 U24917 ( .B1(n19823), .B2(n25145), .C1(N7579), .C2(n22897), .A(
        n25498), .ZN(n4423) );
  INV_X1 U24918 ( .A(n4424), .ZN(n27693) );
  AOI221_X1 U24919 ( .B1(n19825), .B2(n24243), .C1(N7578), .C2(n25850), .A(
        n25498), .ZN(n4424) );
  INV_X1 U24920 ( .A(n4425), .ZN(n27694) );
  AOI221_X1 U24921 ( .B1(n19827), .B2(n26027), .C1(N7577), .C2(n25855), .A(
        n25499), .ZN(n4425) );
  INV_X1 U24922 ( .A(n4426), .ZN(n27695) );
  AOI221_X1 U24923 ( .B1(n19829), .B2(n260301), .C1(N7576), .C2(n22899), .A(
        n19169), .ZN(n4426) );
  INV_X1 U24924 ( .A(n4257), .ZN(n27648) );
  AOI221_X1 U24925 ( .B1(n19903), .B2(n24244), .C1(N6976), .C2(n25817), .A(
        n25480), .ZN(n4257) );
  INV_X1 U24926 ( .A(n4259), .ZN(n27649) );
  AOI221_X1 U24927 ( .B1(n19905), .B2(n26023), .C1(N6975), .C2(n27183), .A(
        n19160), .ZN(n4259) );
  INV_X1 U24928 ( .A(n4260), .ZN(n27650) );
  AOI221_X1 U24929 ( .B1(n19907), .B2(n26026), .C1(N6974), .C2(n25809), .A(
        n25481), .ZN(n4260) );
  INV_X1 U24930 ( .A(n4261), .ZN(n27651) );
  AOI221_X1 U24931 ( .B1(n19909), .B2(n26029), .C1(N6973), .C2(n25813), .A(
        n25480), .ZN(n4261) );
  INV_X1 U24932 ( .A(n4262), .ZN(n27652) );
  AOI221_X1 U24933 ( .B1(n19911), .B2(n19309), .C1(N6972), .C2(n25796), .A(
        n19160), .ZN(n4262) );
  INV_X1 U24934 ( .A(n42630), .ZN(n27653) );
  AOI221_X1 U24935 ( .B1(n19913), .B2(n26024), .C1(N6971), .C2(n27179), .A(
        n25481), .ZN(n42630) );
  INV_X1 U24936 ( .A(n40960), .ZN(n27606) );
  AOI221_X1 U24937 ( .B1(n19987), .B2(n26025), .C1(N6370), .C2(n24528), .A(
        n25470), .ZN(n40960) );
  INV_X1 U24938 ( .A(n40980), .ZN(n27607) );
  AOI221_X1 U24939 ( .B1(n19989), .B2(n26028), .C1(N6369), .C2(n25552), .A(
        n19155), .ZN(n40980) );
  INV_X1 U24940 ( .A(n40990), .ZN(n27608) );
  AOI221_X1 U24941 ( .B1(n19991), .B2(n26022), .C1(N6368), .C2(n25801), .A(
        n25471), .ZN(n40990) );
  INV_X1 U24942 ( .A(n41000), .ZN(n27609) );
  AOI221_X1 U24943 ( .B1(n19993), .B2(n23172), .C1(N6367), .C2(n25805), .A(
        n25470), .ZN(n41000) );
  INV_X1 U24944 ( .A(n41010), .ZN(n27610) );
  AOI221_X1 U24945 ( .B1(n19995), .B2(n21475), .C1(N6366), .C2(n25822), .A(
        n19155), .ZN(n41010) );
  INV_X1 U24946 ( .A(n41020), .ZN(n27611) );
  AOI221_X1 U24947 ( .B1(n19997), .B2(n21478), .C1(N6365), .C2(n25826), .A(
        n25471), .ZN(n41020) );
  INV_X1 U24948 ( .A(n4004), .ZN(n27582) );
  AOI221_X1 U24949 ( .B1(n20035), .B2(n21485), .C1(N6034), .C2(n25840), .A(
        n25462), .ZN(n4004) );
  INV_X1 U24950 ( .A(n40060), .ZN(n27583) );
  AOI221_X1 U24951 ( .B1(n20037), .B2(n21487), .C1(N6033), .C2(n27233), .A(
        n19151), .ZN(n40060) );
  INV_X1 U24952 ( .A(n40070), .ZN(n27584) );
  AOI221_X1 U24953 ( .B1(n20039), .B2(n25127), .C1(N6032), .C2(n22901), .A(
        n25461), .ZN(n40070) );
  INV_X1 U24954 ( .A(n40080), .ZN(n27585) );
  AOI221_X1 U24955 ( .B1(n20041), .B2(n24234), .C1(N6031), .C2(n25836), .A(
        n25461), .ZN(n40080) );
  INV_X1 U24956 ( .A(n40090), .ZN(n27586) );
  AOI221_X1 U24957 ( .B1(n20043), .B2(n26051), .C1(N6030), .C2(n25841), .A(
        n25462), .ZN(n40090) );
  INV_X1 U24958 ( .A(n40100), .ZN(n27587) );
  AOI221_X1 U24959 ( .B1(n20045), .B2(n26054), .C1(N6029), .C2(n22903), .A(
        n19151), .ZN(n40100) );
  INV_X1 U24960 ( .A(n39350), .ZN(n27564) );
  AOI221_X1 U24961 ( .B1(n20071), .B2(n23171), .C1(N5774), .C2(n21420), .A(
        n25451), .ZN(n39350) );
  INV_X1 U24962 ( .A(n39370), .ZN(n27565) );
  AOI221_X1 U24963 ( .B1(n20073), .B2(n22850), .C1(N5773), .C2(n25851), .A(
        n25452), .ZN(n39370) );
  INV_X1 U24964 ( .A(n39380), .ZN(n27566) );
  AOI221_X1 U24965 ( .B1(n20075), .B2(n26027), .C1(N5772), .C2(n25844), .A(
        n19146), .ZN(n39380) );
  INV_X1 U24966 ( .A(n39390), .ZN(n27567) );
  AOI221_X1 U24967 ( .B1(n20077), .B2(n260301), .C1(N5771), .C2(n25852), .A(
        n25451), .ZN(n39390) );
  INV_X1 U24968 ( .A(n39400), .ZN(n27568) );
  AOI221_X1 U24969 ( .B1(n20079), .B2(n26023), .C1(N5770), .C2(n25856), .A(
        n25452), .ZN(n39400) );
  INV_X1 U24970 ( .A(n39410), .ZN(n27569) );
  AOI221_X1 U24971 ( .B1(n20081), .B2(n24244), .C1(N5769), .C2(n25848), .A(
        n19146), .ZN(n39410) );
  INV_X1 U24972 ( .A(n38470), .ZN(n27540) );
  AOI221_X1 U24973 ( .B1(n20119), .B2(n24235), .C1(N5438), .C2(n25783), .A(
        n25443), .ZN(n38470) );
  INV_X1 U24974 ( .A(n38490), .ZN(n27541) );
  AOI221_X1 U24975 ( .B1(n20121), .B2(n26047), .C1(N5437), .C2(n27238), .A(
        n19142), .ZN(n38490) );
  INV_X1 U24976 ( .A(n38500), .ZN(n27542) );
  AOI221_X1 U24977 ( .B1(n20123), .B2(n260501), .C1(N5436), .C2(n25775), .A(
        n25444), .ZN(n38500) );
  INV_X1 U24978 ( .A(n38510), .ZN(n27543) );
  AOI221_X1 U24979 ( .B1(n20125), .B2(n26053), .C1(N5435), .C2(n25779), .A(
        n25443), .ZN(n38510) );
  INV_X1 U24980 ( .A(n38520), .ZN(n27544) );
  AOI221_X1 U24981 ( .B1(n20127), .B2(n19307), .C1(N5434), .C2(n25762), .A(
        n19142), .ZN(n38520) );
  INV_X1 U24982 ( .A(n38530), .ZN(n27545) );
  AOI221_X1 U24983 ( .B1(n20129), .B2(n26048), .C1(N5433), .C2(n27234), .A(
        n25444), .ZN(n38530) );
  INV_X1 U24984 ( .A(n3775), .ZN(n27522) );
  AOI221_X1 U24985 ( .B1(n20155), .B2(n26026), .C1(N5188), .C2(n25818), .A(
        n25441), .ZN(n3775) );
  INV_X1 U24986 ( .A(n3777), .ZN(n27523) );
  AOI221_X1 U24987 ( .B1(n20157), .B2(n26029), .C1(N5187), .C2(n25820), .A(
        n19141), .ZN(n3777) );
  INV_X1 U24988 ( .A(n3778), .ZN(n27524) );
  AOI221_X1 U24989 ( .B1(n20159), .B2(n19309), .C1(N5186), .C2(n25810), .A(
        n25442), .ZN(n3778) );
  INV_X1 U24990 ( .A(n3779), .ZN(n27525) );
  AOI221_X1 U24991 ( .B1(n20161), .B2(n23172), .C1(N5185), .C2(n25814), .A(
        n25441), .ZN(n3779) );
  INV_X1 U24992 ( .A(n3780), .ZN(n27526) );
  AOI221_X1 U24993 ( .B1(n20163), .B2(n26025), .C1(N5184), .C2(n25797), .A(
        n19141), .ZN(n3780) );
  INV_X1 U24994 ( .A(n3781), .ZN(n27527) );
  AOI221_X1 U24995 ( .B1(n20165), .B2(n26028), .C1(N5183), .C2(n25799), .A(
        n25442), .ZN(n3781) );
  INV_X1 U24996 ( .A(n3687), .ZN(n27498) );
  AOI221_X1 U24997 ( .B1(n20203), .B2(n26049), .C1(N4840), .C2(n24534), .A(
        n25433), .ZN(n3687) );
  INV_X1 U24998 ( .A(n3689), .ZN(n27499) );
  AOI221_X1 U24999 ( .B1(n20205), .B2(n26052), .C1(N4839), .C2(n25550), .A(
        n19137), .ZN(n3689) );
  INV_X1 U25000 ( .A(n3690), .ZN(n27500) );
  AOI221_X1 U25001 ( .B1(n20207), .B2(n26046), .C1(N4838), .C2(n25767), .A(
        n25434), .ZN(n3690) );
  INV_X1 U25002 ( .A(n3691), .ZN(n27501) );
  AOI221_X1 U25003 ( .B1(n20209), .B2(n23192), .C1(N4837), .C2(n25771), .A(
        n25433), .ZN(n3691) );
  INV_X1 U25004 ( .A(n3692), .ZN(n27502) );
  AOI221_X1 U25005 ( .B1(n20211), .B2(n21485), .C1(N4836), .C2(n25788), .A(
        n19137), .ZN(n3692) );
  INV_X1 U25006 ( .A(n3693), .ZN(n27503) );
  AOI221_X1 U25007 ( .B1(n20213), .B2(n21488), .C1(N4835), .C2(n25792), .A(
        n25434), .ZN(n3693) );
  INV_X1 U25008 ( .A(n3616), .ZN(n274801) );
  AOI221_X1 U25009 ( .B1(n20239), .B2(n26024), .C1(N4566), .C2(n25553), .A(
        n25423), .ZN(n3616) );
  INV_X1 U25010 ( .A(n3619), .ZN(n27481) );
  AOI221_X1 U25011 ( .B1(n20241), .B2(n267701), .C1(N4565), .C2(n24527), .A(
        n19132), .ZN(n3619) );
  INV_X1 U25012 ( .A(n3620), .ZN(n27482) );
  AOI221_X1 U25013 ( .B1(n20243), .B2(n21476), .C1(N4564), .C2(n25802), .A(
        n25424), .ZN(n3620) );
  INV_X1 U25014 ( .A(n36210), .ZN(n27483) );
  AOI221_X1 U25015 ( .B1(n20245), .B2(n21477), .C1(N4563), .C2(n25806), .A(
        n25423), .ZN(n36210) );
  INV_X1 U25016 ( .A(n36220), .ZN(n27484) );
  AOI221_X1 U25017 ( .B1(n20247), .B2(n267701), .C1(N4562), .C2(n25823), .A(
        n19132), .ZN(n36220) );
  INV_X1 U25018 ( .A(n36230), .ZN(n27485) );
  AOI221_X1 U25019 ( .B1(n20249), .B2(n22849), .C1(N4561), .C2(n25827), .A(
        n25424), .ZN(n36230) );
  INV_X1 U25020 ( .A(n3528), .ZN(n27456) );
  AOI221_X1 U25021 ( .B1(n20287), .B2(n23191), .C1(N4227), .C2(n21417), .A(
        n25415), .ZN(n3528) );
  INV_X1 U25022 ( .A(n3530), .ZN(n27457) );
  AOI221_X1 U25023 ( .B1(n20289), .B2(n22841), .C1(N4226), .C2(n25837), .A(
        n25416), .ZN(n3530) );
  INV_X1 U25024 ( .A(n3531), .ZN(n27458) );
  AOI221_X1 U25025 ( .B1(n20291), .B2(n26051), .C1(N4225), .C2(n25830), .A(
        n19128), .ZN(n3531) );
  INV_X1 U25026 ( .A(n35320), .ZN(n27459) );
  AOI221_X1 U25027 ( .B1(n20293), .B2(n26054), .C1(N4224), .C2(n25838), .A(
        n25415), .ZN(n35320) );
  INV_X1 U25028 ( .A(n35330), .ZN(n274601) );
  AOI221_X1 U25029 ( .B1(n20295), .B2(n26047), .C1(N4223), .C2(n25842), .A(
        n25416), .ZN(n35330) );
  INV_X1 U25030 ( .A(n35340), .ZN(n27461) );
  AOI221_X1 U25031 ( .B1(n20297), .B2(n24235), .C1(N4222), .C2(n25834), .A(
        n19128), .ZN(n35340) );
  INV_X1 U25032 ( .A(n33680), .ZN(n27414) );
  AOI221_X1 U25033 ( .B1(matrix_mul_2D_1__4__20_), .B2(n260501), .C1(N3641), 
        .C2(n25784), .A(n25405), .ZN(n33680) );
  INV_X1 U25034 ( .A(n33700), .ZN(n27415) );
  AOI221_X1 U25035 ( .B1(matrix_mul_2D_1__4__19_), .B2(n26053), .C1(N3640), 
        .C2(n25786), .A(n19123), .ZN(n33700) );
  INV_X1 U25036 ( .A(n33710), .ZN(n27416) );
  AOI221_X1 U25037 ( .B1(matrix_mul_2D_1__4__18_), .B2(n19307), .C1(N3639), 
        .C2(n25776), .A(n25406), .ZN(n33710) );
  INV_X1 U25038 ( .A(n33720), .ZN(n27417) );
  AOI221_X1 U25039 ( .B1(matrix_mul_2D_1__4__17_), .B2(n23192), .C1(N3638), 
        .C2(n25780), .A(n25405), .ZN(n33720) );
  INV_X1 U25040 ( .A(n33730), .ZN(n27418) );
  AOI221_X1 U25041 ( .B1(matrix_mul_2D_1__4__16_), .B2(n26049), .C1(N3637), 
        .C2(n25763), .A(n19123), .ZN(n33730) );
  INV_X1 U25042 ( .A(n33740), .ZN(n27419) );
  AOI221_X1 U25043 ( .B1(matrix_mul_2D_1__4__15_), .B2(n26052), .C1(N3636), 
        .C2(n25765), .A(n25406), .ZN(n33740) );
  INV_X1 U25044 ( .A(n32020), .ZN(n27372) );
  AOI221_X1 U25045 ( .B1(n20407), .B2(n26048), .C1(N3042), .C2(n24561), .A(
        n25387), .ZN(n32020) );
  INV_X1 U25046 ( .A(n32050), .ZN(n27373) );
  AOI221_X1 U25047 ( .B1(n20409), .B2(n26764), .C1(N3041), .C2(n24532), .A(
        n19114), .ZN(n32050) );
  INV_X1 U25048 ( .A(n32060), .ZN(n27374) );
  AOI221_X1 U25049 ( .B1(n20411), .B2(n21486), .C1(N3040), .C2(n25768), .A(
        n25388), .ZN(n32060) );
  INV_X1 U25050 ( .A(n32070), .ZN(n27375) );
  AOI221_X1 U25051 ( .B1(n20413), .B2(n21487), .C1(N3039), .C2(n25772), .A(
        n25387), .ZN(n32070) );
  INV_X1 U25052 ( .A(n32080), .ZN(n27376) );
  AOI221_X1 U25053 ( .B1(n20415), .B2(n26764), .C1(N3038), .C2(n25789), .A(
        n19114), .ZN(n32080) );
  INV_X1 U25054 ( .A(n32090), .ZN(n27377) );
  AOI221_X1 U25055 ( .B1(n20417), .B2(n22840), .C1(N3037), .C2(n25793), .A(
        n25388), .ZN(n32090) );
  INV_X1 U25056 ( .A(n4541), .ZN(n277201) );
  AOI221_X1 U25057 ( .B1(n19759), .B2(n25115), .C1(N7999), .C2(n24444), .A(
        n25504), .ZN(n4541) );
  INV_X1 U25058 ( .A(n4544), .ZN(n27721) );
  AOI221_X1 U25059 ( .B1(n19761), .B2(n19034), .C1(N7998), .C2(n24811), .A(
        n19172), .ZN(n4544) );
  INV_X1 U25060 ( .A(n4545), .ZN(n27722) );
  AOI221_X1 U25061 ( .B1(n19763), .B2(n25116), .C1(N7997), .C2(n24445), .A(
        n25505), .ZN(n4545) );
  INV_X1 U25062 ( .A(n45460), .ZN(n27723) );
  AOI221_X1 U25063 ( .B1(n19765), .B2(n25115), .C1(N7996), .C2(n24447), .A(
        n25504), .ZN(n45460) );
  INV_X1 U25064 ( .A(n45470), .ZN(n27724) );
  AOI221_X1 U25065 ( .B1(n19767), .B2(n19034), .C1(N7995), .C2(n24442), .A(
        n19172), .ZN(n45470) );
  INV_X1 U25066 ( .A(n45480), .ZN(n27725) );
  AOI221_X1 U25067 ( .B1(n19769), .B2(n25116), .C1(N7994), .C2(n24441), .A(
        n25505), .ZN(n45480) );
  INV_X1 U25068 ( .A(n45170), .ZN(n27714) );
  AOI221_X1 U25069 ( .B1(n19771), .B2(n26536), .C1(N7917), .C2(n19242), .A(
        n25506), .ZN(n45170) );
  INV_X1 U25070 ( .A(n45190), .ZN(n27715) );
  AOI221_X1 U25071 ( .B1(n19773), .B2(n22484), .C1(N7916), .C2(n21443), .A(
        n19173), .ZN(n45190) );
  INV_X1 U25072 ( .A(n45200), .ZN(n27716) );
  AOI221_X1 U25073 ( .B1(n19775), .B2(n22480), .C1(N7915), .C2(n20528), .A(
        n25507), .ZN(n45200) );
  INV_X1 U25074 ( .A(n45210), .ZN(n27717) );
  AOI221_X1 U25075 ( .B1(n19777), .B2(n22483), .C1(N7914), .C2(n24738), .A(
        n25506), .ZN(n45210) );
  INV_X1 U25076 ( .A(n45220), .ZN(n27718) );
  AOI221_X1 U25077 ( .B1(n19779), .B2(n26537), .C1(N7913), .C2(n21439), .A(
        n19173), .ZN(n45220) );
  INV_X1 U25078 ( .A(n45230), .ZN(n27719) );
  AOI221_X1 U25079 ( .B1(n19781), .B2(n19268), .C1(N7912), .C2(n25964), .A(
        n25507), .ZN(n45230) );
  INV_X1 U25080 ( .A(n4493), .ZN(n27708) );
  AOI221_X1 U25081 ( .B1(n19783), .B2(n24989), .C1(N7828), .C2(n25704), .A(
        n25500), .ZN(n4493) );
  INV_X1 U25082 ( .A(n4495), .ZN(n27709) );
  AOI221_X1 U25083 ( .B1(n19785), .B2(n17087), .C1(N7827), .C2(n25696), .A(
        n19170), .ZN(n4495) );
  INV_X1 U25084 ( .A(n4496), .ZN(n277101) );
  AOI221_X1 U25085 ( .B1(n19787), .B2(n22749), .C1(N7826), .C2(n25712), .A(
        n25501), .ZN(n4496) );
  INV_X1 U25086 ( .A(n4497), .ZN(n27711) );
  AOI221_X1 U25087 ( .B1(n19789), .B2(n22748), .C1(N7825), .C2(n25732), .A(
        n25500), .ZN(n4497) );
  INV_X1 U25088 ( .A(n4498), .ZN(n27712) );
  AOI221_X1 U25089 ( .B1(n19791), .B2(n20787), .C1(N7824), .C2(n25728), .A(
        n19170), .ZN(n4498) );
  INV_X1 U25090 ( .A(n4499), .ZN(n27713) );
  AOI221_X1 U25091 ( .B1(n19793), .B2(n20780), .C1(N7823), .C2(n25733), .A(
        n25501), .ZN(n4499) );
  INV_X1 U25092 ( .A(n44690), .ZN(n27702) );
  AOI221_X1 U25093 ( .B1(n19795), .B2(n19076), .C1(N7749), .C2(n25750), .A(
        n25502), .ZN(n44690) );
  INV_X1 U25094 ( .A(n44710), .ZN(n27703) );
  AOI221_X1 U25095 ( .B1(n19797), .B2(n19077), .C1(N7748), .C2(n20799), .A(
        n19171), .ZN(n44710) );
  INV_X1 U25096 ( .A(n44720), .ZN(n27704) );
  AOI221_X1 U25097 ( .B1(n19799), .B2(n25304), .C1(N7747), .C2(n19287), .A(
        n25503), .ZN(n44720) );
  INV_X1 U25098 ( .A(n44730), .ZN(n27705) );
  AOI221_X1 U25099 ( .B1(n19801), .B2(n24178), .C1(N7746), .C2(n20523), .A(
        n25502), .ZN(n44730) );
  INV_X1 U25100 ( .A(n44740), .ZN(n27706) );
  AOI221_X1 U25101 ( .B1(n19803), .B2(n25306), .C1(N7745), .C2(n20525), .A(
        n19171), .ZN(n44740) );
  INV_X1 U25102 ( .A(n44750), .ZN(n27707) );
  AOI221_X1 U25103 ( .B1(n19805), .B2(n25308), .C1(N7744), .C2(n20792), .A(
        n25503), .ZN(n44750) );
  INV_X1 U25104 ( .A(n44440), .ZN(n27696) );
  AOI221_X1 U25105 ( .B1(n19807), .B2(n25925), .C1(N7660), .C2(n21215), .A(
        n25496), .ZN(n44440) );
  INV_X1 U25106 ( .A(n44460), .ZN(n27697) );
  AOI221_X1 U25107 ( .B1(n19809), .B2(n25914), .C1(N7659), .C2(n25562), .A(
        n19168), .ZN(n44460) );
  INV_X1 U25108 ( .A(n4447), .ZN(n27698) );
  AOI221_X1 U25109 ( .B1(n19811), .B2(n25596), .C1(N7658), .C2(n24539), .A(
        n25497), .ZN(n4447) );
  INV_X1 U25110 ( .A(n4448), .ZN(n27699) );
  AOI221_X1 U25111 ( .B1(n19813), .B2(n256001), .C1(N7657), .C2(n21224), .A(
        n25496), .ZN(n4448) );
  INV_X1 U25112 ( .A(n4449), .ZN(n277001) );
  AOI221_X1 U25113 ( .B1(n19815), .B2(n25926), .C1(N7656), .C2(n25563), .A(
        n19168), .ZN(n4449) );
  INV_X1 U25114 ( .A(n4450), .ZN(n27701) );
  AOI221_X1 U25115 ( .B1(n19817), .B2(n25915), .C1(N7655), .C2(n19050), .A(
        n25497), .ZN(n4450) );
  INV_X1 U25116 ( .A(n43450), .ZN(n27672) );
  AOI221_X1 U25117 ( .B1(n19855), .B2(n22480), .C1(N7324), .C2(n25965), .A(
        n25488), .ZN(n43450) );
  INV_X1 U25118 ( .A(n43480), .ZN(n27673) );
  AOI221_X1 U25119 ( .B1(n19857), .B2(n22484), .C1(N7323), .C2(n17098), .A(
        n25489), .ZN(n43480) );
  INV_X1 U25120 ( .A(n43490), .ZN(n27674) );
  AOI221_X1 U25121 ( .B1(n19859), .B2(n26537), .C1(N7322), .C2(n20521), .A(
        n19164), .ZN(n43490) );
  INV_X1 U25122 ( .A(n43500), .ZN(n27675) );
  AOI221_X1 U25123 ( .B1(n19861), .B2(n19268), .C1(N7321), .C2(n24741), .A(
        n25488), .ZN(n43500) );
  INV_X1 U25124 ( .A(n43510), .ZN(n27676) );
  AOI221_X1 U25125 ( .B1(n19863), .B2(n22481), .C1(N7320), .C2(n25958), .A(
        n25489), .ZN(n43510) );
  INV_X1 U25126 ( .A(n43520), .ZN(n27677) );
  AOI221_X1 U25127 ( .B1(n19865), .B2(n22483), .C1(N7319), .C2(n20513), .A(
        n19164), .ZN(n43520) );
  INV_X1 U25128 ( .A(n4323), .ZN(n27666) );
  AOI221_X1 U25129 ( .B1(n19867), .B2(n26672), .C1(N7242), .C2(n25729), .A(
        n25490), .ZN(n4323) );
  INV_X1 U25130 ( .A(n4325), .ZN(n27667) );
  AOI221_X1 U25131 ( .B1(n19869), .B2(n26672), .C1(N7241), .C2(n257301), .A(
        n19165), .ZN(n4325) );
  INV_X1 U25132 ( .A(n4326), .ZN(n27668) );
  AOI221_X1 U25133 ( .B1(n19871), .B2(n20787), .C1(N7240), .C2(n25734), .A(
        n25491), .ZN(n4326) );
  INV_X1 U25134 ( .A(n4327), .ZN(n27669) );
  AOI221_X1 U25135 ( .B1(n19873), .B2(n17087), .C1(N7239), .C2(n21159), .A(
        n25490), .ZN(n4327) );
  INV_X1 U25136 ( .A(n4328), .ZN(n276701) );
  AOI221_X1 U25137 ( .B1(n19875), .B2(n19293), .C1(N7238), .C2(n25716), .A(
        n19165), .ZN(n4328) );
  INV_X1 U25138 ( .A(n4329), .ZN(n27671) );
  AOI221_X1 U25139 ( .B1(n19877), .B2(n19293), .C1(N7237), .C2(n25708), .A(
        n25491), .ZN(n4329) );
  INV_X1 U25140 ( .A(n43010), .ZN(n276601) );
  AOI221_X1 U25141 ( .B1(n19879), .B2(n26718), .C1(N7150), .C2(n20796), .A(
        n25484), .ZN(n43010) );
  INV_X1 U25142 ( .A(n43030), .ZN(n27661) );
  AOI221_X1 U25143 ( .B1(n19881), .B2(n24177), .C1(N7149), .C2(n26650), .A(
        n19162), .ZN(n43030) );
  INV_X1 U25144 ( .A(n43040), .ZN(n27662) );
  AOI221_X1 U25145 ( .B1(n19883), .B2(n25305), .C1(N7148), .C2(n24737), .A(
        n25485), .ZN(n43040) );
  INV_X1 U25146 ( .A(n43050), .ZN(n27663) );
  AOI221_X1 U25147 ( .B1(n19885), .B2(n25307), .C1(N7147), .C2(n19032), .A(
        n25484), .ZN(n43050) );
  INV_X1 U25148 ( .A(n43060), .ZN(n27664) );
  AOI221_X1 U25149 ( .B1(n19887), .B2(n25303), .C1(N7146), .C2(n25742), .A(
        n19162), .ZN(n43060) );
  INV_X1 U25150 ( .A(n43070), .ZN(n27665) );
  AOI221_X1 U25151 ( .B1(n19889), .B2(n26718), .C1(N7145), .C2(n26654), .A(
        n25485), .ZN(n43070) );
  INV_X1 U25152 ( .A(n4279), .ZN(n27654) );
  AOI221_X1 U25153 ( .B1(n19891), .B2(n26753), .C1(N7068), .C2(n21201), .A(
        n25486), .ZN(n4279) );
  INV_X1 U25154 ( .A(n4281), .ZN(n27655) );
  AOI221_X1 U25155 ( .B1(n19893), .B2(n24228), .C1(N7067), .C2(n24550), .A(
        n19163), .ZN(n4281) );
  INV_X1 U25156 ( .A(n4282), .ZN(n27656) );
  AOI221_X1 U25157 ( .B1(n19895), .B2(n25923), .C1(N7066), .C2(n25557), .A(
        n25487), .ZN(n4282) );
  INV_X1 U25158 ( .A(n4283), .ZN(n27657) );
  AOI221_X1 U25159 ( .B1(n19897), .B2(n25913), .C1(N7065), .C2(n24537), .A(
        n25486), .ZN(n4283) );
  INV_X1 U25160 ( .A(n4284), .ZN(n27658) );
  AOI221_X1 U25161 ( .B1(n19899), .B2(n25599), .C1(N7064), .C2(n24558), .A(
        n19163), .ZN(n4284) );
  INV_X1 U25162 ( .A(n4285), .ZN(n27659) );
  AOI221_X1 U25163 ( .B1(n19901), .B2(n26751), .C1(N7063), .C2(n25566), .A(
        n25487), .ZN(n4285) );
  INV_X1 U25164 ( .A(n4162), .ZN(n27624) );
  AOI221_X1 U25165 ( .B1(n19951), .B2(n24989), .C1(N6620), .C2(n19182), .A(
        n25472), .ZN(n4162) );
  INV_X1 U25166 ( .A(n4165), .ZN(n27625) );
  AOI221_X1 U25167 ( .B1(n19953), .B2(n20780), .C1(N6619), .C2(n25717), .A(
        n19156), .ZN(n4165) );
  INV_X1 U25168 ( .A(n4166), .ZN(n27626) );
  AOI221_X1 U25169 ( .B1(n19955), .B2(n24100), .C1(N6618), .C2(n25709), .A(
        n25473), .ZN(n4166) );
  INV_X1 U25170 ( .A(n4167), .ZN(n27627) );
  AOI221_X1 U25171 ( .B1(n19957), .B2(n24100), .C1(N6617), .C2(n25705), .A(
        n25472), .ZN(n4167) );
  INV_X1 U25172 ( .A(n4168), .ZN(n27628) );
  AOI221_X1 U25173 ( .B1(n19959), .B2(n20788), .C1(N6616), .C2(n25697), .A(
        n19156), .ZN(n4168) );
  INV_X1 U25174 ( .A(n4169), .ZN(n27629) );
  AOI221_X1 U25175 ( .B1(n19961), .B2(n20781), .C1(N6615), .C2(n25713), .A(
        n25473), .ZN(n4169) );
  INV_X1 U25176 ( .A(n41400), .ZN(n27618) );
  AOI221_X1 U25177 ( .B1(n19963), .B2(n19076), .C1(N6538), .C2(n19244), .A(
        n25474), .ZN(n41400) );
  INV_X1 U25178 ( .A(n41420), .ZN(n27619) );
  AOI221_X1 U25179 ( .B1(n19965), .B2(n19077), .C1(N6537), .C2(n24069), .A(
        n19157), .ZN(n41420) );
  INV_X1 U25180 ( .A(n41430), .ZN(n27620) );
  AOI221_X1 U25181 ( .B1(n19967), .B2(n25302), .C1(N6536), .C2(n25006), .A(
        n25475), .ZN(n41430) );
  INV_X1 U25182 ( .A(n41440), .ZN(n27621) );
  AOI221_X1 U25183 ( .B1(n19969), .B2(n25303), .C1(N6535), .C2(n19289), .A(
        n25474), .ZN(n41440) );
  INV_X1 U25184 ( .A(n41450), .ZN(n27622) );
  AOI221_X1 U25185 ( .B1(n19971), .B2(n25306), .C1(N6534), .C2(n24999), .A(
        n19157), .ZN(n41450) );
  INV_X1 U25186 ( .A(n41460), .ZN(n27623) );
  AOI221_X1 U25187 ( .B1(n19973), .B2(n25308), .C1(N6533), .C2(n24078), .A(
        n25475), .ZN(n41460) );
  INV_X1 U25188 ( .A(n4118), .ZN(n27612) );
  AOI221_X1 U25189 ( .B1(n19975), .B2(n25924), .C1(N6449), .C2(n21207), .A(
        n25468), .ZN(n4118) );
  INV_X1 U25190 ( .A(n4120), .ZN(n27613) );
  AOI221_X1 U25191 ( .B1(n19977), .B2(n25914), .C1(N6448), .C2(n19190), .A(
        n19154), .ZN(n4120) );
  INV_X1 U25192 ( .A(n4121), .ZN(n27614) );
  AOI221_X1 U25193 ( .B1(n19979), .B2(n25597), .C1(N6447), .C2(n24555), .A(
        n25469), .ZN(n4121) );
  INV_X1 U25194 ( .A(n4122), .ZN(n27615) );
  AOI221_X1 U25195 ( .B1(n19981), .B2(n25599), .C1(N6446), .C2(n24553), .A(
        n25468), .ZN(n4122) );
  INV_X1 U25196 ( .A(n4123), .ZN(n27616) );
  AOI221_X1 U25197 ( .B1(n19983), .B2(n25925), .C1(N6445), .C2(n21204), .A(
        n19154), .ZN(n4123) );
  INV_X1 U25198 ( .A(n4124), .ZN(n27617) );
  AOI221_X1 U25199 ( .B1(n19985), .B2(n25915), .C1(N6444), .C2(n19192), .A(
        n25469), .ZN(n4124) );
  INV_X1 U25200 ( .A(n39790), .ZN(n27576) );
  AOI221_X1 U25201 ( .B1(n20047), .B2(n24178), .C1(N5945), .C2(n19033), .A(
        n25455), .ZN(n39790) );
  INV_X1 U25202 ( .A(n3982), .ZN(n27577) );
  AOI221_X1 U25203 ( .B1(n20049), .B2(n25302), .C1(N5944), .C2(n25004), .A(
        n19148), .ZN(n3982) );
  INV_X1 U25204 ( .A(n3983), .ZN(n27578) );
  AOI221_X1 U25205 ( .B1(n20051), .B2(n25305), .C1(N5943), .C2(n17081), .A(
        n25456), .ZN(n3983) );
  INV_X1 U25206 ( .A(n3984), .ZN(n27579) );
  AOI221_X1 U25207 ( .B1(n20053), .B2(n25307), .C1(N5942), .C2(n20801), .A(
        n25455), .ZN(n3984) );
  INV_X1 U25208 ( .A(n3985), .ZN(n27580) );
  AOI221_X1 U25209 ( .B1(n20055), .B2(n26719), .C1(N5941), .C2(n25751), .A(
        n19148), .ZN(n3985) );
  INV_X1 U25210 ( .A(n3986), .ZN(n27581) );
  AOI221_X1 U25211 ( .B1(n20057), .B2(n25301), .C1(N5940), .C2(n24996), .A(
        n25456), .ZN(n3986) );
  INV_X1 U25212 ( .A(n3957), .ZN(n27570) );
  AOI221_X1 U25213 ( .B1(n20059), .B2(n24229), .C1(N5863), .C2(n25176), .A(
        n25457), .ZN(n3957) );
  INV_X1 U25214 ( .A(n3959), .ZN(n27571) );
  AOI221_X1 U25215 ( .B1(n20061), .B2(n25597), .C1(N5862), .C2(n19051), .A(
        n19149), .ZN(n3959) );
  INV_X1 U25216 ( .A(n39600), .ZN(n27572) );
  AOI221_X1 U25217 ( .B1(n20063), .B2(n25926), .C1(N5861), .C2(n22933), .A(
        n25458), .ZN(n39600) );
  INV_X1 U25218 ( .A(n39610), .ZN(n27573) );
  AOI221_X1 U25219 ( .B1(n20065), .B2(n25912), .C1(N5860), .C2(n25181), .A(
        n25457), .ZN(n39610) );
  INV_X1 U25220 ( .A(n39620), .ZN(n27574) );
  AOI221_X1 U25221 ( .B1(n20067), .B2(n24226), .C1(N5859), .C2(n27167), .A(
        n19149), .ZN(n39620) );
  INV_X1 U25222 ( .A(n39630), .ZN(n27575) );
  AOI221_X1 U25223 ( .B1(n20069), .B2(n24229), .C1(N5858), .C2(n19191), .A(
        n25458), .ZN(n39630) );
  INV_X1 U25224 ( .A(n3822), .ZN(n27534) );
  AOI221_X1 U25225 ( .B1(n20131), .B2(n25933), .C1(N5359), .C2(n21211), .A(
        n25445), .ZN(n3822) );
  INV_X1 U25226 ( .A(n3824), .ZN(n27535) );
  AOI221_X1 U25227 ( .B1(n20133), .B2(n25921), .C1(N5358), .C2(n25548), .A(
        n19143), .ZN(n3824) );
  INV_X1 U25228 ( .A(n3825), .ZN(n27536) );
  AOI221_X1 U25229 ( .B1(n20135), .B2(n25601), .C1(N5357), .C2(n24544), .A(
        n25446), .ZN(n3825) );
  INV_X1 U25230 ( .A(n3826), .ZN(n27537) );
  AOI221_X1 U25231 ( .B1(n20137), .B2(n25605), .C1(N5356), .C2(n21218), .A(
        n25445), .ZN(n3826) );
  INV_X1 U25232 ( .A(n3827), .ZN(n27538) );
  AOI221_X1 U25233 ( .B1(n20139), .B2(n25934), .C1(N5355), .C2(n25560), .A(
        n19143), .ZN(n3827) );
  INV_X1 U25234 ( .A(n3828), .ZN(n27539) );
  AOI221_X1 U25235 ( .B1(n20141), .B2(n25922), .C1(N5354), .C2(n19049), .A(
        n25446), .ZN(n3828) );
  INV_X1 U25236 ( .A(n37970), .ZN(n27528) );
  AOI221_X1 U25237 ( .B1(n20143), .B2(n25923), .C1(N5270), .C2(n19197), .A(
        n25439), .ZN(n37970) );
  INV_X1 U25238 ( .A(n38000), .ZN(n27529) );
  AOI221_X1 U25239 ( .B1(n20145), .B2(n25913), .C1(N5269), .C2(n19194), .A(
        n19140), .ZN(n38000) );
  INV_X1 U25240 ( .A(n38010), .ZN(n27530) );
  AOI221_X1 U25241 ( .B1(n20147), .B2(n256001), .C1(N5268), .C2(n25179), .A(
        n25440), .ZN(n38010) );
  INV_X1 U25242 ( .A(n38020), .ZN(n27531) );
  AOI221_X1 U25243 ( .B1(n20149), .B2(n26753), .C1(N5267), .C2(n25167), .A(
        n25439), .ZN(n38020) );
  INV_X1 U25244 ( .A(n38030), .ZN(n27532) );
  AOI221_X1 U25245 ( .B1(n20151), .B2(n25924), .C1(N5266), .C2(n22930), .A(
        n19140), .ZN(n38030) );
  INV_X1 U25246 ( .A(n38040), .ZN(n27533) );
  AOI221_X1 U25247 ( .B1(n20153), .B2(n25912), .C1(N5265), .C2(n27168), .A(
        n25440), .ZN(n38040) );
  INV_X1 U25248 ( .A(n3665), .ZN(n27492) );
  AOI221_X1 U25249 ( .B1(n20215), .B2(n25605), .C1(N4748), .C2(n21192), .A(
        n25427), .ZN(n3665) );
  INV_X1 U25250 ( .A(n36670), .ZN(n27493) );
  AOI221_X1 U25251 ( .B1(n20217), .B2(n267501), .C1(N4747), .C2(n24567), .A(
        n19134), .ZN(n36670) );
  INV_X1 U25252 ( .A(n36680), .ZN(n27494) );
  AOI221_X1 U25253 ( .B1(n20219), .B2(n25932), .C1(N4746), .C2(n25544), .A(
        n25428), .ZN(n36680) );
  INV_X1 U25254 ( .A(n36690), .ZN(n27495) );
  AOI221_X1 U25255 ( .B1(n20221), .B2(n259201), .C1(N4745), .C2(n24542), .A(
        n25427), .ZN(n36690) );
  INV_X1 U25256 ( .A(n36700), .ZN(n27496) );
  AOI221_X1 U25257 ( .B1(n20223), .B2(n24222), .C1(N4744), .C2(n24575), .A(
        n19134), .ZN(n36700) );
  INV_X1 U25258 ( .A(n36710), .ZN(n27497) );
  AOI221_X1 U25259 ( .B1(n20225), .B2(n24225), .C1(N4743), .C2(n25564), .A(
        n25428), .ZN(n36710) );
  INV_X1 U25260 ( .A(n36410), .ZN(n27486) );
  AOI221_X1 U25261 ( .B1(n20227), .B2(n25298), .C1(N4666), .C2(n19031), .A(
        n25429), .ZN(n36410) );
  INV_X1 U25262 ( .A(n3643), .ZN(n27487) );
  AOI221_X1 U25263 ( .B1(n20229), .B2(n25300), .C1(N4665), .C2(n20805), .A(
        n19135), .ZN(n3643) );
  INV_X1 U25264 ( .A(n3644), .ZN(n27488) );
  AOI221_X1 U25265 ( .B1(n20231), .B2(n25296), .C1(N4664), .C2(n19286), .A(
        n25430), .ZN(n3644) );
  INV_X1 U25266 ( .A(n3645), .ZN(n27489) );
  AOI221_X1 U25267 ( .B1(n20233), .B2(n24183), .C1(N4663), .C2(n20807), .A(
        n25429), .ZN(n3645) );
  INV_X1 U25268 ( .A(n3646), .ZN(n27490) );
  AOI221_X1 U25269 ( .B1(n20235), .B2(n19073), .C1(N4662), .C2(n20518), .A(
        n19135), .ZN(n3646) );
  INV_X1 U25270 ( .A(n3647), .ZN(n27491) );
  AOI221_X1 U25271 ( .B1(n20237), .B2(n19074), .C1(N4661), .C2(n20803), .A(
        n25430), .ZN(n3647) );
  INV_X1 U25272 ( .A(n35060), .ZN(n274501) );
  AOI221_X1 U25273 ( .B1(n20299), .B2(n25931), .C1(N4148), .C2(n21198), .A(
        n25417), .ZN(n35060) );
  INV_X1 U25274 ( .A(n35080), .ZN(n27451) );
  AOI221_X1 U25275 ( .B1(n20301), .B2(n25919), .C1(N4147), .C2(n19186), .A(
        n19129), .ZN(n35080) );
  INV_X1 U25276 ( .A(n35090), .ZN(n27452) );
  AOI221_X1 U25277 ( .B1(n20303), .B2(n24225), .C1(N4146), .C2(n24572), .A(
        n25418), .ZN(n35090) );
  INV_X1 U25278 ( .A(n35100), .ZN(n27453) );
  AOI221_X1 U25279 ( .B1(n20305), .B2(n25602), .C1(N4145), .C2(n24570), .A(
        n25417), .ZN(n35100) );
  INV_X1 U25280 ( .A(n35110), .ZN(n27454) );
  AOI221_X1 U25281 ( .B1(n20307), .B2(n25934), .C1(N4144), .C2(n21195), .A(
        n19129), .ZN(n35110) );
  INV_X1 U25282 ( .A(n35120), .ZN(n27455) );
  AOI221_X1 U25283 ( .B1(n20309), .B2(n25922), .C1(N4143), .C2(n19188), .A(
        n25418), .ZN(n35120) );
  INV_X1 U25284 ( .A(n3484), .ZN(n27444) );
  AOI221_X1 U25285 ( .B1(n20311), .B2(n26721), .C1(N4059), .C2(n25109), .A(
        n25411), .ZN(n3484) );
  INV_X1 U25286 ( .A(n3486), .ZN(n27445) );
  AOI221_X1 U25287 ( .B1(n20313), .B2(n24182), .C1(N4058), .C2(n26649), .A(
        n19126), .ZN(n3486) );
  INV_X1 U25288 ( .A(n3487), .ZN(n27446) );
  AOI221_X1 U25289 ( .B1(n20315), .B2(n25297), .C1(N4057), .C2(n25737), .A(
        n25412), .ZN(n3487) );
  INV_X1 U25290 ( .A(n3488), .ZN(n27447) );
  AOI221_X1 U25291 ( .B1(n20317), .B2(n25299), .C1(N4056), .C2(n25738), .A(
        n25411), .ZN(n3488) );
  INV_X1 U25292 ( .A(n3489), .ZN(n27448) );
  AOI221_X1 U25293 ( .B1(n20319), .B2(n25295), .C1(N4055), .C2(n257401), .A(
        n19126), .ZN(n3489) );
  INV_X1 U25294 ( .A(n3490), .ZN(n27449) );
  AOI221_X1 U25295 ( .B1(n20321), .B2(n26721), .C1(N4054), .C2(n26648), .A(
        n25412), .ZN(n3490) );
  INV_X1 U25296 ( .A(n34590), .ZN(n27438) );
  AOI221_X1 U25297 ( .B1(n20323), .B2(n20783), .C1(N3980), .C2(n25691), .A(
        n25413), .ZN(n34590) );
  INV_X1 U25298 ( .A(n34610), .ZN(n27439) );
  AOI221_X1 U25299 ( .B1(n20325), .B2(n20774), .C1(N3979), .C2(n25683), .A(
        n19127), .ZN(n34610) );
  INV_X1 U25300 ( .A(n34620), .ZN(n274401) );
  AOI221_X1 U25301 ( .B1(n20327), .B2(n22753), .C1(N3978), .C2(n257001), .A(
        n25414), .ZN(n34620) );
  INV_X1 U25302 ( .A(n34630), .ZN(n27441) );
  AOI221_X1 U25303 ( .B1(n20329), .B2(n22752), .C1(N3977), .C2(n25724), .A(
        n25413), .ZN(n34630) );
  INV_X1 U25304 ( .A(n34640), .ZN(n27442) );
  AOI221_X1 U25305 ( .B1(n20331), .B2(n17088), .C1(N3976), .C2(n257201), .A(
        n19127), .ZN(n34640) );
  INV_X1 U25306 ( .A(n34650), .ZN(n27443) );
  AOI221_X1 U25307 ( .B1(n20333), .B2(n24985), .C1(N3975), .C2(n25725), .A(
        n25414), .ZN(n34650) );
  INV_X1 U25308 ( .A(n33460), .ZN(n27408) );
  AOI221_X1 U25309 ( .B1(matrix_mul_2D_1__3__20_), .B2(n25602), .C1(N3552), 
        .C2(n25174), .A(n25399), .ZN(n33460) );
  INV_X1 U25310 ( .A(n3348), .ZN(n27409) );
  AOI221_X1 U25311 ( .B1(matrix_mul_2D_1__3__19_), .B2(n25604), .C1(N3551), 
        .C2(n19048), .A(n19120), .ZN(n3348) );
  INV_X1 U25312 ( .A(n3349), .ZN(n274101) );
  AOI221_X1 U25313 ( .B1(matrix_mul_2D_1__3__18_), .B2(n25933), .C1(N3550), 
        .C2(n22939), .A(n25400), .ZN(n3349) );
  INV_X1 U25314 ( .A(n3350), .ZN(n27411) );
  AOI221_X1 U25315 ( .B1(matrix_mul_2D_1__3__17_), .B2(n25921), .C1(N3549), 
        .C2(n25171), .A(n25399), .ZN(n3350) );
  INV_X1 U25316 ( .A(n3351), .ZN(n27412) );
  AOI221_X1 U25317 ( .B1(matrix_mul_2D_1__3__16_), .B2(n25604), .C1(N3548), 
        .C2(n27255), .A(n19120), .ZN(n3351) );
  INV_X1 U25318 ( .A(n3352), .ZN(n27413) );
  AOI221_X1 U25319 ( .B1(matrix_mul_2D_1__3__15_), .B2(n26748), .C1(N3547), 
        .C2(n19187), .A(n25400), .ZN(n3352) );
  INV_X1 U25320 ( .A(n3324), .ZN(n27402) );
  AOI221_X1 U25321 ( .B1(matrix_mul_2D_1__2__20_), .B2(n19073), .C1(N3473), 
        .C2(n25103), .A(n25401), .ZN(n3324) );
  INV_X1 U25322 ( .A(n3326), .ZN(n27403) );
  AOI221_X1 U25323 ( .B1(matrix_mul_2D_1__2__19_), .B2(n19074), .C1(N3472), 
        .C2(n24064), .A(n19121), .ZN(n3326) );
  INV_X1 U25324 ( .A(n3327), .ZN(n27404) );
  AOI221_X1 U25325 ( .B1(matrix_mul_2D_1__2__18_), .B2(n25294), .C1(N3471), 
        .C2(n22714), .A(n25402), .ZN(n3327) );
  INV_X1 U25326 ( .A(n3328), .ZN(n27405) );
  AOI221_X1 U25327 ( .B1(matrix_mul_2D_1__2__17_), .B2(n25295), .C1(N3470), 
        .C2(n19285), .A(n25401), .ZN(n3328) );
  INV_X1 U25328 ( .A(n3329), .ZN(n27406) );
  AOI221_X1 U25329 ( .B1(matrix_mul_2D_1__2__16_), .B2(n25298), .C1(N3469), 
        .C2(n25736), .A(n19121), .ZN(n3329) );
  INV_X1 U25330 ( .A(n3330), .ZN(n27407) );
  AOI221_X1 U25331 ( .B1(matrix_mul_2D_1__2__15_), .B2(n25300), .C1(N3468), 
        .C2(n24059), .A(n25402), .ZN(n3330) );
  INV_X1 U25332 ( .A(n33020), .ZN(n27396) );
  AOI221_X1 U25333 ( .B1(n20359), .B2(n26673), .C1(N3384), .C2(n25721), .A(
        n25395), .ZN(n33020) );
  INV_X1 U25334 ( .A(n33040), .ZN(n27397) );
  AOI221_X1 U25335 ( .B1(n20361), .B2(n26673), .C1(N3383), .C2(n25722), .A(
        n19118), .ZN(n33040) );
  INV_X1 U25336 ( .A(n33050), .ZN(n27398) );
  AOI221_X1 U25337 ( .B1(n20363), .B2(n20783), .C1(N3382), .C2(n25726), .A(
        n25396), .ZN(n33050) );
  INV_X1 U25338 ( .A(n3306), .ZN(n27399) );
  AOI221_X1 U25339 ( .B1(n20365), .B2(n24985), .C1(N3381), .C2(n21153), .A(
        n25395), .ZN(n3306) );
  INV_X1 U25340 ( .A(n3307), .ZN(n274001) );
  AOI221_X1 U25341 ( .B1(n20367), .B2(n19294), .C1(N3380), .C2(n25687), .A(
        n19118), .ZN(n3307) );
  INV_X1 U25342 ( .A(n3308), .ZN(n27401) );
  AOI221_X1 U25343 ( .B1(n20369), .B2(n19294), .C1(N3379), .C2(n25678), .A(
        n25396), .ZN(n3308) );
  INV_X1 U25344 ( .A(n3277), .ZN(n273901) );
  AOI221_X1 U25345 ( .B1(n20371), .B2(n26539), .C1(N3305), .C2(n19243), .A(
        n25397), .ZN(n3277) );
  INV_X1 U25346 ( .A(n3279), .ZN(n27391) );
  AOI221_X1 U25347 ( .B1(n20373), .B2(n19269), .C1(N3304), .C2(n21445), .A(
        n19119), .ZN(n3279) );
  INV_X1 U25348 ( .A(n3280), .ZN(n27392) );
  AOI221_X1 U25349 ( .B1(n20375), .B2(n22486), .C1(N3303), .C2(n20531), .A(
        n25398), .ZN(n3280) );
  INV_X1 U25350 ( .A(n3281), .ZN(n27393) );
  AOI221_X1 U25351 ( .B1(n20377), .B2(n22489), .C1(N3302), .C2(n24739), .A(
        n25397), .ZN(n3281) );
  INV_X1 U25352 ( .A(n3282), .ZN(n27394) );
  AOI221_X1 U25353 ( .B1(n20379), .B2(n26538), .C1(N3301), .C2(n21441), .A(
        n19119), .ZN(n3282) );
  INV_X1 U25354 ( .A(n3283), .ZN(n27395) );
  AOI221_X1 U25355 ( .B1(n20381), .B2(n22490), .C1(N3300), .C2(n25967), .A(
        n25398), .ZN(n3283) );
  INV_X1 U25356 ( .A(n31770), .ZN(n27366) );
  AOI221_X1 U25357 ( .B1(n20419), .B2(n25932), .C1(N2960), .C2(n19195), .A(
        n25389), .ZN(n31770) );
  INV_X1 U25358 ( .A(n3180), .ZN(n27367) );
  AOI221_X1 U25359 ( .B1(n20421), .B2(n259201), .C1(N2959), .C2(n19193), .A(
        n19115), .ZN(n3180) );
  INV_X1 U25360 ( .A(n3181), .ZN(n27368) );
  AOI221_X1 U25361 ( .B1(n20423), .B2(n267501), .C1(N2958), .C2(n25177), .A(
        n25390), .ZN(n3181) );
  INV_X1 U25362 ( .A(n3182), .ZN(n27369) );
  AOI221_X1 U25363 ( .B1(n20425), .B2(n24224), .C1(N2957), .C2(n25163), .A(
        n25389), .ZN(n3182) );
  INV_X1 U25364 ( .A(n3183), .ZN(n273701) );
  AOI221_X1 U25365 ( .B1(n20427), .B2(n25931), .C1(N2956), .C2(n22936), .A(
        n19115), .ZN(n3183) );
  INV_X1 U25366 ( .A(n3184), .ZN(n27371) );
  AOI221_X1 U25367 ( .B1(n20429), .B2(n25919), .C1(N2955), .C2(n27256), .A(
        n25390), .ZN(n3184) );
  INV_X1 U25368 ( .A(n3152), .ZN(n273601) );
  AOI221_X1 U25369 ( .B1(n20431), .B2(n24183), .C1(N2868), .C2(n19284), .A(
        n25383), .ZN(n3152) );
  INV_X1 U25370 ( .A(n3155), .ZN(n27361) );
  AOI221_X1 U25371 ( .B1(n20433), .B2(n25294), .C1(N2867), .C2(n25010), .A(
        n19112), .ZN(n3155) );
  INV_X1 U25372 ( .A(n3156), .ZN(n27362) );
  AOI221_X1 U25373 ( .B1(n20435), .B2(n25297), .C1(N2866), .C2(n19027), .A(
        n25384), .ZN(n3156) );
  INV_X1 U25374 ( .A(n3157), .ZN(n27363) );
  AOI221_X1 U25375 ( .B1(n20437), .B2(n25299), .C1(N2865), .C2(n27261), .A(
        n25383), .ZN(n3157) );
  INV_X1 U25376 ( .A(n3158), .ZN(n27364) );
  AOI221_X1 U25377 ( .B1(n20439), .B2(n26722), .C1(N2864), .C2(n24733), .A(
        n19112), .ZN(n3158) );
  INV_X1 U25378 ( .A(n3159), .ZN(n27365) );
  AOI221_X1 U25379 ( .B1(n20441), .B2(n25293), .C1(N2863), .C2(n25008), .A(
        n25384), .ZN(n3159) );
  INV_X1 U25380 ( .A(n31270), .ZN(n27354) );
  AOI221_X1 U25381 ( .B1(n20443), .B2(n17088), .C1(N2786), .C2(n19180), .A(
        n25385), .ZN(n31270) );
  INV_X1 U25382 ( .A(n31300), .ZN(n27355) );
  AOI221_X1 U25383 ( .B1(n20445), .B2(n20774), .C1(N2785), .C2(n25688), .A(
        n19113), .ZN(n31300) );
  INV_X1 U25384 ( .A(n31310), .ZN(n27356) );
  AOI221_X1 U25385 ( .B1(n20447), .B2(n24102), .C1(N2784), .C2(n25679), .A(
        n25386), .ZN(n31310) );
  INV_X1 U25386 ( .A(n31320), .ZN(n27357) );
  AOI221_X1 U25387 ( .B1(n20449), .B2(n24102), .C1(N2783), .C2(n25692), .A(
        n25385), .ZN(n31320) );
  INV_X1 U25388 ( .A(n31330), .ZN(n27358) );
  AOI221_X1 U25389 ( .B1(n20451), .B2(n20784), .C1(N2782), .C2(n25684), .A(
        n19113), .ZN(n31330) );
  INV_X1 U25390 ( .A(n31340), .ZN(n27359) );
  AOI221_X1 U25391 ( .B1(n20453), .B2(n20775), .C1(N2781), .C2(n25701), .A(
        n25386), .ZN(n31340) );
  INV_X1 U25392 ( .A(n3102), .ZN(n27348) );
  AOI221_X1 U25393 ( .B1(n20455), .B2(n22486), .C1(N2694), .C2(n25968), .A(
        n25379), .ZN(n3102) );
  INV_X1 U25394 ( .A(n3105), .ZN(n27349) );
  AOI221_X1 U25395 ( .B1(n20457), .B2(n22490), .C1(N2693), .C2(n17101), .A(
        n25380), .ZN(n3105) );
  INV_X1 U25396 ( .A(n3106), .ZN(n273501) );
  AOI221_X1 U25397 ( .B1(n20459), .B2(n26539), .C1(N2692), .C2(n20516), .A(
        n19110), .ZN(n3106) );
  INV_X1 U25398 ( .A(n3107), .ZN(n27351) );
  AOI221_X1 U25399 ( .B1(n20461), .B2(n19269), .C1(N2691), .C2(n24743), .A(
        n25379), .ZN(n3107) );
  INV_X1 U25400 ( .A(n3108), .ZN(n27352) );
  AOI221_X1 U25401 ( .B1(n20463), .B2(n22487), .C1(N2690), .C2(n25961), .A(
        n25380), .ZN(n3108) );
  INV_X1 U25402 ( .A(n3109), .ZN(n27353) );
  AOI221_X1 U25403 ( .B1(n20465), .B2(n22489), .C1(N2689), .C2(n20509), .A(
        n19110), .ZN(n3109) );
  INV_X1 U25404 ( .A(n3070), .ZN(n27342) );
  AOI221_X1 U25405 ( .B1(n20467), .B2(n25117), .C1(N2612), .C2(n21392), .A(
        n25381), .ZN(n3070) );
  INV_X1 U25406 ( .A(n3073), .ZN(n27343) );
  AOI221_X1 U25407 ( .B1(n20469), .B2(n19035), .C1(N2611), .C2(n21395), .A(
        n19111), .ZN(n3073) );
  INV_X1 U25408 ( .A(n3074), .ZN(n27344) );
  AOI221_X1 U25409 ( .B1(n20471), .B2(n25118), .C1(N2610), .C2(n21385), .A(
        n25382), .ZN(n3074) );
  INV_X1 U25410 ( .A(n3075), .ZN(n27345) );
  AOI221_X1 U25411 ( .B1(n20473), .B2(n25117), .C1(N2609), .C2(n19240), .A(
        n25381), .ZN(n3075) );
  INV_X1 U25412 ( .A(n3076), .ZN(n27346) );
  AOI221_X1 U25413 ( .B1(n20475), .B2(n19035), .C1(N2608), .C2(n19241), .A(
        n19111), .ZN(n3076) );
  INV_X1 U25414 ( .A(n3077), .ZN(n27347) );
  AOI221_X1 U25415 ( .B1(n20477), .B2(n25118), .C1(N2607), .C2(n19239), .A(
        n25382), .ZN(n3077) );
  INV_X1 U25416 ( .A(n50960), .ZN(n27785) );
  AOI22_X1 U25417 ( .A1(n17899), .A2(n21509), .B1(n17923), .B2(n26326), .ZN(
        n50960) );
  INV_X1 U25418 ( .A(n50920), .ZN(n27784) );
  AOI22_X1 U25419 ( .A1(n17897), .A2(n21511), .B1(n17921), .B2(n21873), .ZN(
        n50920) );
  INV_X1 U25420 ( .A(n5100), .ZN(n27786) );
  AOI22_X1 U25421 ( .A1(n17901), .A2(n26084), .B1(n17925), .B2(n26328), .ZN(
        n5100) );
  INV_X1 U25422 ( .A(n5104), .ZN(n27787) );
  AOI22_X1 U25423 ( .A1(n17903), .A2(n26085), .B1(n17927), .B2(n26327), .ZN(
        n5104) );
  INV_X1 U25424 ( .A(n47970), .ZN(n27762) );
  AOI22_X1 U25425 ( .A1(n17707), .A2(n26148), .B1(n17695), .B2(n26373), .ZN(
        n47970) );
  INV_X1 U25426 ( .A(n47930), .ZN(n27761) );
  AOI22_X1 U25427 ( .A1(n17705), .A2(n21630), .B1(n17693), .B2(n21945), .ZN(
        n47930) );
  INV_X1 U25428 ( .A(n4786), .ZN(n277601) );
  AOI22_X1 U25429 ( .A1(n17703), .A2(n21631), .B1(n17691), .B2(n18431), .ZN(
        n4786) );
  INV_X1 U25430 ( .A(n48010), .ZN(n27763) );
  AOI22_X1 U25431 ( .A1(n17709), .A2(n26147), .B1(n17697), .B2(n26376), .ZN(
        n48010) );
  INV_X1 U25432 ( .A(n4809), .ZN(n27764) );
  AOI22_X1 U25433 ( .A1(n17711), .A2(n26148), .B1(n17699), .B2(n26375), .ZN(
        n4809) );
  INV_X1 U25434 ( .A(n4813), .ZN(n27765) );
  AOI22_X1 U25435 ( .A1(n17713), .A2(n21629), .B1(n17701), .B2(n21945), .ZN(
        n4813) );
  INV_X1 U25436 ( .A(n552), .ZN(n27301) );
  INV_X1 U25437 ( .A(n454), .ZN(n27300) );
  OAI21_X1 U25438 ( .B1(n20885), .B2(n18514), .A(n27305), .ZN(r899_B_2_) );
  INV_X1 U25439 ( .A(n467), .ZN(n27302) );
  OAI21_X1 U25440 ( .B1(n22952), .B2(n27303), .A(n27304), .ZN(r899_B_1_) );
  INV_X1 U25441 ( .A(n455), .ZN(n27303) );
  AOI21_X1 U25442 ( .B1(n876), .B2(n543), .A(n20886), .ZN(n4029) );
  AOI221_X1 U25443 ( .B1(n25941), .B2(matrix_mul_2D_0__4__0_), .C1(
        matrix_mul_2D_0__3__0_), .C2(n25315), .A(n54210), .ZN(n54200) );
  OAI22_X1 U25444 ( .A1(n1970), .A2(n22745), .B1(n1940), .B2(n19283), .ZN(
        n54210) );
  AOI221_X1 U25445 ( .B1(n25951), .B2(matrix_mul_2D_0__4__1_), .C1(
        matrix_mul_2D_0__3__1_), .C2(n21023), .A(n50880), .ZN(n50870) );
  OAI22_X1 U25446 ( .A1(n1969), .A2(n24099), .B1(n1939), .B2(n24051), .ZN(
        n50880) );
  AOI221_X1 U25447 ( .B1(n259401), .B2(matrix_mul_2D_0__4__2_), .C1(
        matrix_mul_2D_0__3__2_), .C2(n25311), .A(n5042), .ZN(n5041) );
  OAI22_X1 U25448 ( .A1(n1968), .A2(n24987), .B1(n1938), .B2(n24054), .ZN(
        n5042) );
  AOI221_X1 U25449 ( .B1(n25952), .B2(matrix_mul_2D_0__4__3_), .C1(
        matrix_mul_2D_0__3__3_), .C2(n25313), .A(n49980), .ZN(n49970) );
  OAI22_X1 U25450 ( .A1(n1967), .A2(n22744), .B1(n1937), .B2(n26645), .ZN(
        n49980) );
  AOI221_X1 U25451 ( .B1(n25944), .B2(matrix_mul_2D_0__4__4_), .C1(
        matrix_mul_2D_0__3__4_), .C2(n22795), .A(n4946), .ZN(n4945) );
  OAI22_X1 U25452 ( .A1(n1966), .A2(n26671), .B1(n1936), .B2(n22712), .ZN(
        n4946) );
  AOI221_X1 U25453 ( .B1(n25937), .B2(matrix_mul_2D_0__4__5_), .C1(
        matrix_mul_2D_0__3__5_), .C2(n25314), .A(n49020), .ZN(n4901) );
  OAI22_X1 U25454 ( .A1(n1965), .A2(n19292), .B1(n1935), .B2(n26645), .ZN(
        n49020) );
  AOI221_X1 U25455 ( .B1(n259501), .B2(matrix_mul_2D_0__4__6_), .C1(
        matrix_mul_2D_0__3__6_), .C2(n22794), .A(n4851), .ZN(n4850) );
  OAI22_X1 U25456 ( .A1(n1964), .A2(n24098), .B1(n1934), .B2(n24052), .ZN(
        n4851) );
  AOI221_X1 U25457 ( .B1(n17126), .B2(matrix_mul_2D_0__4__7_), .C1(
        matrix_mul_2D_0__3__7_), .C2(n26717), .A(n4805), .ZN(n4804) );
  OAI22_X1 U25458 ( .A1(n1963), .A2(n24099), .B1(n1933), .B2(n24051), .ZN(
        n4805) );
  AOI221_X1 U25459 ( .B1(n25938), .B2(matrix_mul_2D_0__4__8_), .C1(
        matrix_mul_2D_0__3__8_), .C2(n22795), .A(n4758), .ZN(n4757) );
  OAI22_X1 U25460 ( .A1(n1962), .A2(n20786), .B1(n1932), .B2(n24055), .ZN(
        n4758) );
  AOI221_X1 U25461 ( .B1(n25951), .B2(matrix_mul_2D_0__4__9_), .C1(
        matrix_mul_2D_0__3__9_), .C2(n19078), .A(n47040), .ZN(n47020) );
  OAI22_X1 U25462 ( .A1(n1961), .A2(n26670), .B1(n1931), .B2(n22711), .ZN(
        n47040) );
  AOI221_X1 U25463 ( .B1(n25939), .B2(matrix_mul_2D_0__4__10_), .C1(
        matrix_mul_2D_0__3__10_), .C2(n25315), .A(n5374), .ZN(n5373) );
  OAI22_X1 U25464 ( .A1(n1960), .A2(n24096), .B1(n1930), .B2(n24048), .ZN(
        n5374) );
  AOI221_X1 U25465 ( .B1(n25952), .B2(matrix_mul_2D_0__4__11_), .C1(
        matrix_mul_2D_0__3__11_), .C2(n21024), .A(n5330), .ZN(n5329) );
  OAI22_X1 U25466 ( .A1(n1959), .A2(n24098), .B1(n1929), .B2(n24052), .ZN(
        n5330) );
  AOI221_X1 U25467 ( .B1(n25943), .B2(matrix_mul_2D_0__4__12_), .C1(
        matrix_mul_2D_0__3__12_), .C2(n21024), .A(n5280), .ZN(n5279) );
  OAI22_X1 U25468 ( .A1(n1958), .A2(n24987), .B1(n1928), .B2(n24055), .ZN(
        n5280) );
  AOI221_X1 U25469 ( .B1(n259401), .B2(matrix_mul_2D_0__4__13_), .C1(
        matrix_mul_2D_0__3__13_), .C2(n25309), .A(n5236), .ZN(n5235) );
  OAI22_X1 U25470 ( .A1(n1957), .A2(n20785), .B1(n1927), .B2(n24054), .ZN(
        n5236) );
  AOI221_X1 U25471 ( .B1(n25949), .B2(matrix_mul_2D_0__4__14_), .C1(
        matrix_mul_2D_0__3__14_), .C2(n25312), .A(n51880), .ZN(n51870) );
  OAI22_X1 U25472 ( .A1(n1956), .A2(n26671), .B1(n1926), .B2(n24048), .ZN(
        n51880) );
  AOI221_X1 U25473 ( .B1(n26332), .B2(matrix_mul_2D_1__0__0_), .C1(n21886), 
        .C2(matrix_mul_2D_1__1__0_), .A(n50770), .ZN(n50760) );
  OAI22_X1 U25474 ( .A1(n2042), .A2(n21247), .B1(n2021), .B2(n21244), .ZN(
        n50770) );
  AOI221_X1 U25475 ( .B1(n26330), .B2(matrix_mul_2D_1__0__1_), .C1(n26335), 
        .C2(matrix_mul_2D_1__1__1_), .A(n5073), .ZN(n5072) );
  OAI22_X1 U25476 ( .A1(n2041), .A2(n21249), .B1(n2020), .B2(n21233), .ZN(
        n5073) );
  AOI221_X1 U25477 ( .B1(n26108), .B2(matrix_mul_2D_1__0__2_), .C1(n21539), 
        .C2(matrix_mul_2D_1__1__2_), .A(n5069), .ZN(n5068) );
  OAI22_X1 U25478 ( .A1(n2040), .A2(n21240), .B1(n2019), .B2(n21236), .ZN(
        n5069) );
  AOI221_X1 U25479 ( .B1(n21552), .B2(matrix_mul_2D_1__0__3_), .C1(n261001), 
        .C2(matrix_mul_2D_1__1__3_), .A(n5065), .ZN(n5064) );
  OAI22_X1 U25480 ( .A1(n2039), .A2(n25574), .B1(n2018), .B2(n25573), .ZN(
        n5065) );
  AOI221_X1 U25481 ( .B1(n26331), .B2(matrix_mul_2D_1__0__4_), .C1(n26335), 
        .C2(matrix_mul_2D_1__1__4_), .A(n5061), .ZN(n5060) );
  OAI22_X1 U25482 ( .A1(n2038), .A2(n25575), .B1(n2017), .B2(n21244), .ZN(
        n5061) );
  AOI221_X1 U25483 ( .B1(n21878), .B2(matrix_mul_2D_1__0__5_), .C1(n26334), 
        .C2(matrix_mul_2D_1__1__5_), .A(n50570), .ZN(n50560) );
  OAI22_X1 U25484 ( .A1(n2037), .A2(n19202), .B1(n2016), .B2(n19201), .ZN(
        n50570) );
  AOI221_X1 U25485 ( .B1(n26108), .B2(matrix_mul_2D_1__0__6_), .C1(n21541), 
        .C2(matrix_mul_2D_1__1__6_), .A(n50530), .ZN(n50520) );
  OAI22_X1 U25486 ( .A1(n2036), .A2(n25574), .B1(n2015), .B2(n25573), .ZN(
        n50530) );
  AOI221_X1 U25487 ( .B1(n21553), .B2(matrix_mul_2D_1__0__7_), .C1(n21540), 
        .C2(matrix_mul_2D_1__1__7_), .A(n50490), .ZN(n50480) );
  OAI22_X1 U25488 ( .A1(n2035), .A2(n25575), .B1(n2014), .B2(n21237), .ZN(
        n50490) );
  AOI221_X1 U25489 ( .B1(n21877), .B2(matrix_mul_2D_1__0__8_), .C1(n21885), 
        .C2(matrix_mul_2D_1__1__8_), .A(n50450), .ZN(n50440) );
  OAI22_X1 U25490 ( .A1(n2034), .A2(n25571), .B1(n2013), .B2(n25570), .ZN(
        n50450) );
  AOI221_X1 U25491 ( .B1(n21880), .B2(matrix_mul_2D_1__0__9_), .C1(n21882), 
        .C2(matrix_mul_2D_1__1__9_), .A(n5037), .ZN(n5036) );
  OAI22_X1 U25492 ( .A1(n2033), .A2(n19203), .B1(n2012), .B2(n21233), .ZN(
        n5037) );
  AOI221_X1 U25493 ( .B1(n21551), .B2(matrix_mul_2D_1__0__10_), .C1(n21538), 
        .C2(matrix_mul_2D_1__1__10_), .A(n5033), .ZN(n5032) );
  OAI22_X1 U25494 ( .A1(n2032), .A2(n21249), .B1(n2011), .B2(n21232), .ZN(
        n5033) );
  AOI221_X1 U25495 ( .B1(n26107), .B2(matrix_mul_2D_1__0__11_), .C1(n26101), 
        .C2(matrix_mul_2D_1__1__11_), .A(n5029), .ZN(n5028) );
  OAI22_X1 U25496 ( .A1(n2031), .A2(n25571), .B1(n2010), .B2(n25570), .ZN(
        n5029) );
  AOI221_X1 U25497 ( .B1(n21881), .B2(matrix_mul_2D_1__0__12_), .C1(n21883), 
        .C2(matrix_mul_2D_1__1__12_), .A(n5025), .ZN(n5024) );
  OAI22_X1 U25498 ( .A1(n2030), .A2(n21246), .B1(n2009), .B2(n21243), .ZN(
        n5025) );
  AOI221_X1 U25499 ( .B1(n26332), .B2(matrix_mul_2D_1__0__13_), .C1(n26333), 
        .C2(matrix_mul_2D_1__1__13_), .A(n5021), .ZN(n5020) );
  OAI22_X1 U25500 ( .A1(n2029), .A2(n19204), .B1(n2008), .B2(n19200), .ZN(
        n5021) );
  AOI221_X1 U25501 ( .B1(n21554), .B2(matrix_mul_2D_1__0__14_), .C1(n26101), 
        .C2(matrix_mul_2D_1__1__14_), .A(n5017), .ZN(n5016) );
  OAI22_X1 U25502 ( .A1(n2028), .A2(n21239), .B1(n2007), .B2(n21237), .ZN(
        n5017) );
  OAI22_X1 U25503 ( .A1(n28520), .A2(n25525), .B1(n2837), .B2(n20753), .ZN(
        n5202) );
  OAI22_X1 U25504 ( .A1(n28510), .A2(n24639), .B1(n2836), .B2(n20746), .ZN(
        n5196) );
  OAI22_X1 U25505 ( .A1(n28500), .A2(n24633), .B1(n2835), .B2(n24968), .ZN(
        n5192) );
  OAI22_X1 U25506 ( .A1(n28490), .A2(n25668), .B1(n2834), .B2(n24141), .ZN(
        n51840) );
  OAI22_X1 U25507 ( .A1(n28480), .A2(n256701), .B1(n2833), .B2(n24973), .ZN(
        n51800) );
  OAI22_X1 U25508 ( .A1(n2847), .A2(n25669), .B1(n2832), .B2(n26676), .ZN(
        n51760) );
  OAI22_X1 U25509 ( .A1(n2846), .A2(n25671), .B1(n2831), .B2(n22757), .ZN(
        n51720) );
  OAI22_X1 U25510 ( .A1(n2845), .A2(n24632), .B1(n28300), .B2(n24141), .ZN(
        n51680) );
  OAI22_X1 U25511 ( .A1(n2844), .A2(n24638), .B1(n28290), .B2(n20752), .ZN(
        n5164) );
  OAI22_X1 U25512 ( .A1(n2843), .A2(n24635), .B1(n28280), .B2(n19295), .ZN(
        n5160) );
  OAI22_X1 U25513 ( .A1(n2842), .A2(n24636), .B1(n28270), .B2(n20747), .ZN(
        n5156) );
  OAI22_X1 U25514 ( .A1(n2841), .A2(n25666), .B1(n28260), .B2(n26677), .ZN(
        n5152) );
  OAI22_X1 U25515 ( .A1(n2840), .A2(n25672), .B1(n28250), .B2(n22756), .ZN(
        n51480) );
  OAI22_X1 U25516 ( .A1(n2839), .A2(n25667), .B1(n28240), .B2(n24973), .ZN(
        n51400) );
  OAI22_X1 U25517 ( .A1(n2838), .A2(n25673), .B1(n28230), .B2(n24968), .ZN(
        n5134) );
  OAI22_X1 U25518 ( .A1(n2588), .A2(n26517), .B1(n257300), .B2(n26678), .ZN(
        n53940) );
  OAI22_X1 U25519 ( .A1(n2581), .A2(n22948), .B1(n256600), .B2(n20744), .ZN(
        n5362) );
  OAI22_X1 U25520 ( .A1(n2580), .A2(n23450), .B1(n256500), .B2(n20748), .ZN(
        n53580) );
  OAI22_X1 U25521 ( .A1(n257400), .A2(n22466), .B1(n255900), .B2(n22760), .ZN(
        n5334) );
  OAI22_X1 U25522 ( .A1(n2587), .A2(n22450), .B1(n257200), .B2(n20740), .ZN(
        n53900) );
  OAI22_X1 U25523 ( .A1(n2586), .A2(n24662), .B1(n257100), .B2(n26683), .ZN(
        n53860) );
  OAI22_X1 U25524 ( .A1(n2585), .A2(n26519), .B1(n257000), .B2(n25347), .ZN(
        n5382) );
  OAI22_X1 U25525 ( .A1(n2583), .A2(n22462), .B1(n256800), .B2(n25345), .ZN(
        n5370) );
  OAI22_X1 U25526 ( .A1(n2579), .A2(n24655), .B1(n256400), .B2(n20742), .ZN(
        n53540) );
  OAI22_X1 U25527 ( .A1(n2578), .A2(n24668), .B1(n256300), .B2(n19177), .ZN(
        n53500) );
  OAI22_X1 U25528 ( .A1(n2577), .A2(n22453), .B1(n256200), .B2(n22762), .ZN(
        n53460) );
  OAI22_X1 U25529 ( .A1(n2575), .A2(n22949), .B1(n256000), .B2(n19179), .ZN(
        n5338) );
  OAI22_X1 U25530 ( .A1(n2584), .A2(n26525), .B1(n256900), .B2(n21141), .ZN(
        n5378) );
  OAI22_X1 U25531 ( .A1(n2582), .A2(n22465), .B1(n256700), .B2(n21151), .ZN(
        n5366) );
  OAI22_X1 U25532 ( .A1(n2576), .A2(n23451), .B1(n256100), .B2(n25520), .ZN(
        n53420) );
  OAI22_X1 U25533 ( .A1(n2462), .A2(n24961), .B1(n2447), .B2(n22509), .ZN(
        n4782) );
  OAI22_X1 U25534 ( .A1(n2461), .A2(n25094), .B1(n2446), .B2(n22510), .ZN(
        n4778) );
  OAI22_X1 U25535 ( .A1(n2460), .A2(n25093), .B1(n2445), .B2(n22506), .ZN(
        n4774) );
  OAI22_X1 U25536 ( .A1(n2459), .A2(n26681), .B1(n2444), .B2(n26533), .ZN(
        n4770) );
  OAI22_X1 U25537 ( .A1(n2458), .A2(n25522), .B1(n2443), .B2(n26522), .ZN(
        n4766) );
  OAI22_X1 U25538 ( .A1(n2457), .A2(n24966), .B1(n2442), .B2(n23686), .ZN(
        n4762) );
  OAI22_X1 U25539 ( .A1(n2456), .A2(n24965), .B1(n2441), .B2(n22474), .ZN(
        n4754) );
  OAI22_X1 U25540 ( .A1(n2455), .A2(n26685), .B1(n2440), .B2(n22503), .ZN(
        n4750) );
  OAI22_X1 U25541 ( .A1(n2454), .A2(n24963), .B1(n2439), .B2(n26554), .ZN(
        n47460) );
  OAI22_X1 U25542 ( .A1(n2453), .A2(n25344), .B1(n2438), .B2(n26535), .ZN(
        n47420) );
  OAI22_X1 U25543 ( .A1(n2452), .A2(n24959), .B1(n2437), .B2(n22456), .ZN(
        n47380) );
  OAI22_X1 U25544 ( .A1(n2451), .A2(n19092), .B1(n2436), .B2(n22477), .ZN(
        n47340) );
  OAI22_X1 U25545 ( .A1(n2450), .A2(n21147), .B1(n2435), .B2(n26524), .ZN(
        n47300) );
  OAI22_X1 U25546 ( .A1(n2449), .A2(n24970), .B1(n2434), .B2(n22459), .ZN(
        n4726) );
  OAI22_X1 U25547 ( .A1(n2448), .A2(n25516), .B1(n2433), .B2(n23680), .ZN(
        n4720) );
  OAI22_X1 U25548 ( .A1(n2084), .A2(n21259), .B1(n2063), .B2(n21222), .ZN(
        n50800) );
  OAI22_X1 U25549 ( .A1(n2083), .A2(n21267), .B1(n2062), .B2(n21230), .ZN(
        n5074) );
  OAI22_X1 U25550 ( .A1(n2082), .A2(n21265), .B1(n2061), .B2(n21227), .ZN(
        n5070) );
  OAI22_X1 U25551 ( .A1(n2081), .A2(n25582), .B1(n2060), .B2(n25565), .ZN(
        n5066) );
  OAI22_X1 U25552 ( .A1(n2080), .A2(n25585), .B1(n2059), .B2(n25568), .ZN(
        n5062) );
  OAI22_X1 U25553 ( .A1(n2079), .A2(n19208), .B1(n2058), .B2(n19198), .ZN(
        n50580) );
  OAI22_X1 U25554 ( .A1(n2078), .A2(n25582), .B1(n2057), .B2(n25565), .ZN(
        n50540) );
  OAI22_X1 U25555 ( .A1(n2077), .A2(n25585), .B1(n2056), .B2(n25568), .ZN(
        n50500) );
  OAI22_X1 U25556 ( .A1(n2076), .A2(n25584), .B1(n2055), .B2(n25567), .ZN(
        n50460) );
  OAI22_X1 U25557 ( .A1(n2075), .A2(n19206), .B1(n2054), .B2(n19196), .ZN(
        n5038) );
  OAI22_X1 U25558 ( .A1(n2074), .A2(n21267), .B1(n2053), .B2(n21230), .ZN(
        n5034) );
  OAI22_X1 U25559 ( .A1(n2073), .A2(n25584), .B1(n2052), .B2(n25567), .ZN(
        n5030) );
  OAI22_X1 U25560 ( .A1(n2072), .A2(n21258), .B1(n2051), .B2(n21221), .ZN(
        n5026) );
  OAI22_X1 U25561 ( .A1(n2071), .A2(n19209), .B1(n2050), .B2(n19199), .ZN(
        n5022) );
  OAI22_X1 U25562 ( .A1(n2070), .A2(n21264), .B1(n2049), .B2(n21228), .ZN(
        n5018) );
  OAI22_X1 U25563 ( .A1(n273500), .A2(n25524), .B1(n2705), .B2(n26517), .ZN(
        n5298) );
  OAI22_X1 U25564 ( .A1(n273400), .A2(n24639), .B1(n2704), .B2(n22465), .ZN(
        n5292) );
  OAI22_X1 U25565 ( .A1(n273300), .A2(n25669), .B1(n2703), .B2(n24655), .ZN(
        n5288) );
  OAI22_X1 U25566 ( .A1(n2732), .A2(n256701), .B1(n2702), .B2(n22453), .ZN(
        n5284) );
  OAI22_X1 U25567 ( .A1(n2731), .A2(n25668), .B1(n2701), .B2(n26525), .ZN(
        n5276) );
  OAI22_X1 U25568 ( .A1(n2730), .A2(n25672), .B1(n2700), .B2(n24661), .ZN(
        n5272) );
  OAI22_X1 U25569 ( .A1(n272900), .A2(n25525), .B1(n2699), .B2(n22450), .ZN(
        n52680) );
  OAI22_X1 U25570 ( .A1(n2728), .A2(n24638), .B1(n2698), .B2(n19267), .ZN(
        n52640) );
  OAI22_X1 U25571 ( .A1(n2727), .A2(n24633), .B1(n2697), .B2(n23450), .ZN(
        n52600) );
  OAI22_X1 U25572 ( .A1(n2726), .A2(n24635), .B1(n2696), .B2(n22462), .ZN(
        n52560) );
  OAI22_X1 U25573 ( .A1(n2725), .A2(n25666), .B1(n2695), .B2(n22948), .ZN(
        n52520) );
  OAI22_X1 U25574 ( .A1(n2724), .A2(n25673), .B1(n269400), .B2(n24664), .ZN(
        n5248) );
  OAI22_X1 U25575 ( .A1(n2723), .A2(n25667), .B1(n269300), .B2(n24667), .ZN(
        n5244) );
  OAI22_X1 U25576 ( .A1(n2722), .A2(n25671), .B1(n269200), .B2(n24665), .ZN(
        n5240) );
  OAI22_X1 U25577 ( .A1(n2721), .A2(n24636), .B1(n269100), .B2(n26519), .ZN(
        n52320) );
  AOI22_X1 U25578 ( .A1(n26511), .A2(matrix_mul_2D_0__0__0_), .B1(n25320), 
        .B2(matrix_mul_2D_0__2__0_), .ZN(n54190) );
  AOI22_X1 U25579 ( .A1(n26324), .A2(matrix_mul_2D_0__0__1_), .B1(n19301), 
        .B2(matrix_mul_2D_0__2__1_), .ZN(n50860) );
  AOI22_X1 U25580 ( .A1(n26325), .A2(matrix_mul_2D_0__0__2_), .B1(n24932), 
        .B2(matrix_mul_2D_0__2__2_), .ZN(n5040) );
  AOI22_X1 U25581 ( .A1(n22441), .A2(matrix_mul_2D_0__0__3_), .B1(n25327), 
        .B2(matrix_mul_2D_0__2__3_), .ZN(n49960) );
  AOI22_X1 U25582 ( .A1(n26324), .A2(matrix_mul_2D_0__0__4_), .B1(n24929), 
        .B2(matrix_mul_2D_0__2__4_), .ZN(n4944) );
  AOI22_X1 U25583 ( .A1(n22445), .A2(matrix_mul_2D_0__0__5_), .B1(n19081), 
        .B2(matrix_mul_2D_0__2__5_), .ZN(n4900) );
  AOI22_X1 U25584 ( .A1(n265101), .A2(matrix_mul_2D_0__0__6_), .B1(n24929), 
        .B2(matrix_mul_2D_0__2__6_), .ZN(n4849) );
  AOI22_X1 U25585 ( .A1(n26512), .A2(matrix_mul_2D_0__0__7_), .B1(n22786), 
        .B2(matrix_mul_2D_0__2__7_), .ZN(n4803) );
  AOI22_X1 U25586 ( .A1(n26325), .A2(matrix_mul_2D_0__0__8_), .B1(n25326), 
        .B2(matrix_mul_2D_0__2__8_), .ZN(n4756) );
  AOI22_X1 U25587 ( .A1(n21871), .A2(matrix_mul_2D_0__0__9_), .B1(n26711), 
        .B2(matrix_mul_2D_0__2__9_), .ZN(n47010) );
  AOI22_X1 U25588 ( .A1(n17118), .A2(matrix_mul_2D_0__0__10_), .B1(n25321), 
        .B2(matrix_mul_2D_0__2__10_), .ZN(n5372) );
  AOI22_X1 U25589 ( .A1(n22442), .A2(matrix_mul_2D_0__0__11_), .B1(n19084), 
        .B2(matrix_mul_2D_0__2__11_), .ZN(n5328) );
  AOI22_X1 U25590 ( .A1(n21870), .A2(matrix_mul_2D_0__0__12_), .B1(n24931), 
        .B2(matrix_mul_2D_0__2__12_), .ZN(n5278) );
  AOI22_X1 U25591 ( .A1(n22444), .A2(matrix_mul_2D_0__0__13_), .B1(n25321), 
        .B2(matrix_mul_2D_0__2__13_), .ZN(n5234) );
  AOI22_X1 U25592 ( .A1(n22442), .A2(matrix_mul_2D_0__0__14_), .B1(n25327), 
        .B2(matrix_mul_2D_0__2__14_), .ZN(n51860) );
  OR4_X1 U25593 ( .A1(n453), .A2(n541), .A3(n464), .A4(n538), .ZN(n4570) );
  INV_X1 U25594 ( .A(cycle_num[6]), .ZN(n27299) );
  OR2_X1 U25595 ( .A1(n27306), .A2(cycle_num[4]), .ZN(n26973) );
  INV_X1 U25596 ( .A(n24657), .ZN(n26978) );
  INV_X1 U25597 ( .A(n24656), .ZN(n26979) );
  INV_X1 U25598 ( .A(n24657), .ZN(n26980) );
  INV_X1 U25599 ( .A(n24656), .ZN(n26981) );
  INV_X1 U25600 ( .A(n24659), .ZN(n26982) );
  INV_X1 U25601 ( .A(n24659), .ZN(n26983) );
  INV_X1 U25602 ( .A(n24658), .ZN(n26984) );
  INV_X1 U25603 ( .A(n26977), .ZN(n26985) );
  INV_X1 U25604 ( .A(n26977), .ZN(n26986) );
  INV_X1 U25605 ( .A(n27001), .ZN(n27003) );
  INV_X1 U25606 ( .A(n27002), .ZN(n27004) );
  INV_X1 U25607 ( .A(n27001), .ZN(n27005) );
  INV_X1 U25608 ( .A(n24501), .ZN(n27006) );
  INV_X1 U25609 ( .A(n24502), .ZN(n27007) );
  INV_X1 U25610 ( .A(n24502), .ZN(n27008) );
  INV_X1 U25611 ( .A(n24501), .ZN(n27009) );
  INV_X1 U25612 ( .A(n24504), .ZN(n27010) );
  INV_X1 U25613 ( .A(n24504), .ZN(n27011) );
  INV_X1 U25614 ( .A(n24505), .ZN(n27012) );
  INV_X1 U25615 ( .A(n24505), .ZN(n27013) );
  INV_X1 U25616 ( .A(n24507), .ZN(n27016) );
  INV_X1 U25617 ( .A(n24506), .ZN(n27017) );
  INV_X1 U25618 ( .A(n24507), .ZN(n27018) );
  INV_X1 U25619 ( .A(n24506), .ZN(n27019) );
  INV_X1 U25620 ( .A(n24509), .ZN(n27020) );
  INV_X1 U25621 ( .A(n24510), .ZN(n27021) );
  INV_X1 U25622 ( .A(n24510), .ZN(n27022) );
  INV_X1 U25623 ( .A(n24509), .ZN(n27023) );
  INV_X1 U25624 ( .A(n27015), .ZN(n27024) );
  INV_X1 U25625 ( .A(n27014), .ZN(n27025) );
  INV_X1 U25626 ( .A(n27015), .ZN(n27026) );
  INV_X1 U25627 ( .A(n24597), .ZN(n27032) );
  INV_X1 U25628 ( .A(n24596), .ZN(n27033) );
  INV_X1 U25629 ( .A(n24597), .ZN(n27034) );
  INV_X1 U25630 ( .A(n24596), .ZN(n27035) );
  INV_X1 U25631 ( .A(n27030), .ZN(n27036) );
  INV_X1 U25632 ( .A(n27031), .ZN(n27037) );
  INV_X1 U25633 ( .A(n27030), .ZN(n27038) );
  INV_X1 U25634 ( .A(n24600), .ZN(n27039) );
  INV_X1 U25635 ( .A(n24599), .ZN(n27040) );
  INV_X1 U25636 ( .A(n24599), .ZN(n27041) );
  INV_X1 U25637 ( .A(n24600), .ZN(n27042) );
  INV_X1 U25638 ( .A(n27048), .ZN(n27050) );
  INV_X1 U25639 ( .A(n27049), .ZN(n27051) );
  INV_X1 U25640 ( .A(n27048), .ZN(n27052) );
  INV_X1 U25641 ( .A(n24591), .ZN(n27053) );
  INV_X1 U25642 ( .A(n24592), .ZN(n27054) );
  INV_X1 U25643 ( .A(n24592), .ZN(n27055) );
  INV_X1 U25644 ( .A(n24591), .ZN(n27056) );
  INV_X1 U25645 ( .A(n24594), .ZN(n27057) );
  INV_X1 U25646 ( .A(n24594), .ZN(n27058) );
  INV_X1 U25647 ( .A(n24595), .ZN(n27059) );
  INV_X1 U25648 ( .A(n24595), .ZN(n27060) );
  INV_X1 U25649 ( .A(n24586), .ZN(n27063) );
  INV_X1 U25650 ( .A(n24585), .ZN(n27064) );
  INV_X1 U25651 ( .A(n24586), .ZN(n27065) );
  INV_X1 U25652 ( .A(n24585), .ZN(n27066) );
  INV_X1 U25653 ( .A(n24589), .ZN(n27067) );
  INV_X1 U25654 ( .A(n24590), .ZN(n27068) );
  INV_X1 U25655 ( .A(n24590), .ZN(n27069) );
  INV_X1 U25656 ( .A(n24589), .ZN(n27070) );
  INV_X1 U25657 ( .A(n27062), .ZN(n27071) );
  INV_X1 U25658 ( .A(n27062), .ZN(n27072) );
  INV_X1 U25659 ( .A(n27073), .ZN(n27076) );
  INV_X1 U25660 ( .A(n26966), .ZN(n27077) );
  INV_X1 U25661 ( .A(n22942), .ZN(n27078) );
  INV_X1 U25662 ( .A(n27075), .ZN(n27079) );
  INV_X1 U25663 ( .A(n27074), .ZN(n27080) );
  INV_X1 U25664 ( .A(n27075), .ZN(n27081) );
  INV_X1 U25665 ( .A(n22942), .ZN(n27082) );
  INV_X1 U25666 ( .A(n27074), .ZN(n27083) );
  INV_X1 U25667 ( .A(n26966), .ZN(n27084) );
  INV_X1 U25668 ( .A(n24497), .ZN(n27087) );
  INV_X1 U25669 ( .A(n24496), .ZN(n27088) );
  INV_X1 U25670 ( .A(n24497), .ZN(n27089) );
  INV_X1 U25671 ( .A(n24496), .ZN(n27090) );
  INV_X1 U25672 ( .A(n27085), .ZN(n27091) );
  INV_X1 U25673 ( .A(n27086), .ZN(n27092) );
  INV_X1 U25674 ( .A(n27085), .ZN(n27093) );
  INV_X1 U25675 ( .A(n24499), .ZN(n27094) );
  INV_X1 U25676 ( .A(n24499), .ZN(n27095) );
  INV_X1 U25677 ( .A(n24500), .ZN(n27096) );
  INV_X1 U25678 ( .A(n24500), .ZN(n27097) );
  INV_X1 U25679 ( .A(n24584), .ZN(n27100) );
  INV_X1 U25680 ( .A(n24583), .ZN(n27101) );
  INV_X1 U25681 ( .A(n24584), .ZN(n27102) );
  INV_X1 U25682 ( .A(n24583), .ZN(n27103) );
  INV_X1 U25683 ( .A(n24587), .ZN(n27104) );
  INV_X1 U25684 ( .A(n24588), .ZN(n27105) );
  INV_X1 U25685 ( .A(n24588), .ZN(n27106) );
  INV_X1 U25686 ( .A(n24587), .ZN(n27107) );
  INV_X1 U25687 ( .A(n27099), .ZN(n27108) );
  INV_X1 U25688 ( .A(n27099), .ZN(n27109) );
  INV_X1 U25689 ( .A(n25089), .ZN(n27128) );
  INV_X1 U25690 ( .A(n25089), .ZN(n27129) );
  INV_X1 U25691 ( .A(n20898), .ZN(n27130) );
  INV_X1 U25692 ( .A(n19319), .ZN(n27131) );
  INV_X1 U25693 ( .A(n27130), .ZN(n27132) );
  INV_X1 U25694 ( .A(n27128), .ZN(n27133) );
  INV_X1 U25695 ( .A(n27129), .ZN(n27134) );
  INV_X1 U25696 ( .A(n27128), .ZN(n27135) );
  INV_X1 U25697 ( .A(n22968), .ZN(n27136) );
  INV_X1 U25698 ( .A(n22969), .ZN(n27137) );
  INV_X1 U25699 ( .A(n19319), .ZN(n27138) );
  INV_X1 U25700 ( .A(n27130), .ZN(n27139) );
  INV_X1 U25701 ( .A(n24670), .ZN(n27140) );
  INV_X1 U25702 ( .A(n22968), .ZN(n27141) );
  INV_X1 U25703 ( .A(n24671), .ZN(n27142) );
  INV_X1 U25704 ( .A(n24670), .ZN(n27143) );
  INV_X1 U25705 ( .A(n24671), .ZN(n27144) );
  INV_X1 U25706 ( .A(n25086), .ZN(n27276) );
  INV_X1 U25707 ( .A(n25086), .ZN(n27277) );
  INV_X1 U25708 ( .A(n20894), .ZN(n27278) );
  INV_X1 U25709 ( .A(n19322), .ZN(n27279) );
  INV_X1 U25710 ( .A(n27278), .ZN(n27280) );
  INV_X1 U25711 ( .A(n27276), .ZN(n27281) );
  INV_X1 U25712 ( .A(n27277), .ZN(n27282) );
  INV_X1 U25713 ( .A(n27276), .ZN(n27283) );
  INV_X1 U25714 ( .A(n22971), .ZN(n27284) );
  INV_X1 U25715 ( .A(n22972), .ZN(n27285) );
  INV_X1 U25716 ( .A(n19322), .ZN(n27286) );
  INV_X1 U25717 ( .A(n27278), .ZN(n27287) );
  INV_X1 U25718 ( .A(n24673), .ZN(n27288) );
  INV_X1 U25719 ( .A(n22971), .ZN(n27289) );
  INV_X1 U25720 ( .A(n24674), .ZN(n272901) );
  INV_X1 U25721 ( .A(n24673), .ZN(n27291) );
  INV_X1 U25722 ( .A(n24674), .ZN(n27292) );
  NOR2_X1 U25723 ( .A1(cycle_num[1]), .A2(n875), .ZN(n27293) );
  NOR2_X1 U25724 ( .A1(n27304), .A2(n466), .ZN(n27294) );
  NOR2_X1 U25725 ( .A1(n27305), .A2(n551), .ZN(n27295) );
  NOR2_X1 U25726 ( .A1(n26973), .A2(n540), .ZN(n27297) );
  AOI21_X1 U25727 ( .B1(n17998), .B2(n459), .A(n17999), .ZN(n27296) );
  OAI21_X1 U25728 ( .B1(n460), .B2(n24680), .A(n465), .ZN(n27298) );
  NAND3_X1 U25729 ( .A1(n23742), .A2(n26509), .A3(n23953), .ZN(n27308) );
  NOR4_X1 U25730 ( .A1(n18823), .A2(n17071), .A3(n26604), .A4(n23944), .ZN(
        n27307) );
  NAND3_X1 U25731 ( .A1(n27311), .A2(n27308), .A3(n27307), .ZN(N7942) );
  NOR2_X1 U25732 ( .A1(n23738), .A2(n23958), .ZN(n27311) );
  OAI211_X1 U25733 ( .C1(n17122), .C2(n22436), .A(n22545), .B(n23950), .ZN(
        n27310) );
  NOR4_X1 U25734 ( .A1(n18823), .A2(n17070), .A3(n23941), .A4(n23946), .ZN(
        n27309) );
  NAND3_X1 U25735 ( .A1(n27311), .A2(n27310), .A3(n27309), .ZN(N7267) );
  AOI211_X1 U25736 ( .C1(n23952), .C2(n22544), .A(n26593), .B(n23959), .ZN(
        n27313) );
  NOR4_X1 U25737 ( .A1(n24015), .A2(n17070), .A3(n26604), .A4(r899_B_6_), .ZN(
        n27312) );
  NAND2_X1 U25738 ( .A1(n27313), .A2(n27312), .ZN(N6563) );
  AOI21_X1 U25739 ( .B1(n22437), .B2(n19176), .A(n22542), .ZN(n27315) );
  NOR2_X1 U25740 ( .A1(n26594), .A2(n26613), .ZN(n27314) );
  OAI211_X1 U25741 ( .C1(n27315), .C2(n18818), .A(n27314), .B(n27327), .ZN(
        N5888) );
  NOR2_X1 U25742 ( .A1(n26594), .A2(n26612), .ZN(n27317) );
  OAI21_X1 U25743 ( .B1(n26509), .B2(n22545), .A(n23953), .ZN(n27316) );
  NAND3_X1 U25744 ( .A1(n27317), .A2(n27316), .A3(n27323), .ZN(N5213) );
  OR3_X1 U25745 ( .A1(n22541), .A2(n22436), .A3(n25513), .ZN(n27318) );
  AOI211_X1 U25746 ( .C1(n26608), .C2(n27318), .A(n23735), .B(n23955), .ZN(
        n27319) );
  NAND2_X1 U25747 ( .A1(n27319), .A2(n27309), .ZN(N4509) );
  OR4_X1 U25748 ( .A1(n23940), .A2(n23943), .A3(n17105), .A4(n23936), .ZN(
        n27320) );
  OR4_X1 U25749 ( .A1(n26595), .A2(n23956), .A3(n26609), .A4(n27320), .ZN(
        r948_LT_LE) );
  AND3_X1 U25750 ( .A1(n26507), .A2(n19176), .A3(n23741), .ZN(n27321) );
  NOR4_X1 U25751 ( .A1(n23739), .A2(r899_B_4_), .A3(n23950), .A4(n27321), .ZN(
        n27322) );
  NAND2_X1 U25752 ( .A1(n27322), .A2(n27307), .ZN(r929_LT_LE) );
  AOI21_X1 U25753 ( .B1(n22544), .B2(n22440), .A(n26607), .ZN(n27325) );
  NOR2_X1 U25754 ( .A1(n23735), .A2(n23955), .ZN(n27324) );
  NOR4_X1 U25755 ( .A1(n17068), .A2(n17072), .A3(n17069), .A4(n23944), .ZN(
        n27323) );
  NAND3_X1 U25756 ( .A1(n27325), .A2(n27324), .A3(n27323), .ZN(r924_LT_LE) );
  OAI21_X1 U25757 ( .B1(n25514), .B2(n22439), .A(n19271), .ZN(n27326) );
  NAND4_X1 U25758 ( .A1(n27326), .A2(n18818), .A3(n27314), .A4(n27312), .ZN(
        N2985) );
  NOR4_X1 U25759 ( .A1(n23736), .A2(n26611), .A3(n26606), .A4(n22542), .ZN(
        n27328) );
  NOR4_X1 U25760 ( .A1(n17105), .A2(n23936), .A3(n23940), .A4(n26605), .ZN(
        n27327) );
  NAND2_X1 U25761 ( .A1(n27328), .A2(n27327), .ZN(N2903) );
  AOI21_X1 U25762 ( .B1(n26508), .B2(n17122), .A(n23742), .ZN(n273301) );
  NOR2_X1 U25763 ( .A1(n23958), .A2(n23952), .ZN(n27329) );
  NAND4_X1 U25764 ( .A1(n273301), .A2(n27329), .A3(n27334), .A4(n27333), .ZN(
        N2811) );
  NOR2_X1 U25765 ( .A1(n23943), .A2(n23738), .ZN(n27332) );
  NOR4_X1 U25766 ( .A1(n26613), .A2(n26608), .A3(n22541), .A4(n26508), .ZN(
        n27331) );
  NAND3_X1 U25767 ( .A1(n27332), .A2(n17130), .A3(n27331), .ZN(N2729) );
  NOR2_X1 U25768 ( .A1(n22439), .A2(n25514), .ZN(n27336) );
  NOR3_X1 U25769 ( .A1(n23741), .A2(n23956), .A3(n26609), .ZN(n27335) );
  NOR2_X1 U25770 ( .A1(n23946), .A2(n23736), .ZN(n27334) );
  NOR3_X1 U25771 ( .A1(n23941), .A2(n24015), .A3(n23937), .ZN(n27333) );
  NAND4_X1 U25772 ( .A1(n27336), .A2(n27335), .A3(n27334), .A4(n17130), .ZN(
        N2637) );
  OR4_X1 U25773 ( .A1(n543), .A2(n452), .A3(n552), .A4(n466), .ZN(n27337) );
  AOI21_X1 U25774 ( .B1(n542), .B2(n27337), .A(n541), .ZN(n27339) );
  NOR3_X1 U25775 ( .A1(n453), .A2(n464), .A3(n460), .ZN(n27338) );
  OR3_X1 U25776 ( .A1(n467), .A2(n455), .A3(n876), .ZN(n273401) );
  AOI211_X1 U25777 ( .C1(n551), .C2(n273401), .A(n459), .B(n454), .ZN(n27341)
         );
endmodule


module systolic_controll_ARRAY_SIZE8_DW01_inc_1 ( A, SUM );
  input [8:0] A;
  output [8:0] SUM;

  wire   [8:2] carry;

  HA_X1 U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  HA_X1 U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2_X1 U1 ( .A(carry[8]), .B(A[8]), .Z(SUM[8]) );
  INV_X1 U2 ( .A(A[0]), .ZN(SUM[0]) );
endmodule


module systolic_controll_ARRAY_SIZE8_DW01_inc_2 ( A, SUM_6_, SUM_5_, SUM_4_, 
        SUM_3_, SUM_2_, SUM_1_ );
  input [6:0] A;
  output SUM_6_, SUM_5_, SUM_4_, SUM_3_, SUM_2_, SUM_1_;

  wire   [6:2] carry;

  HA_X1 U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM_5_) );
  HA_X1 U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM_4_) );
  HA_X1 U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM_3_) );
  HA_X1 U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM_2_) );
  HA_X1 U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM_1_) );
  XOR2_X1 U1 ( .A(carry[6]), .B(A[6]), .Z(SUM_6_) );
endmodule


module systolic_controll_ARRAY_SIZE8 ( clk, srstn, tpu_start, 
        sram_write_enable, addr_serial_num, alu_start, cycle_num, matrix_index, 
        data_set, tpu_done );
  output [6:0] addr_serial_num;
  output [8:0] cycle_num;
  output [5:0] matrix_index;
  output [1:0] data_set;
  input clk, srstn, tpu_start;
  output sram_write_enable, alu_start, tpu_done;
  wire   n235, n236, n237, n238, n239, n240, n241, n242, n243, n244, n245,
         n246, n247, n248, n249, n250, n251, n252, n253, n254, n255, n256,
         n257, n258, N25, N26, N27, N37, N38, N39, N40, N41, N42, N43, N44,
         N50, N83, N84, N85, N86, N87, N88, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N125, N126, N127, N128, N129, N130, n22, n23,
         n270, n29, n30, n34, n35, n36, n370, n380, n390, n400, n410, n440,
         n45, n46, n47, n48, n49, n500, n51, n52, n53, n54, n56, n57, n58, n1,
         n4, n5, n6, n7, n8, n9, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n24, n259, n260, n28, n31, n32, n33, n420, n430, n55, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n78, n79, n80, n81, n82, n830, n840, n850, n860, n870, n89, n90,
         n91, n92, n93, n94, n95, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n1110, n1120, n1130, n1140, n1150,
         n1160, n1170, n1180, n1190, n121, n123, n1250, n1260, n1270, n1280,
         n1290, n1300, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n146, n147, n148, n150, n152, n153,
         n155, n157, n158, n159, n160, n162, n163, n164, n165, n167, n168,
         n169, n170, n171, n172, n173, n175, n176, n177, n178, n179, n180,
         n181, n182, n184, n185, n186, n187, n188, n190, n192, n193, n194,
         n195, n196, n198, n199, n200, n201, n202, n203, n204, n206, n207,
         n208, n209, n210, n212, n213, n214, n215, n216, n217, n218, n219,
         n220, n221, n222, n223, n224, n225, n226, n227, n228, n229, n230,
         n231, n232, n233, n234;
  wire   [1:0] state;
  wire   [5:2] add_166_carry;

  DFF_X1 matrix_index_reg_1_ ( .D(N38), .CK(clk), .Q(n255), .QN(n188) );
  DFF_X1 matrix_index_reg_2_ ( .D(N39), .CK(clk), .Q(n254), .QN(n155) );
  DFF_X1 matrix_index_reg_3_ ( .D(N40), .CK(clk), .Q(n253), .QN(n210) );
  DFF_X1 matrix_index_reg_4_ ( .D(N41), .CK(clk), .Q(n252), .QN(n204) );
  DFF_X1 matrix_index_reg_5_ ( .D(n9), .CK(clk), .Q(n251), .QN(n173) );
  DFF_X1 data_set_reg_1_ ( .D(N27), .CK(clk), .Q(n257), .QN(n78) );
  DFF_X1 tpu_done_reg ( .D(N50), .CK(clk), .Q(tpu_done) );
  DFF_X1 addr_serial_num_reg_2_ ( .D(n232), .CK(clk), .Q(n239), .QN(n89) );
  DFF_X1 addr_serial_num_reg_3_ ( .D(n231), .CK(clk), .Q(n238), .QN(n93) );
  DFF_X1 addr_serial_num_reg_4_ ( .D(n230), .CK(clk), .Q(n237), .QN(n91) );
  DFF_X1 addr_serial_num_reg_5_ ( .D(n229), .CK(clk), .Q(n236), .QN(n175) );
  DFF_X1 addr_serial_num_reg_6_ ( .D(n8), .CK(clk), .Q(n235), .QN(n146) );
  OAI33_X1 U67 ( .A1(n134), .A2(n227), .A3(n101), .B1(n104), .B2(n97), .B3(n99), .ZN(N26) );
  systolic_controll_ARRAY_SIZE8_DW01_inc_1 add_159 ( .A({n177, n185, n158, 
        n181, n195, n201, n163, n179, n98}), .SUM({N119, N118, N117, N116, 
        N115, N114, N113, N112, N111}) );
  systolic_controll_ARRAY_SIZE8_DW01_inc_2 add_121 ( .A({n235, n199, n1120, 
        n170, n165, n240, n160}), .SUM_6_(N88), .SUM_5_(N87), .SUM_4_(N86), 
        .SUM_3_(N85), .SUM_2_(N84), .SUM_1_(N83) );
  HA_X1 add_166_U1_1_1 ( .A(n203), .B(n198), .CO(add_166_carry[2]), .S(N126)
         );
  HA_X1 add_166_U1_1_2 ( .A(n187), .B(add_166_carry[2]), .CO(add_166_carry[3]), 
        .S(N127) );
  HA_X1 add_166_U1_1_3 ( .A(n213), .B(add_166_carry[3]), .CO(add_166_carry[4]), 
        .S(N128) );
  HA_X1 add_166_U1_1_4 ( .A(n208), .B(add_166_carry[4]), .CO(add_166_carry[5]), 
        .S(N129) );
  DFF_X1 state_reg_0_ ( .D(n69), .CK(clk), .Q(state[0]), .QN(n29) );
  DFF_X1 cycle_num_reg_8_ ( .D(n20), .CK(clk), .Q(n242), .QN(n121) );
  DFF_X1 cycle_num_reg_7_ ( .D(n221), .CK(clk), .Q(n243), .QN(n153) );
  DFF_X1 cycle_num_reg_6_ ( .D(n220), .CK(clk), .Q(n244), .QN(n870) );
  DFF_X1 cycle_num_reg_5_ ( .D(n219), .CK(clk), .Q(n245), .QN(n148) );
  DFF_X1 cycle_num_reg_4_ ( .D(n218), .CK(clk), .Q(n246), .QN(n144) );
  DFF_X1 cycle_num_reg_3_ ( .D(n217), .CK(clk), .Q(n247), .QN(n182) );
  DFF_X1 cycle_num_reg_2_ ( .D(n216), .CK(clk), .Q(n248), .QN(n1190) );
  DFF_X1 cycle_num_reg_1_ ( .D(n215), .CK(clk), .Q(n249), .QN(n150) );
  DFF_X1 cycle_num_reg_0_ ( .D(n1), .CK(clk), .Q(n250), .QN(n190) );
  DFF_X1 state_reg_1_ ( .D(n66), .CK(clk), .Q(state[1]), .QN(n270) );
  DFF_X1 data_set_reg_0_ ( .D(n33), .CK(clk), .Q(n258), .QN(n30) );
  DFF_X1 addr_serial_num_reg_0_ ( .D(n420), .CK(clk), .Q(n241), .QN(n23) );
  DFF_X1 matrix_index_reg_0_ ( .D(n61), .CK(clk), .Q(n256), .QN(N125) );
  DFF_X1 addr_serial_num_reg_1_ ( .D(n21), .CK(clk), .Q(n240), .QN(n22) );
  INV_X2 U3 ( .A(n89), .ZN(n90) );
  BUF_X1 U4 ( .A(n214), .Z(n1) );
  INV_X2 U5 ( .A(n241), .ZN(n159) );
  INV_X1 U6 ( .A(n91), .ZN(n92) );
  INV_X1 U7 ( .A(n93), .ZN(n94) );
  INV_X1 U8 ( .A(n15), .ZN(addr_serial_num[5]) );
  INV_X1 U9 ( .A(n16), .ZN(addr_serial_num[6]) );
  AND2_X1 U10 ( .A1(n139), .A2(n29), .ZN(n4) );
  AND4_X1 U11 ( .A1(n187), .A2(n203), .A3(n213), .A4(n58), .ZN(n5) );
  BUF_X1 U12 ( .A(srstn), .Z(n6) );
  INV_X1 U13 ( .A(n860), .ZN(n7) );
  BUF_X1 U14 ( .A(n228), .Z(n8) );
  INV_X2 U15 ( .A(n78), .ZN(n79) );
  OAI21_X2 U16 ( .B1(n137), .B2(n104), .A(n53), .ZN(N27) );
  INV_X2 U17 ( .A(n257), .ZN(n123) );
  BUF_X1 U18 ( .A(N42), .Z(n9) );
  AND2_X2 U19 ( .A1(N129), .A2(n172), .ZN(N41) );
  AND2_X2 U20 ( .A1(N128), .A2(n171), .ZN(N40) );
  AND2_X2 U21 ( .A1(N127), .A2(n171), .ZN(N39) );
  AND2_X2 U22 ( .A1(N126), .A2(n82), .ZN(N38) );
  AND2_X2 U23 ( .A1(N115), .A2(n131), .ZN(n218) );
  AND2_X2 U24 ( .A1(N114), .A2(n1280), .ZN(n217) );
  BUF_X1 U25 ( .A(n90), .Z(addr_serial_num[2]) );
  BUF_X1 U26 ( .A(n94), .Z(addr_serial_num[3]) );
  BUF_X1 U27 ( .A(n92), .Z(addr_serial_num[4]) );
  CLKBUF_X1 U28 ( .A(n175), .Z(n13) );
  INV_X1 U29 ( .A(n13), .ZN(n14) );
  INV_X1 U30 ( .A(n14), .ZN(n15) );
  INV_X1 U31 ( .A(n19), .ZN(n16) );
  INV_X1 U32 ( .A(n16), .ZN(n17) );
  INV_X1 U33 ( .A(n147), .ZN(n18) );
  INV_X1 U34 ( .A(n18), .ZN(n19) );
  BUF_X1 U35 ( .A(n222), .Z(n20) );
  BUF_X1 U36 ( .A(n28), .Z(n21) );
  INV_X1 U37 ( .A(n22), .ZN(n24) );
  INV_X1 U38 ( .A(n24), .ZN(n259) );
  INV_X1 U39 ( .A(N44), .ZN(n260) );
  INV_X1 U40 ( .A(n260), .ZN(n28) );
  INV_X2 U41 ( .A(N26), .ZN(n32) );
  BUF_X1 U42 ( .A(n100), .Z(n31) );
  INV_X1 U43 ( .A(n32), .ZN(n33) );
  BUF_X1 U44 ( .A(n55), .Z(n420) );
  INV_X1 U45 ( .A(n60), .ZN(n430) );
  INV_X1 U46 ( .A(n430), .ZN(n55) );
  INV_X1 U47 ( .A(N43), .ZN(n59) );
  INV_X1 U48 ( .A(n59), .ZN(n60) );
  BUF_X1 U49 ( .A(n63), .Z(n61) );
  INV_X1 U50 ( .A(n65), .ZN(n62) );
  INV_X1 U51 ( .A(n62), .ZN(n63) );
  INV_X1 U52 ( .A(N37), .ZN(n64) );
  INV_X1 U53 ( .A(n64), .ZN(n65) );
  BUF_X1 U54 ( .A(n68), .Z(n66) );
  INV_X1 U55 ( .A(N25), .ZN(n67) );
  INV_X1 U56 ( .A(n67), .ZN(n68) );
  AND2_X2 U57 ( .A1(N113), .A2(n830), .ZN(n216) );
  AND2_X2 U58 ( .A1(N112), .A2(n1260), .ZN(n215) );
  AND2_X2 U59 ( .A1(N118), .A2(n1290), .ZN(n221) );
  BUF_X1 U60 ( .A(n71), .Z(n69) );
  INV_X1 U61 ( .A(n223), .ZN(n70) );
  INV_X1 U62 ( .A(n70), .ZN(n71) );
  AND2_X2 U63 ( .A1(N116), .A2(n1170), .ZN(n219) );
  AND2_X2 U64 ( .A1(N117), .A2(n209), .ZN(n220) );
  CLKBUF_X1 U65 ( .A(n6), .Z(n72) );
  CLKBUF_X1 U66 ( .A(n410), .Z(n73) );
  CLKBUF_X1 U68 ( .A(n81), .Z(n74) );
  CLKBUF_X1 U69 ( .A(n233), .Z(n75) );
  CLKBUF_X1 U70 ( .A(n1160), .Z(n76) );
  CLKBUF_X1 U71 ( .A(n234), .Z(alu_start) );
  CLKBUF_X1 U72 ( .A(n34), .Z(n80) );
  CLKBUF_X1 U73 ( .A(n410), .Z(n81) );
  CLKBUF_X1 U74 ( .A(n51), .Z(n82) );
  CLKBUF_X1 U75 ( .A(n75), .Z(n830) );
  CLKBUF_X1 U76 ( .A(n5), .Z(n840) );
  INV_X1 U77 ( .A(n72), .ZN(n850) );
  INV_X1 U78 ( .A(n72), .ZN(n860) );
  INV_X1 U79 ( .A(n870), .ZN(cycle_num[6]) );
  INV_X1 U80 ( .A(n258), .ZN(n95) );
  INV_X1 U81 ( .A(n95), .ZN(data_set[0]) );
  INV_X1 U82 ( .A(n95), .ZN(n97) );
  INV_X1 U83 ( .A(n206), .ZN(n98) );
  INV_X1 U84 ( .A(n5), .ZN(n99) );
  INV_X1 U85 ( .A(n30), .ZN(n100) );
  INV_X1 U86 ( .A(n31), .ZN(n101) );
  INV_X1 U87 ( .A(n31), .ZN(n102) );
  INV_X1 U88 ( .A(n52), .ZN(n103) );
  INV_X1 U89 ( .A(n103), .ZN(n104) );
  INV_X1 U90 ( .A(n4), .ZN(n105) );
  INV_X1 U91 ( .A(n74), .ZN(n106) );
  INV_X1 U92 ( .A(n74), .ZN(n107) );
  INV_X1 U93 ( .A(n164), .ZN(n108) );
  INV_X1 U94 ( .A(n108), .ZN(n109) );
  INV_X1 U95 ( .A(n168), .ZN(n110) );
  INV_X1 U96 ( .A(n110), .ZN(n1110) );
  INV_X1 U97 ( .A(n110), .ZN(n1120) );
  INV_X1 U98 ( .A(n170), .ZN(n1130) );
  INV_X1 U99 ( .A(n1130), .ZN(n1140) );
  INV_X1 U100 ( .A(n51), .ZN(n1150) );
  INV_X1 U101 ( .A(n75), .ZN(n1160) );
  INV_X1 U102 ( .A(n76), .ZN(n1170) );
  INV_X1 U103 ( .A(n76), .ZN(n1180) );
  INV_X1 U104 ( .A(n1190), .ZN(cycle_num[2]) );
  INV_X1 U105 ( .A(n121), .ZN(cycle_num[8]) );
  INV_X1 U106 ( .A(n123), .ZN(data_set[1]) );
  INV_X1 U107 ( .A(n123), .ZN(n1250) );
  CLKBUF_X1 U108 ( .A(n233), .Z(n1260) );
  INV_X1 U109 ( .A(n1170), .ZN(n1270) );
  INV_X1 U110 ( .A(n1270), .ZN(n1280) );
  INV_X1 U111 ( .A(n1270), .ZN(n1290) );
  INV_X1 U112 ( .A(n80), .ZN(n1300) );
  INV_X1 U113 ( .A(n80), .ZN(n131) );
  INV_X1 U114 ( .A(n34), .ZN(n132) );
  INV_X1 U115 ( .A(n132), .ZN(n133) );
  INV_X1 U116 ( .A(n132), .ZN(n134) );
  INV_X1 U117 ( .A(n35), .ZN(n135) );
  INV_X1 U118 ( .A(n135), .ZN(n136) );
  INV_X1 U119 ( .A(n135), .ZN(n137) );
  INV_X1 U120 ( .A(state[1]), .ZN(n138) );
  INV_X1 U121 ( .A(n138), .ZN(n139) );
  INV_X1 U122 ( .A(n138), .ZN(n140) );
  INV_X1 U123 ( .A(state[0]), .ZN(n141) );
  INV_X1 U124 ( .A(n141), .ZN(n142) );
  INV_X1 U125 ( .A(n141), .ZN(n143) );
  INV_X1 U126 ( .A(n144), .ZN(cycle_num[4]) );
  INV_X1 U127 ( .A(n146), .ZN(n147) );
  INV_X1 U128 ( .A(n148), .ZN(cycle_num[5]) );
  INV_X1 U129 ( .A(n150), .ZN(cycle_num[1]) );
  INV_X1 U130 ( .A(n81), .ZN(n152) );
  INV_X1 U131 ( .A(n153), .ZN(cycle_num[7]) );
  INV_X1 U132 ( .A(n155), .ZN(matrix_index[2]) );
  INV_X1 U133 ( .A(n244), .ZN(n157) );
  INV_X1 U134 ( .A(n157), .ZN(n158) );
  INV_X1 U135 ( .A(n159), .ZN(n160) );
  INV_X1 U136 ( .A(n159), .ZN(addr_serial_num[0]) );
  INV_X1 U137 ( .A(n248), .ZN(n162) );
  INV_X1 U138 ( .A(n162), .ZN(n163) );
  INV_X1 U139 ( .A(n239), .ZN(n164) );
  INV_X1 U140 ( .A(n109), .ZN(n165) );
  INV_X1 U141 ( .A(n259), .ZN(addr_serial_num[1]) );
  INV_X1 U142 ( .A(n237), .ZN(n167) );
  INV_X1 U143 ( .A(n167), .ZN(n168) );
  INV_X1 U144 ( .A(n238), .ZN(n169) );
  INV_X1 U145 ( .A(n169), .ZN(n170) );
  INV_X1 U146 ( .A(n1150), .ZN(n171) );
  INV_X1 U147 ( .A(n1150), .ZN(n172) );
  INV_X1 U148 ( .A(n173), .ZN(matrix_index[5]) );
  INV_X1 U149 ( .A(n242), .ZN(n176) );
  INV_X1 U150 ( .A(n176), .ZN(n177) );
  INV_X1 U151 ( .A(n249), .ZN(n178) );
  INV_X1 U152 ( .A(n178), .ZN(n179) );
  INV_X1 U153 ( .A(n245), .ZN(n180) );
  INV_X1 U154 ( .A(n180), .ZN(n181) );
  INV_X1 U155 ( .A(n182), .ZN(cycle_num[3]) );
  INV_X1 U156 ( .A(n243), .ZN(n184) );
  INV_X1 U157 ( .A(n184), .ZN(n185) );
  INV_X1 U158 ( .A(n254), .ZN(n186) );
  INV_X1 U159 ( .A(n186), .ZN(n187) );
  INV_X1 U160 ( .A(n188), .ZN(matrix_index[1]) );
  INV_X1 U161 ( .A(n190), .ZN(cycle_num[0]) );
  INV_X1 U162 ( .A(n251), .ZN(n192) );
  INV_X1 U163 ( .A(n192), .ZN(n193) );
  INV_X1 U164 ( .A(n246), .ZN(n194) );
  INV_X1 U165 ( .A(n194), .ZN(n195) );
  INV_X1 U166 ( .A(n256), .ZN(n196) );
  INV_X1 U167 ( .A(n196), .ZN(matrix_index[0]) );
  INV_X1 U168 ( .A(n196), .ZN(n198) );
  INV_X1 U169 ( .A(n15), .ZN(n199) );
  INV_X1 U170 ( .A(n247), .ZN(n200) );
  INV_X1 U171 ( .A(n200), .ZN(n201) );
  INV_X1 U172 ( .A(n255), .ZN(n202) );
  INV_X1 U173 ( .A(n202), .ZN(n203) );
  INV_X1 U174 ( .A(n204), .ZN(matrix_index[4]) );
  INV_X1 U175 ( .A(n250), .ZN(n206) );
  INV_X1 U176 ( .A(n252), .ZN(n207) );
  INV_X1 U177 ( .A(n207), .ZN(n208) );
  INV_X1 U178 ( .A(n1160), .ZN(n209) );
  INV_X1 U179 ( .A(n210), .ZN(matrix_index[3]) );
  INV_X1 U180 ( .A(n253), .ZN(n212) );
  INV_X1 U181 ( .A(n212), .ZN(n213) );
  AND2_X1 U182 ( .A1(N111), .A2(n131), .ZN(n214) );
  AND2_X1 U183 ( .A1(N119), .A2(n1300), .ZN(n222) );
  NOR2_X1 U184 ( .A1(n57), .A2(n850), .ZN(n223) );
  INV_X1 U185 ( .A(n500), .ZN(n234) );
  INV_X1 U186 ( .A(n133), .ZN(n233) );
  NOR2_X1 U187 ( .A1(n52), .A2(n840), .ZN(n51) );
  NOR2_X1 U188 ( .A1(n134), .A2(n136), .ZN(N50) );
  AND2_X1 U189 ( .A1(N120), .A2(alu_start), .ZN(sram_write_enable) );
  NAND2_X1 U190 ( .A1(n840), .A2(N120), .ZN(n54) );
  INV_X1 U191 ( .A(n54), .ZN(n227) );
  OAI21_X1 U192 ( .B1(n46), .B2(n47), .A(n7), .ZN(n410) );
  NOR4_X1 U193 ( .A1(n48), .A2(n49), .A3(n500), .A4(n23), .ZN(n47) );
  NOR3_X1 U194 ( .A1(n143), .A2(tpu_start), .A3(n140), .ZN(n46) );
  NAND2_X1 U195 ( .A1(n90), .A2(n24), .ZN(n49) );
  AOI221_X1 U196 ( .B1(tpu_start), .B2(n29), .C1(n140), .C2(n136), .A(n4), 
        .ZN(n57) );
  OAI221_X1 U197 ( .B1(n23), .B2(n73), .C1(n133), .C2(n160), .A(n45), .ZN(N43)
         );
  NAND3_X1 U198 ( .A1(n143), .A2(n270), .A3(n7), .ZN(n45) );
  OAI221_X1 U199 ( .B1(n259), .B2(n73), .C1(n860), .C2(n105), .A(n440), .ZN(
        N44) );
  NAND2_X1 U200 ( .A1(N83), .A2(n209), .ZN(n440) );
  INV_X1 U201 ( .A(n370), .ZN(n229) );
  AOI22_X1 U202 ( .A1(n1290), .A2(N87), .B1(n199), .B2(n106), .ZN(n370) );
  INV_X1 U203 ( .A(n36), .ZN(n228) );
  AOI22_X1 U204 ( .A1(n1300), .A2(N88), .B1(n17), .B2(n152), .ZN(n36) );
  INV_X1 U205 ( .A(n380), .ZN(n230) );
  AOI22_X1 U206 ( .A1(n1180), .A2(N86), .B1(n1110), .B2(n107), .ZN(n380) );
  INV_X1 U207 ( .A(n390), .ZN(n231) );
  AOI22_X1 U208 ( .A1(n1260), .A2(N85), .B1(n1140), .B2(n152), .ZN(n390) );
  INV_X1 U209 ( .A(n400), .ZN(n232) );
  AOI22_X1 U210 ( .A1(n1280), .A2(N84), .B1(n165), .B2(n106), .ZN(n400) );
  NAND2_X1 U211 ( .A1(n139), .A2(n142), .ZN(n500) );
  NAND2_X1 U212 ( .A1(srstn), .A2(n234), .ZN(n34) );
  NAND2_X1 U213 ( .A1(sram_write_enable), .A2(n6), .ZN(n52) );
  AOI21_X1 U214 ( .B1(n105), .B2(n56), .A(n850), .ZN(N25) );
  OAI21_X1 U215 ( .B1(n270), .B2(n137), .A(n142), .ZN(n56) );
  OAI211_X1 U216 ( .C1(n102), .C2(n54), .A(n830), .B(n1250), .ZN(n53) );
  AND2_X1 U217 ( .A1(N130), .A2(n82), .ZN(N42) );
  AND2_X1 U218 ( .A1(N125), .A2(n172), .ZN(N37) );
  NOR3_X1 U219 ( .A1(N125), .A2(n193), .A3(n208), .ZN(n58) );
  NAND4_X1 U220 ( .A1(n235), .A2(n236), .A3(n1110), .A4(n94), .ZN(n48) );
  OR3_X1 U221 ( .A1(n99), .A2(n79), .A3(n101), .ZN(n35) );
  XOR2_X1 U222 ( .A(add_166_carry[5]), .B(n193), .Z(N130) );
  OR3_X1 U223 ( .A1(n163), .A2(n179), .A3(n250), .ZN(n224) );
  AOI211_X1 U224 ( .C1(n201), .C2(n224), .A(n181), .B(n195), .ZN(n226) );
  NOR3_X1 U225 ( .A1(n158), .A2(n177), .A3(n185), .ZN(n225) );
  NAND2_X1 U226 ( .A1(n226), .A2(n225), .ZN(N120) );
endmodule


module write_out_ARRAY_SIZE8_OUTPUT_DATA_WIDTH16 ( clk, srstn, 
        sram_write_enable, data_set, matrix_index, quantized_data, 
        sram_write_enable_a0, sram_wdata_a, sram_waddr_a, sram_write_enable_b0, 
        sram_wdata_b, sram_waddr_b, sram_write_enable_c0, sram_wdata_c, 
        sram_waddr_c );
  input [1:0] data_set;
  input [5:0] matrix_index;
  input [127:0] quantized_data;
  output [127:0] sram_wdata_a;
  output [5:0] sram_waddr_a;
  output [127:0] sram_wdata_b;
  output [5:0] sram_waddr_b;
  output [127:0] sram_wdata_c;
  output [5:0] sram_waddr_c;
  input clk, srstn, sram_write_enable;
  output sram_write_enable_a0, sram_write_enable_b0, sram_write_enable_c0;
  wire   N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N121,
         N122, N123, N124, N125, N126, N127, N128, N129, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N499, N500, N501,
         N502, N503, N504, N924, N925, N926, N927, N928, N929, N930, N931,
         N932, N933, N934, N935, N936, N937, N938, N939, N1228, N1229, N1539,
         N1547, N1548, N1549, N1550, N1551, N1552, N1553, N1554, N1555, N1556,
         N1557, N1558, N1559, N1560, N1561, N1562, N1581, N1582, N1583, N1584,
         N1585, N1586, N1587, N1588, N1589, N1590, N1591, N1592, N1593, N1594,
         N1595, N1596, N1623, N1624, N1625, N1626, N1627, N1628, N1629, N1630,
         N1631, N1632, N1633, N1634, N1635, N1636, N1637, N1638, r290_B_3_,
         r298_carry_5_, r317_carry_2_, r317_carry_3_, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n10000, n10100, n10200,
         n10300, n10400, n10500, n10600, n10700, n10800, n10900, n11000,
         n11100, n11200, n11300, n11400, n11500, n11600, n11700, n11800,
         n11900, n12000, n12100, n12200, n12300, n12400, n12500, n12600,
         n12700, n12800, n12900, n13000, n13100, n13200, n13300, n13400,
         n13500, n13600, n13700, n13800, n13900, n14000, n14100, n14200,
         n14300, n14400, n14500, n14600, n14700, n14800, n14900, n15000,
         n15100, n15200, n15300, n15400, n15510, n15630, n15700, n15800,
         n15970, n16000, n16100, n16200, n16390, n16400, n16500, n16600,
         n16700, n16800, n16900, n17000, n17100, n17200, n17300, n17400,
         n17500, n17600, n17700, n17800, n17900, n18000, n18100, n18200,
         n18300, n18400, n18500, n18600, n18700, n18800, n18900, n19000,
         n19100, n19200, n19300, n19400, n19500, n19600, n19700, n19800,
         n19900, n20000, n20100, n20200, n20300, n20400, n20500, n20600,
         n20700, n20800, n20900, n21000, n21100, n21200, n21300, n21400,
         n21500, n21600, n21700, n21800, n21900, n22000, n22100, n22200,
         n22300, n22400, n22500, n22600, n22700, n22800, n22900, n23000,
         n23100, n23200, n23300, n23400, n23500, n23600, n23700, n23800,
         n23900, n24000, n24100, n24200, n24300, n24400, n24500, n24600,
         n24700, n24800, n24900, n25000, n25100, n25200, n25300, n25400,
         n25500, n25600, n25700, n25800, n25900, n26000, n26100, n26200,
         n26300, n26400, n26500, n26600, n26700, n26800, n26900, n27000,
         n27100, n27200, n27300, n27400, n27500, n27600, n27700, n27800,
         n27900, n28000, n28100, n28200, n28300, n28400, n28500, n28600,
         n28700, n28800, n28900, n29000, n29100, n29200, n29300, n29400,
         n29500, n29600, n29700, n29800, n29900, n30000, n30100, n30200,
         n30300, n30400, n30500, n30600, n30700, n30800, n30900, n31000,
         n31100, n31200, n31300, n31400, n31500, n31600, n31700, n31800,
         n31900, n32000, n32100, n32200, n32300, n32400, n32500, n32600,
         n32700, n32800, n32900, n33000, n33100, n33200, n33300, n33400,
         n33500, n33600, n33700, n33800, n33900, n34000, n34100, n34200,
         n34300, n34400, n34500, n34600, n34700, n34800, n34900, n35000,
         n35100, n35200, n35300, n35400, n35500, n35600, n35700, n35800,
         n35900, n36000, n36100, n36200, n36300, n36400, n36500, n36600,
         n36700, n36800, n36900, n37000, n37100, n37200, n37300, n37400,
         n37500, n37600, n37700, n37800, n37900, n38000, n38100, n38200,
         n38300, n38400, n38500, n38600, n38700, n38800, n38900, n39000,
         n39100, n39200, n39300, n39400, n39500, n39600, n39700, n39800,
         n39900, n40000, n40100, n40200, n40300, n40400, n40500, n40600,
         n40700, n40800, n40900, n41000, n41100, n41200, n41300, n41400,
         n41500, n41600, n41700, n41800, n41900, n42000, n42100, n42200,
         n42300, n42400, n42500, n42600, n42700, n42800, n42900, n43000,
         n43100, n43200, n43300, n43400, n43500, n43600, n43700, n43800,
         n43900, n44000, n44100, n44200, n44300, n44400, n44500, n44600,
         n44700, n44800, n44900, n45000, n45100, n45200, n45300, n45400,
         n45500, n45600, n45700, n45800, n45900, n46000, n46100, n46200,
         n46300, n46400, n46500, n46600, n46700, n46800, n46900, n4700, n4710,
         n4720, n4730, n4740, n4750, n4760, n4770, n4780, n4790, n4800, n4810,
         n4820, n4830, n4840, n4850, n4860, n4870, n4880, n4890, n4900, n4910,
         n4920, n493, n494, n495, n496, n497, n498, n4990, n5000, n5010, n5020,
         n5030, n5040, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n9240, n9250, n9260, n9270, n9280, n9290, n9300,
         n9310, n9320, n9330, n9340, n9350, n9360, n9370, n9380, n9390, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n10001, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n10101, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n10201, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n10301, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n10401, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n10501, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n10601, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n10701, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n10801, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n10901, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n11001, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n11101, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n11201, n1121, n1122, n1123, n1124, n1125,
         n1126, n1127, n1128, n1129, n11301, n1131, n1132, n1133, n1134, n1135,
         n1136, n1137, n1138, n1139, n11401, n1141, n1142, n1143, n1144, n1145,
         n1146, n1147, n1148, n1149, n11501, n1151, n1152, n1153, n1154, n1155,
         n1156, n1157, n1158, n1159, n11601, n1161, n1162, n1163, n1164, n1165,
         n1166, n1167, n1168, n1169, n11701, n1171, n1172, n1173, n1174, n1175,
         n1176, n1177, n1178, n1179, n11801, n1181, n1182, n1183, n1184, n1185,
         n1186, n1187, n1188, n1189, n11901, n1191, n1192, n1193, n1194, n1195,
         n1196, n1197, n1198, n1199, n12001, n1201, n1202, n1203, n1204, n1205,
         n1206, n1207, n1208, n1209, n12101, n1211, n1212, n1213, n1214, n1215,
         n1216, n1217, n1218, n1219, n12201, n1221, n1222, n1223, n1224,
         n12250, n12260, n1227, n12280, n12290, n12301, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n12401, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n12501, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n12601, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n12701, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n12801, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n12901, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n13001, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n13101, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n13201, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n13301, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n13401, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n13501, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n13601, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n13701, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n13801, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n13901, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n14001, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n14101, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n14201, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n14301, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n14401, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n14501, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n14601, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n14701, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n14801, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n14901, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n15001, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n15101, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n15201, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n15301, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n15390, n15401, n1541, n1542,
         n1543, n1544, n1545, n1546, n15470, n15480, n15490, n15500, n15511,
         n15520, n15530, n15540, n15550, n15560, n15570, n15580, n15590,
         n15600, n15610, n15620, n15631, n1564, n1565, n1566, n1567, n1568,
         n1569, n15701, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n15801, n15810, n15820, n15830, n15840, n15850, n15860, n15870,
         n15880, n15890, n15900, n15910, n15920, n15930, n15940, n15950,
         n15960, n15971, n1598, n1599, n16001, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n16101, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n16201, n1621, n1622, n16230,
         n16240, n16250, n16260, n16270, n16280, n16290, n16300, n16310,
         n16320, n16330, n16340, n16350, n16360, n16370, n16380, n16391,
         n16401, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n16501, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n16601, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n16701, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n16801, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n16901, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n17001, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n17101, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n17201, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n17301, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n17401, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n17501, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n17601, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n17701, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n17801, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n17901, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n18001, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n18101, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n18201, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n18301, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n18401, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n18501, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n18601, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n18701, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n18801, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n18901, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n19001, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n19101, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n19201, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n19301, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n19401, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n19501, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n19601, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n19701, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n19801, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n19901, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n20001, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n20101, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n20201, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n20301, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n20401, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n20501, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n20601, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n20701, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n20801, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n20901, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n21001, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n21101, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n21201, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n21301, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n21401, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n21501, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n21601, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n21701, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n21801, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n21901, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n22001, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n22101, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n22201, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n22301, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n22401, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n22501, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n22601, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n22701, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n22801, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n22901, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n23001, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n23101, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n23201, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n23301, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n23401, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n23501, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n23601, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n23701, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n23801, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n23901, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n24001, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n24101, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n24201, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n24301, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n24401, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n24501, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n24601, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n24701, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n24801, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n24901, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n25001, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n25101, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n25201, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n25301, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539,
         n25401, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549,
         n25501, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559,
         n25601, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569,
         n25701, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579,
         n25801, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589,
         n25901, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599,
         n26001, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609,
         n26101, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619,
         n26201, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629,
         n26301, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639,
         n26401, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649,
         n26501, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659,
         n26601, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669,
         n26701, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679,
         n26801, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689,
         n26901, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699,
         n27001, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709,
         n27101, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719,
         n27201, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729,
         n27301, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739,
         n27401, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749,
         n27501, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759,
         n27601, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769,
         n27701, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779,
         n27801, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789,
         n27901, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799,
         n28001, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809,
         n28101, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819,
         n28201, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829,
         n28301, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839,
         n28401, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849,
         n28501, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859,
         n28601, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869,
         n28701, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879,
         n28801, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889,
         n28901, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899,
         n29001, n2901, n29020, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n29101, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n29201, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n29301, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n29401, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n29501, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n29601, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n29701, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n29801, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n29901, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n30001, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n30101, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n30201, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n30301, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n30401, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n30501, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n30601, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n30701, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n30801, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n30901, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n31001, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n31101, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n31201, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n31301, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n31401, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n31501, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n31601, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n31701, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n31801, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n31901, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n32001, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n32101, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n32201, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n32301, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n32401, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n32501, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n32601, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n32701, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n32801, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n32901, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n33001, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n33101, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n33201, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n33301, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n33401, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n33501, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n33601, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n33701, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n33801, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n33901, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n34001, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n34101, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n34201, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n34301, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n34401, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n34501, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n34601, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n34701, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n34801, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n34901, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n35001, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n35101, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n35201, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n35301, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n35401, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n35501, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n35601, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n35701, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n35801, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n35901, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n36001, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n36101, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n36201, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n36301, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n36401, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n36501, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n36601, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n36701, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n36801, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n36901, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n37001, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n37101, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n37201, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n37301, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n37401, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n37501, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n37601, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n37701, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n37801, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n37901, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n38001, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n38101, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n38201, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n38301, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n38401, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n38501, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n38601, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n38701, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n38801, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n38901, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n39001, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n39101, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n39201, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n39301, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n39401, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n39501, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n39601, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n39701, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n39801, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n39901, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n40001, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n40101, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n40201, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n40301, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n40401, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n40501, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n40601, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n40701, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n40801, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n40901, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n41001, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n41101, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n41201, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n41301, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n41401, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n41501, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n41601, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n41701, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n41801, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n41901, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n42001, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n42101, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n42201, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n42301, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n42401, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n42501, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n42601, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n42701, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n42801, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n42901, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n43001, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n43101, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n43201, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n43301, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n43401, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n43501, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n43601, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n43701, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n43801, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n43901, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n44001, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n44101, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n44201, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n44301, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n44401, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n44501, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n44601, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n44701, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n44801, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n44901, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n45001, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n45101, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n45201, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n45301, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n45401, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n45501, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n45601, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n45701, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n45801, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n45901, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n46001, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n46101, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n46201, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n46301, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n46401, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n46501, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n46601, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n46701, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n46801, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n46901;

  DFF_X1 sram_waddr_b_reg_5_ ( .D(n4686), .CK(clk), .Q(sram_waddr_b[5]) );
  DFF_X1 sram_waddr_b_reg_4_ ( .D(n4687), .CK(clk), .Q(sram_waddr_b[4]) );
  DFF_X1 sram_waddr_b_reg_3_ ( .D(n4689), .CK(clk), .Q(sram_waddr_b[3]) );
  DFF_X1 sram_waddr_b_reg_2_ ( .D(n4688), .CK(clk), .Q(sram_waddr_b[2]) );
  DFF_X1 sram_waddr_b_reg_1_ ( .D(n4685), .CK(clk), .Q(sram_waddr_b[1]) );
  DFF_X1 sram_waddr_b_reg_0_ ( .D(n46901), .CK(clk), .Q(sram_waddr_b[0]) );
  DFF_X1 sram_waddr_c_reg_5_ ( .D(N504), .CK(clk), .Q(sram_waddr_c[5]) );
  DFF_X1 sram_waddr_c_reg_4_ ( .D(N503), .CK(clk), .Q(sram_waddr_c[4]) );
  DFF_X1 sram_waddr_c_reg_3_ ( .D(N502), .CK(clk), .Q(sram_waddr_c[3]) );
  DFF_X1 sram_waddr_c_reg_2_ ( .D(N501), .CK(clk), .Q(sram_waddr_c[2]) );
  DFF_X1 sram_waddr_c_reg_1_ ( .D(N500), .CK(clk), .Q(sram_waddr_c[1]) );
  DFF_X1 sram_waddr_c_reg_0_ ( .D(N499), .CK(clk), .Q(sram_waddr_c[0]) );
  DFF_X1 sram_write_enable_a0_reg ( .D(n1532), .CK(clk), .Q(
        sram_write_enable_a0) );
  DFF_X1 sram_write_enable_b0_reg ( .D(N101), .CK(clk), .Q(
        sram_write_enable_b0) );
  DFF_X1 sram_write_enable_c0_reg ( .D(n1527), .CK(clk), .Q(
        sram_write_enable_c0) );
  DFF_X1 sram_wdata_a_reg_127_ ( .D(N230), .CK(clk), .Q(sram_wdata_a[127]) );
  DFF_X1 sram_wdata_a_reg_126_ ( .D(N229), .CK(clk), .Q(sram_wdata_a[126]) );
  DFF_X1 sram_wdata_a_reg_125_ ( .D(N228), .CK(clk), .Q(sram_wdata_a[125]) );
  DFF_X1 sram_wdata_a_reg_124_ ( .D(N227), .CK(clk), .Q(sram_wdata_a[124]) );
  DFF_X1 sram_wdata_a_reg_123_ ( .D(N226), .CK(clk), .Q(sram_wdata_a[123]) );
  DFF_X1 sram_wdata_a_reg_122_ ( .D(N225), .CK(clk), .Q(sram_wdata_a[122]) );
  DFF_X1 sram_wdata_a_reg_121_ ( .D(N224), .CK(clk), .Q(sram_wdata_a[121]) );
  DFF_X1 sram_wdata_a_reg_120_ ( .D(N223), .CK(clk), .Q(sram_wdata_a[120]) );
  DFF_X1 sram_wdata_a_reg_119_ ( .D(N222), .CK(clk), .Q(sram_wdata_a[119]) );
  DFF_X1 sram_wdata_a_reg_118_ ( .D(N221), .CK(clk), .Q(sram_wdata_a[118]) );
  DFF_X1 sram_wdata_a_reg_117_ ( .D(N220), .CK(clk), .Q(sram_wdata_a[117]) );
  DFF_X1 sram_wdata_a_reg_116_ ( .D(N219), .CK(clk), .Q(sram_wdata_a[116]) );
  DFF_X1 sram_wdata_a_reg_115_ ( .D(N218), .CK(clk), .Q(sram_wdata_a[115]) );
  DFF_X1 sram_wdata_a_reg_114_ ( .D(N217), .CK(clk), .Q(sram_wdata_a[114]) );
  DFF_X1 sram_wdata_a_reg_113_ ( .D(N216), .CK(clk), .Q(sram_wdata_a[113]) );
  DFF_X1 sram_wdata_a_reg_112_ ( .D(N215), .CK(clk), .Q(sram_wdata_a[112]) );
  DFF_X1 sram_wdata_a_reg_111_ ( .D(N214), .CK(clk), .Q(sram_wdata_a[111]) );
  DFF_X1 sram_wdata_a_reg_110_ ( .D(N213), .CK(clk), .Q(sram_wdata_a[110]) );
  DFF_X1 sram_wdata_a_reg_109_ ( .D(N212), .CK(clk), .Q(sram_wdata_a[109]) );
  DFF_X1 sram_wdata_a_reg_108_ ( .D(N211), .CK(clk), .Q(sram_wdata_a[108]) );
  DFF_X1 sram_wdata_a_reg_107_ ( .D(N210), .CK(clk), .Q(sram_wdata_a[107]) );
  DFF_X1 sram_wdata_a_reg_106_ ( .D(N209), .CK(clk), .Q(sram_wdata_a[106]) );
  DFF_X1 sram_wdata_a_reg_105_ ( .D(N208), .CK(clk), .Q(sram_wdata_a[105]) );
  DFF_X1 sram_wdata_a_reg_104_ ( .D(N207), .CK(clk), .Q(sram_wdata_a[104]) );
  DFF_X1 sram_wdata_a_reg_103_ ( .D(N206), .CK(clk), .Q(sram_wdata_a[103]) );
  DFF_X1 sram_wdata_a_reg_102_ ( .D(N205), .CK(clk), .Q(sram_wdata_a[102]) );
  DFF_X1 sram_wdata_a_reg_101_ ( .D(N204), .CK(clk), .Q(sram_wdata_a[101]) );
  DFF_X1 sram_wdata_a_reg_100_ ( .D(N203), .CK(clk), .Q(sram_wdata_a[100]) );
  DFF_X1 sram_wdata_a_reg_99_ ( .D(N202), .CK(clk), .Q(sram_wdata_a[99]) );
  DFF_X1 sram_wdata_a_reg_98_ ( .D(N201), .CK(clk), .Q(sram_wdata_a[98]) );
  DFF_X1 sram_wdata_a_reg_97_ ( .D(N200), .CK(clk), .Q(sram_wdata_a[97]) );
  DFF_X1 sram_wdata_a_reg_96_ ( .D(N199), .CK(clk), .Q(sram_wdata_a[96]) );
  DFF_X1 sram_wdata_a_reg_95_ ( .D(N198), .CK(clk), .Q(sram_wdata_a[95]) );
  DFF_X1 sram_wdata_a_reg_94_ ( .D(N197), .CK(clk), .Q(sram_wdata_a[94]) );
  DFF_X1 sram_wdata_a_reg_93_ ( .D(N196), .CK(clk), .Q(sram_wdata_a[93]) );
  DFF_X1 sram_wdata_a_reg_92_ ( .D(N195), .CK(clk), .Q(sram_wdata_a[92]) );
  DFF_X1 sram_wdata_a_reg_91_ ( .D(N194), .CK(clk), .Q(sram_wdata_a[91]) );
  DFF_X1 sram_wdata_a_reg_90_ ( .D(N193), .CK(clk), .Q(sram_wdata_a[90]) );
  DFF_X1 sram_wdata_a_reg_89_ ( .D(N192), .CK(clk), .Q(sram_wdata_a[89]) );
  DFF_X1 sram_wdata_a_reg_88_ ( .D(N191), .CK(clk), .Q(sram_wdata_a[88]) );
  DFF_X1 sram_wdata_a_reg_87_ ( .D(N190), .CK(clk), .Q(sram_wdata_a[87]) );
  DFF_X1 sram_wdata_a_reg_86_ ( .D(N189), .CK(clk), .Q(sram_wdata_a[86]) );
  DFF_X1 sram_wdata_a_reg_85_ ( .D(N188), .CK(clk), .Q(sram_wdata_a[85]) );
  DFF_X1 sram_wdata_a_reg_84_ ( .D(N187), .CK(clk), .Q(sram_wdata_a[84]) );
  DFF_X1 sram_wdata_a_reg_83_ ( .D(N186), .CK(clk), .Q(sram_wdata_a[83]) );
  DFF_X1 sram_wdata_a_reg_82_ ( .D(N185), .CK(clk), .Q(sram_wdata_a[82]) );
  DFF_X1 sram_wdata_a_reg_81_ ( .D(N184), .CK(clk), .Q(sram_wdata_a[81]) );
  DFF_X1 sram_wdata_a_reg_80_ ( .D(N183), .CK(clk), .Q(sram_wdata_a[80]) );
  DFF_X1 sram_wdata_a_reg_79_ ( .D(N182), .CK(clk), .Q(sram_wdata_a[79]) );
  DFF_X1 sram_wdata_a_reg_78_ ( .D(N181), .CK(clk), .Q(sram_wdata_a[78]) );
  DFF_X1 sram_wdata_a_reg_77_ ( .D(N180), .CK(clk), .Q(sram_wdata_a[77]) );
  DFF_X1 sram_wdata_a_reg_76_ ( .D(N179), .CK(clk), .Q(sram_wdata_a[76]) );
  DFF_X1 sram_wdata_a_reg_75_ ( .D(N178), .CK(clk), .Q(sram_wdata_a[75]) );
  DFF_X1 sram_wdata_a_reg_74_ ( .D(N177), .CK(clk), .Q(sram_wdata_a[74]) );
  DFF_X1 sram_wdata_a_reg_73_ ( .D(N176), .CK(clk), .Q(sram_wdata_a[73]) );
  DFF_X1 sram_wdata_a_reg_72_ ( .D(N175), .CK(clk), .Q(sram_wdata_a[72]) );
  DFF_X1 sram_wdata_a_reg_71_ ( .D(N174), .CK(clk), .Q(sram_wdata_a[71]) );
  DFF_X1 sram_wdata_a_reg_70_ ( .D(N173), .CK(clk), .Q(sram_wdata_a[70]) );
  DFF_X1 sram_wdata_a_reg_69_ ( .D(N172), .CK(clk), .Q(sram_wdata_a[69]) );
  DFF_X1 sram_wdata_a_reg_68_ ( .D(N171), .CK(clk), .Q(sram_wdata_a[68]) );
  DFF_X1 sram_wdata_a_reg_67_ ( .D(N170), .CK(clk), .Q(sram_wdata_a[67]) );
  DFF_X1 sram_wdata_a_reg_66_ ( .D(N169), .CK(clk), .Q(sram_wdata_a[66]) );
  DFF_X1 sram_wdata_a_reg_65_ ( .D(N168), .CK(clk), .Q(sram_wdata_a[65]) );
  DFF_X1 sram_wdata_a_reg_64_ ( .D(N167), .CK(clk), .Q(sram_wdata_a[64]) );
  DFF_X1 sram_wdata_a_reg_63_ ( .D(N166), .CK(clk), .Q(sram_wdata_a[63]) );
  DFF_X1 sram_wdata_a_reg_62_ ( .D(N165), .CK(clk), .Q(sram_wdata_a[62]) );
  DFF_X1 sram_wdata_a_reg_61_ ( .D(N164), .CK(clk), .Q(sram_wdata_a[61]) );
  DFF_X1 sram_wdata_a_reg_60_ ( .D(N163), .CK(clk), .Q(sram_wdata_a[60]) );
  DFF_X1 sram_wdata_a_reg_59_ ( .D(N162), .CK(clk), .Q(sram_wdata_a[59]) );
  DFF_X1 sram_wdata_a_reg_58_ ( .D(N161), .CK(clk), .Q(sram_wdata_a[58]) );
  DFF_X1 sram_wdata_a_reg_57_ ( .D(N160), .CK(clk), .Q(sram_wdata_a[57]) );
  DFF_X1 sram_wdata_a_reg_56_ ( .D(N159), .CK(clk), .Q(sram_wdata_a[56]) );
  DFF_X1 sram_wdata_a_reg_55_ ( .D(N158), .CK(clk), .Q(sram_wdata_a[55]) );
  DFF_X1 sram_wdata_a_reg_54_ ( .D(N157), .CK(clk), .Q(sram_wdata_a[54]) );
  DFF_X1 sram_wdata_a_reg_53_ ( .D(N156), .CK(clk), .Q(sram_wdata_a[53]) );
  DFF_X1 sram_wdata_a_reg_52_ ( .D(N155), .CK(clk), .Q(sram_wdata_a[52]) );
  DFF_X1 sram_wdata_a_reg_51_ ( .D(N154), .CK(clk), .Q(sram_wdata_a[51]) );
  DFF_X1 sram_wdata_a_reg_50_ ( .D(N153), .CK(clk), .Q(sram_wdata_a[50]) );
  DFF_X1 sram_wdata_a_reg_49_ ( .D(N152), .CK(clk), .Q(sram_wdata_a[49]) );
  DFF_X1 sram_wdata_a_reg_48_ ( .D(N151), .CK(clk), .Q(sram_wdata_a[48]) );
  DFF_X1 sram_wdata_a_reg_47_ ( .D(N150), .CK(clk), .Q(sram_wdata_a[47]) );
  DFF_X1 sram_wdata_a_reg_46_ ( .D(N149), .CK(clk), .Q(sram_wdata_a[46]) );
  DFF_X1 sram_wdata_a_reg_45_ ( .D(N148), .CK(clk), .Q(sram_wdata_a[45]) );
  DFF_X1 sram_wdata_a_reg_44_ ( .D(N147), .CK(clk), .Q(sram_wdata_a[44]) );
  DFF_X1 sram_wdata_a_reg_43_ ( .D(N146), .CK(clk), .Q(sram_wdata_a[43]) );
  DFF_X1 sram_wdata_a_reg_42_ ( .D(N145), .CK(clk), .Q(sram_wdata_a[42]) );
  DFF_X1 sram_wdata_a_reg_41_ ( .D(N144), .CK(clk), .Q(sram_wdata_a[41]) );
  DFF_X1 sram_wdata_a_reg_40_ ( .D(N143), .CK(clk), .Q(sram_wdata_a[40]) );
  DFF_X1 sram_wdata_a_reg_39_ ( .D(N142), .CK(clk), .Q(sram_wdata_a[39]) );
  DFF_X1 sram_wdata_a_reg_38_ ( .D(N141), .CK(clk), .Q(sram_wdata_a[38]) );
  DFF_X1 sram_wdata_a_reg_37_ ( .D(N140), .CK(clk), .Q(sram_wdata_a[37]) );
  DFF_X1 sram_wdata_a_reg_36_ ( .D(N139), .CK(clk), .Q(sram_wdata_a[36]) );
  DFF_X1 sram_wdata_a_reg_35_ ( .D(N138), .CK(clk), .Q(sram_wdata_a[35]) );
  DFF_X1 sram_wdata_a_reg_34_ ( .D(N137), .CK(clk), .Q(sram_wdata_a[34]) );
  DFF_X1 sram_wdata_a_reg_33_ ( .D(N136), .CK(clk), .Q(sram_wdata_a[33]) );
  DFF_X1 sram_wdata_a_reg_32_ ( .D(N135), .CK(clk), .Q(sram_wdata_a[32]) );
  DFF_X1 sram_wdata_a_reg_31_ ( .D(N134), .CK(clk), .Q(sram_wdata_a[31]) );
  DFF_X1 sram_wdata_a_reg_30_ ( .D(N133), .CK(clk), .Q(sram_wdata_a[30]) );
  DFF_X1 sram_wdata_a_reg_29_ ( .D(N132), .CK(clk), .Q(sram_wdata_a[29]) );
  DFF_X1 sram_wdata_a_reg_28_ ( .D(N131), .CK(clk), .Q(sram_wdata_a[28]) );
  DFF_X1 sram_wdata_a_reg_27_ ( .D(N130), .CK(clk), .Q(sram_wdata_a[27]) );
  DFF_X1 sram_wdata_a_reg_26_ ( .D(N129), .CK(clk), .Q(sram_wdata_a[26]) );
  DFF_X1 sram_wdata_a_reg_25_ ( .D(N128), .CK(clk), .Q(sram_wdata_a[25]) );
  DFF_X1 sram_wdata_a_reg_24_ ( .D(N127), .CK(clk), .Q(sram_wdata_a[24]) );
  DFF_X1 sram_wdata_a_reg_23_ ( .D(N126), .CK(clk), .Q(sram_wdata_a[23]) );
  DFF_X1 sram_wdata_a_reg_22_ ( .D(N125), .CK(clk), .Q(sram_wdata_a[22]) );
  DFF_X1 sram_wdata_a_reg_21_ ( .D(N124), .CK(clk), .Q(sram_wdata_a[21]) );
  DFF_X1 sram_wdata_a_reg_20_ ( .D(N123), .CK(clk), .Q(sram_wdata_a[20]) );
  DFF_X1 sram_wdata_a_reg_19_ ( .D(N122), .CK(clk), .Q(sram_wdata_a[19]) );
  DFF_X1 sram_wdata_a_reg_18_ ( .D(N121), .CK(clk), .Q(sram_wdata_a[18]) );
  DFF_X1 sram_wdata_a_reg_17_ ( .D(N120), .CK(clk), .Q(sram_wdata_a[17]) );
  DFF_X1 sram_wdata_a_reg_16_ ( .D(N119), .CK(clk), .Q(sram_wdata_a[16]) );
  DFF_X1 sram_wdata_a_reg_15_ ( .D(N118), .CK(clk), .Q(sram_wdata_a[15]) );
  DFF_X1 sram_wdata_a_reg_14_ ( .D(N117), .CK(clk), .Q(sram_wdata_a[14]) );
  DFF_X1 sram_wdata_a_reg_13_ ( .D(N116), .CK(clk), .Q(sram_wdata_a[13]) );
  DFF_X1 sram_wdata_a_reg_12_ ( .D(N115), .CK(clk), .Q(sram_wdata_a[12]) );
  DFF_X1 sram_wdata_a_reg_11_ ( .D(N114), .CK(clk), .Q(sram_wdata_a[11]) );
  DFF_X1 sram_wdata_a_reg_10_ ( .D(N113), .CK(clk), .Q(sram_wdata_a[10]) );
  DFF_X1 sram_wdata_a_reg_9_ ( .D(N112), .CK(clk), .Q(sram_wdata_a[9]) );
  DFF_X1 sram_wdata_a_reg_8_ ( .D(N111), .CK(clk), .Q(sram_wdata_a[8]) );
  DFF_X1 sram_wdata_a_reg_7_ ( .D(N110), .CK(clk), .Q(sram_wdata_a[7]) );
  DFF_X1 sram_wdata_a_reg_6_ ( .D(N109), .CK(clk), .Q(sram_wdata_a[6]) );
  DFF_X1 sram_wdata_a_reg_5_ ( .D(N108), .CK(clk), .Q(sram_wdata_a[5]) );
  DFF_X1 sram_wdata_a_reg_4_ ( .D(N107), .CK(clk), .Q(sram_wdata_a[4]) );
  DFF_X1 sram_wdata_a_reg_3_ ( .D(N106), .CK(clk), .Q(sram_wdata_a[3]) );
  DFF_X1 sram_wdata_a_reg_2_ ( .D(N105), .CK(clk), .Q(sram_wdata_a[2]) );
  DFF_X1 sram_wdata_a_reg_1_ ( .D(N104), .CK(clk), .Q(sram_wdata_a[1]) );
  DFF_X1 sram_wdata_a_reg_0_ ( .D(N103), .CK(clk), .Q(sram_wdata_a[0]) );
  DFF_X1 sram_wdata_b_reg_127_ ( .D(N358), .CK(clk), .Q(sram_wdata_b[127]) );
  DFF_X1 sram_wdata_b_reg_126_ ( .D(N357), .CK(clk), .Q(sram_wdata_b[126]) );
  DFF_X1 sram_wdata_b_reg_125_ ( .D(N356), .CK(clk), .Q(sram_wdata_b[125]) );
  DFF_X1 sram_wdata_b_reg_124_ ( .D(N355), .CK(clk), .Q(sram_wdata_b[124]) );
  DFF_X1 sram_wdata_b_reg_123_ ( .D(N354), .CK(clk), .Q(sram_wdata_b[123]) );
  DFF_X1 sram_wdata_b_reg_122_ ( .D(N353), .CK(clk), .Q(sram_wdata_b[122]) );
  DFF_X1 sram_wdata_b_reg_121_ ( .D(N352), .CK(clk), .Q(sram_wdata_b[121]) );
  DFF_X1 sram_wdata_b_reg_120_ ( .D(N351), .CK(clk), .Q(sram_wdata_b[120]) );
  DFF_X1 sram_wdata_b_reg_119_ ( .D(N350), .CK(clk), .Q(sram_wdata_b[119]) );
  DFF_X1 sram_wdata_b_reg_118_ ( .D(N349), .CK(clk), .Q(sram_wdata_b[118]) );
  DFF_X1 sram_wdata_b_reg_117_ ( .D(N348), .CK(clk), .Q(sram_wdata_b[117]) );
  DFF_X1 sram_wdata_b_reg_116_ ( .D(N347), .CK(clk), .Q(sram_wdata_b[116]) );
  DFF_X1 sram_wdata_b_reg_115_ ( .D(N346), .CK(clk), .Q(sram_wdata_b[115]) );
  DFF_X1 sram_wdata_b_reg_114_ ( .D(N345), .CK(clk), .Q(sram_wdata_b[114]) );
  DFF_X1 sram_wdata_b_reg_113_ ( .D(N344), .CK(clk), .Q(sram_wdata_b[113]) );
  DFF_X1 sram_wdata_b_reg_112_ ( .D(N343), .CK(clk), .Q(sram_wdata_b[112]) );
  DFF_X1 sram_wdata_b_reg_111_ ( .D(N342), .CK(clk), .Q(sram_wdata_b[111]) );
  DFF_X1 sram_wdata_b_reg_110_ ( .D(N341), .CK(clk), .Q(sram_wdata_b[110]) );
  DFF_X1 sram_wdata_b_reg_109_ ( .D(N340), .CK(clk), .Q(sram_wdata_b[109]) );
  DFF_X1 sram_wdata_b_reg_108_ ( .D(N339), .CK(clk), .Q(sram_wdata_b[108]) );
  DFF_X1 sram_wdata_b_reg_107_ ( .D(N338), .CK(clk), .Q(sram_wdata_b[107]) );
  DFF_X1 sram_wdata_b_reg_106_ ( .D(N337), .CK(clk), .Q(sram_wdata_b[106]) );
  DFF_X1 sram_wdata_b_reg_105_ ( .D(N336), .CK(clk), .Q(sram_wdata_b[105]) );
  DFF_X1 sram_wdata_b_reg_104_ ( .D(N335), .CK(clk), .Q(sram_wdata_b[104]) );
  DFF_X1 sram_wdata_b_reg_103_ ( .D(N334), .CK(clk), .Q(sram_wdata_b[103]) );
  DFF_X1 sram_wdata_b_reg_102_ ( .D(N333), .CK(clk), .Q(sram_wdata_b[102]) );
  DFF_X1 sram_wdata_b_reg_101_ ( .D(N332), .CK(clk), .Q(sram_wdata_b[101]) );
  DFF_X1 sram_wdata_b_reg_100_ ( .D(N331), .CK(clk), .Q(sram_wdata_b[100]) );
  DFF_X1 sram_wdata_b_reg_99_ ( .D(N330), .CK(clk), .Q(sram_wdata_b[99]) );
  DFF_X1 sram_wdata_b_reg_98_ ( .D(N329), .CK(clk), .Q(sram_wdata_b[98]) );
  DFF_X1 sram_wdata_b_reg_97_ ( .D(N328), .CK(clk), .Q(sram_wdata_b[97]) );
  DFF_X1 sram_wdata_b_reg_96_ ( .D(N327), .CK(clk), .Q(sram_wdata_b[96]) );
  DFF_X1 sram_wdata_b_reg_95_ ( .D(N326), .CK(clk), .Q(sram_wdata_b[95]) );
  DFF_X1 sram_wdata_b_reg_94_ ( .D(N325), .CK(clk), .Q(sram_wdata_b[94]) );
  DFF_X1 sram_wdata_b_reg_93_ ( .D(N324), .CK(clk), .Q(sram_wdata_b[93]) );
  DFF_X1 sram_wdata_b_reg_92_ ( .D(N323), .CK(clk), .Q(sram_wdata_b[92]) );
  DFF_X1 sram_wdata_b_reg_91_ ( .D(N322), .CK(clk), .Q(sram_wdata_b[91]) );
  DFF_X1 sram_wdata_b_reg_90_ ( .D(N321), .CK(clk), .Q(sram_wdata_b[90]) );
  DFF_X1 sram_wdata_b_reg_89_ ( .D(N320), .CK(clk), .Q(sram_wdata_b[89]) );
  DFF_X1 sram_wdata_b_reg_88_ ( .D(N319), .CK(clk), .Q(sram_wdata_b[88]) );
  DFF_X1 sram_wdata_b_reg_87_ ( .D(N318), .CK(clk), .Q(sram_wdata_b[87]) );
  DFF_X1 sram_wdata_b_reg_86_ ( .D(N317), .CK(clk), .Q(sram_wdata_b[86]) );
  DFF_X1 sram_wdata_b_reg_85_ ( .D(N316), .CK(clk), .Q(sram_wdata_b[85]) );
  DFF_X1 sram_wdata_b_reg_84_ ( .D(N315), .CK(clk), .Q(sram_wdata_b[84]) );
  DFF_X1 sram_wdata_b_reg_83_ ( .D(N314), .CK(clk), .Q(sram_wdata_b[83]) );
  DFF_X1 sram_wdata_b_reg_82_ ( .D(N313), .CK(clk), .Q(sram_wdata_b[82]) );
  DFF_X1 sram_wdata_b_reg_81_ ( .D(N312), .CK(clk), .Q(sram_wdata_b[81]) );
  DFF_X1 sram_wdata_b_reg_80_ ( .D(N311), .CK(clk), .Q(sram_wdata_b[80]) );
  DFF_X1 sram_wdata_b_reg_79_ ( .D(N310), .CK(clk), .Q(sram_wdata_b[79]) );
  DFF_X1 sram_wdata_b_reg_78_ ( .D(N309), .CK(clk), .Q(sram_wdata_b[78]) );
  DFF_X1 sram_wdata_b_reg_77_ ( .D(N308), .CK(clk), .Q(sram_wdata_b[77]) );
  DFF_X1 sram_wdata_b_reg_76_ ( .D(N307), .CK(clk), .Q(sram_wdata_b[76]) );
  DFF_X1 sram_wdata_b_reg_75_ ( .D(N306), .CK(clk), .Q(sram_wdata_b[75]) );
  DFF_X1 sram_wdata_b_reg_74_ ( .D(N305), .CK(clk), .Q(sram_wdata_b[74]) );
  DFF_X1 sram_wdata_b_reg_73_ ( .D(N304), .CK(clk), .Q(sram_wdata_b[73]) );
  DFF_X1 sram_wdata_b_reg_72_ ( .D(N303), .CK(clk), .Q(sram_wdata_b[72]) );
  DFF_X1 sram_wdata_b_reg_71_ ( .D(N302), .CK(clk), .Q(sram_wdata_b[71]) );
  DFF_X1 sram_wdata_b_reg_70_ ( .D(N301), .CK(clk), .Q(sram_wdata_b[70]) );
  DFF_X1 sram_wdata_b_reg_69_ ( .D(N300), .CK(clk), .Q(sram_wdata_b[69]) );
  DFF_X1 sram_wdata_b_reg_68_ ( .D(N299), .CK(clk), .Q(sram_wdata_b[68]) );
  DFF_X1 sram_wdata_b_reg_67_ ( .D(N298), .CK(clk), .Q(sram_wdata_b[67]) );
  DFF_X1 sram_wdata_b_reg_66_ ( .D(N297), .CK(clk), .Q(sram_wdata_b[66]) );
  DFF_X1 sram_wdata_b_reg_65_ ( .D(N296), .CK(clk), .Q(sram_wdata_b[65]) );
  DFF_X1 sram_wdata_b_reg_64_ ( .D(N295), .CK(clk), .Q(sram_wdata_b[64]) );
  DFF_X1 sram_wdata_b_reg_63_ ( .D(N294), .CK(clk), .Q(sram_wdata_b[63]) );
  DFF_X1 sram_wdata_b_reg_62_ ( .D(N293), .CK(clk), .Q(sram_wdata_b[62]) );
  DFF_X1 sram_wdata_b_reg_61_ ( .D(N292), .CK(clk), .Q(sram_wdata_b[61]) );
  DFF_X1 sram_wdata_b_reg_60_ ( .D(N291), .CK(clk), .Q(sram_wdata_b[60]) );
  DFF_X1 sram_wdata_b_reg_59_ ( .D(N290), .CK(clk), .Q(sram_wdata_b[59]) );
  DFF_X1 sram_wdata_b_reg_58_ ( .D(N289), .CK(clk), .Q(sram_wdata_b[58]) );
  DFF_X1 sram_wdata_b_reg_57_ ( .D(N288), .CK(clk), .Q(sram_wdata_b[57]) );
  DFF_X1 sram_wdata_b_reg_56_ ( .D(N287), .CK(clk), .Q(sram_wdata_b[56]) );
  DFF_X1 sram_wdata_b_reg_55_ ( .D(N286), .CK(clk), .Q(sram_wdata_b[55]) );
  DFF_X1 sram_wdata_b_reg_54_ ( .D(N285), .CK(clk), .Q(sram_wdata_b[54]) );
  DFF_X1 sram_wdata_b_reg_53_ ( .D(N284), .CK(clk), .Q(sram_wdata_b[53]) );
  DFF_X1 sram_wdata_b_reg_52_ ( .D(N283), .CK(clk), .Q(sram_wdata_b[52]) );
  DFF_X1 sram_wdata_b_reg_51_ ( .D(N282), .CK(clk), .Q(sram_wdata_b[51]) );
  DFF_X1 sram_wdata_b_reg_50_ ( .D(N281), .CK(clk), .Q(sram_wdata_b[50]) );
  DFF_X1 sram_wdata_b_reg_49_ ( .D(N280), .CK(clk), .Q(sram_wdata_b[49]) );
  DFF_X1 sram_wdata_b_reg_48_ ( .D(N279), .CK(clk), .Q(sram_wdata_b[48]) );
  DFF_X1 sram_wdata_b_reg_47_ ( .D(N278), .CK(clk), .Q(sram_wdata_b[47]) );
  DFF_X1 sram_wdata_b_reg_46_ ( .D(N277), .CK(clk), .Q(sram_wdata_b[46]) );
  DFF_X1 sram_wdata_b_reg_45_ ( .D(N276), .CK(clk), .Q(sram_wdata_b[45]) );
  DFF_X1 sram_wdata_b_reg_44_ ( .D(N275), .CK(clk), .Q(sram_wdata_b[44]) );
  DFF_X1 sram_wdata_b_reg_43_ ( .D(N274), .CK(clk), .Q(sram_wdata_b[43]) );
  DFF_X1 sram_wdata_b_reg_42_ ( .D(N273), .CK(clk), .Q(sram_wdata_b[42]) );
  DFF_X1 sram_wdata_b_reg_41_ ( .D(N272), .CK(clk), .Q(sram_wdata_b[41]) );
  DFF_X1 sram_wdata_b_reg_40_ ( .D(N271), .CK(clk), .Q(sram_wdata_b[40]) );
  DFF_X1 sram_wdata_b_reg_39_ ( .D(N270), .CK(clk), .Q(sram_wdata_b[39]) );
  DFF_X1 sram_wdata_b_reg_38_ ( .D(N269), .CK(clk), .Q(sram_wdata_b[38]) );
  DFF_X1 sram_wdata_b_reg_37_ ( .D(N268), .CK(clk), .Q(sram_wdata_b[37]) );
  DFF_X1 sram_wdata_b_reg_36_ ( .D(N267), .CK(clk), .Q(sram_wdata_b[36]) );
  DFF_X1 sram_wdata_b_reg_35_ ( .D(N266), .CK(clk), .Q(sram_wdata_b[35]) );
  DFF_X1 sram_wdata_b_reg_34_ ( .D(N265), .CK(clk), .Q(sram_wdata_b[34]) );
  DFF_X1 sram_wdata_b_reg_33_ ( .D(N264), .CK(clk), .Q(sram_wdata_b[33]) );
  DFF_X1 sram_wdata_b_reg_32_ ( .D(N263), .CK(clk), .Q(sram_wdata_b[32]) );
  DFF_X1 sram_wdata_b_reg_31_ ( .D(N262), .CK(clk), .Q(sram_wdata_b[31]) );
  DFF_X1 sram_wdata_b_reg_30_ ( .D(N261), .CK(clk), .Q(sram_wdata_b[30]) );
  DFF_X1 sram_wdata_b_reg_29_ ( .D(N260), .CK(clk), .Q(sram_wdata_b[29]) );
  DFF_X1 sram_wdata_b_reg_28_ ( .D(N259), .CK(clk), .Q(sram_wdata_b[28]) );
  DFF_X1 sram_wdata_b_reg_27_ ( .D(N258), .CK(clk), .Q(sram_wdata_b[27]) );
  DFF_X1 sram_wdata_b_reg_26_ ( .D(N257), .CK(clk), .Q(sram_wdata_b[26]) );
  DFF_X1 sram_wdata_b_reg_25_ ( .D(N256), .CK(clk), .Q(sram_wdata_b[25]) );
  DFF_X1 sram_wdata_b_reg_24_ ( .D(N255), .CK(clk), .Q(sram_wdata_b[24]) );
  DFF_X1 sram_wdata_b_reg_23_ ( .D(N254), .CK(clk), .Q(sram_wdata_b[23]) );
  DFF_X1 sram_wdata_b_reg_22_ ( .D(N253), .CK(clk), .Q(sram_wdata_b[22]) );
  DFF_X1 sram_wdata_b_reg_21_ ( .D(N252), .CK(clk), .Q(sram_wdata_b[21]) );
  DFF_X1 sram_wdata_b_reg_20_ ( .D(N251), .CK(clk), .Q(sram_wdata_b[20]) );
  DFF_X1 sram_wdata_b_reg_19_ ( .D(N250), .CK(clk), .Q(sram_wdata_b[19]) );
  DFF_X1 sram_wdata_b_reg_18_ ( .D(N249), .CK(clk), .Q(sram_wdata_b[18]) );
  DFF_X1 sram_wdata_b_reg_17_ ( .D(N248), .CK(clk), .Q(sram_wdata_b[17]) );
  DFF_X1 sram_wdata_b_reg_16_ ( .D(N247), .CK(clk), .Q(sram_wdata_b[16]) );
  DFF_X1 sram_wdata_b_reg_15_ ( .D(N246), .CK(clk), .Q(sram_wdata_b[15]) );
  DFF_X1 sram_wdata_b_reg_14_ ( .D(N245), .CK(clk), .Q(sram_wdata_b[14]) );
  DFF_X1 sram_wdata_b_reg_13_ ( .D(N244), .CK(clk), .Q(sram_wdata_b[13]) );
  DFF_X1 sram_wdata_b_reg_12_ ( .D(N243), .CK(clk), .Q(sram_wdata_b[12]) );
  DFF_X1 sram_wdata_b_reg_11_ ( .D(N242), .CK(clk), .Q(sram_wdata_b[11]) );
  DFF_X1 sram_wdata_b_reg_10_ ( .D(N241), .CK(clk), .Q(sram_wdata_b[10]) );
  DFF_X1 sram_wdata_b_reg_9_ ( .D(N240), .CK(clk), .Q(sram_wdata_b[9]) );
  DFF_X1 sram_wdata_b_reg_8_ ( .D(N239), .CK(clk), .Q(sram_wdata_b[8]) );
  DFF_X1 sram_wdata_b_reg_7_ ( .D(N238), .CK(clk), .Q(sram_wdata_b[7]) );
  DFF_X1 sram_wdata_b_reg_6_ ( .D(N237), .CK(clk), .Q(sram_wdata_b[6]) );
  DFF_X1 sram_wdata_b_reg_5_ ( .D(N236), .CK(clk), .Q(sram_wdata_b[5]) );
  DFF_X1 sram_wdata_b_reg_4_ ( .D(N235), .CK(clk), .Q(sram_wdata_b[4]) );
  DFF_X1 sram_wdata_b_reg_3_ ( .D(N234), .CK(clk), .Q(sram_wdata_b[3]) );
  DFF_X1 sram_wdata_b_reg_2_ ( .D(N233), .CK(clk), .Q(sram_wdata_b[2]) );
  DFF_X1 sram_wdata_b_reg_1_ ( .D(N232), .CK(clk), .Q(sram_wdata_b[1]) );
  DFF_X1 sram_wdata_b_reg_0_ ( .D(N231), .CK(clk), .Q(sram_wdata_b[0]) );
  DFF_X1 sram_wdata_c_reg_127_ ( .D(N486), .CK(clk), .Q(sram_wdata_c[127]) );
  DFF_X1 sram_wdata_c_reg_126_ ( .D(N485), .CK(clk), .Q(sram_wdata_c[126]) );
  DFF_X1 sram_wdata_c_reg_125_ ( .D(N484), .CK(clk), .Q(sram_wdata_c[125]) );
  DFF_X1 sram_wdata_c_reg_124_ ( .D(N483), .CK(clk), .Q(sram_wdata_c[124]) );
  DFF_X1 sram_wdata_c_reg_123_ ( .D(N482), .CK(clk), .Q(sram_wdata_c[123]) );
  DFF_X1 sram_wdata_c_reg_122_ ( .D(N481), .CK(clk), .Q(sram_wdata_c[122]) );
  DFF_X1 sram_wdata_c_reg_121_ ( .D(N480), .CK(clk), .Q(sram_wdata_c[121]) );
  DFF_X1 sram_wdata_c_reg_120_ ( .D(N479), .CK(clk), .Q(sram_wdata_c[120]) );
  DFF_X1 sram_wdata_c_reg_119_ ( .D(N478), .CK(clk), .Q(sram_wdata_c[119]) );
  DFF_X1 sram_wdata_c_reg_118_ ( .D(N477), .CK(clk), .Q(sram_wdata_c[118]) );
  DFF_X1 sram_wdata_c_reg_117_ ( .D(N476), .CK(clk), .Q(sram_wdata_c[117]) );
  DFF_X1 sram_wdata_c_reg_116_ ( .D(N475), .CK(clk), .Q(sram_wdata_c[116]) );
  DFF_X1 sram_wdata_c_reg_115_ ( .D(N474), .CK(clk), .Q(sram_wdata_c[115]) );
  DFF_X1 sram_wdata_c_reg_114_ ( .D(N473), .CK(clk), .Q(sram_wdata_c[114]) );
  DFF_X1 sram_wdata_c_reg_113_ ( .D(N472), .CK(clk), .Q(sram_wdata_c[113]) );
  DFF_X1 sram_wdata_c_reg_112_ ( .D(N471), .CK(clk), .Q(sram_wdata_c[112]) );
  DFF_X1 sram_wdata_c_reg_111_ ( .D(N470), .CK(clk), .Q(sram_wdata_c[111]) );
  DFF_X1 sram_wdata_c_reg_110_ ( .D(N469), .CK(clk), .Q(sram_wdata_c[110]) );
  DFF_X1 sram_wdata_c_reg_109_ ( .D(N468), .CK(clk), .Q(sram_wdata_c[109]) );
  DFF_X1 sram_wdata_c_reg_108_ ( .D(N467), .CK(clk), .Q(sram_wdata_c[108]) );
  DFF_X1 sram_wdata_c_reg_107_ ( .D(N466), .CK(clk), .Q(sram_wdata_c[107]) );
  DFF_X1 sram_wdata_c_reg_106_ ( .D(N465), .CK(clk), .Q(sram_wdata_c[106]) );
  DFF_X1 sram_wdata_c_reg_105_ ( .D(N464), .CK(clk), .Q(sram_wdata_c[105]) );
  DFF_X1 sram_wdata_c_reg_104_ ( .D(N463), .CK(clk), .Q(sram_wdata_c[104]) );
  DFF_X1 sram_wdata_c_reg_103_ ( .D(N462), .CK(clk), .Q(sram_wdata_c[103]) );
  DFF_X1 sram_wdata_c_reg_102_ ( .D(N461), .CK(clk), .Q(sram_wdata_c[102]) );
  DFF_X1 sram_wdata_c_reg_101_ ( .D(N460), .CK(clk), .Q(sram_wdata_c[101]) );
  DFF_X1 sram_wdata_c_reg_100_ ( .D(N459), .CK(clk), .Q(sram_wdata_c[100]) );
  DFF_X1 sram_wdata_c_reg_99_ ( .D(N458), .CK(clk), .Q(sram_wdata_c[99]) );
  DFF_X1 sram_wdata_c_reg_98_ ( .D(N457), .CK(clk), .Q(sram_wdata_c[98]) );
  DFF_X1 sram_wdata_c_reg_97_ ( .D(N456), .CK(clk), .Q(sram_wdata_c[97]) );
  DFF_X1 sram_wdata_c_reg_96_ ( .D(N455), .CK(clk), .Q(sram_wdata_c[96]) );
  DFF_X1 sram_wdata_c_reg_95_ ( .D(N454), .CK(clk), .Q(sram_wdata_c[95]) );
  DFF_X1 sram_wdata_c_reg_94_ ( .D(N453), .CK(clk), .Q(sram_wdata_c[94]) );
  DFF_X1 sram_wdata_c_reg_93_ ( .D(N452), .CK(clk), .Q(sram_wdata_c[93]) );
  DFF_X1 sram_wdata_c_reg_92_ ( .D(N451), .CK(clk), .Q(sram_wdata_c[92]) );
  DFF_X1 sram_wdata_c_reg_91_ ( .D(N450), .CK(clk), .Q(sram_wdata_c[91]) );
  DFF_X1 sram_wdata_c_reg_90_ ( .D(N449), .CK(clk), .Q(sram_wdata_c[90]) );
  DFF_X1 sram_wdata_c_reg_89_ ( .D(N448), .CK(clk), .Q(sram_wdata_c[89]) );
  DFF_X1 sram_wdata_c_reg_88_ ( .D(N447), .CK(clk), .Q(sram_wdata_c[88]) );
  DFF_X1 sram_wdata_c_reg_87_ ( .D(N446), .CK(clk), .Q(sram_wdata_c[87]) );
  DFF_X1 sram_wdata_c_reg_86_ ( .D(N445), .CK(clk), .Q(sram_wdata_c[86]) );
  DFF_X1 sram_wdata_c_reg_85_ ( .D(N444), .CK(clk), .Q(sram_wdata_c[85]) );
  DFF_X1 sram_wdata_c_reg_84_ ( .D(N443), .CK(clk), .Q(sram_wdata_c[84]) );
  DFF_X1 sram_wdata_c_reg_83_ ( .D(N442), .CK(clk), .Q(sram_wdata_c[83]) );
  DFF_X1 sram_wdata_c_reg_82_ ( .D(N441), .CK(clk), .Q(sram_wdata_c[82]) );
  DFF_X1 sram_wdata_c_reg_81_ ( .D(N440), .CK(clk), .Q(sram_wdata_c[81]) );
  DFF_X1 sram_wdata_c_reg_80_ ( .D(N439), .CK(clk), .Q(sram_wdata_c[80]) );
  DFF_X1 sram_wdata_c_reg_79_ ( .D(N438), .CK(clk), .Q(sram_wdata_c[79]) );
  DFF_X1 sram_wdata_c_reg_78_ ( .D(N437), .CK(clk), .Q(sram_wdata_c[78]) );
  DFF_X1 sram_wdata_c_reg_77_ ( .D(N436), .CK(clk), .Q(sram_wdata_c[77]) );
  DFF_X1 sram_wdata_c_reg_76_ ( .D(N435), .CK(clk), .Q(sram_wdata_c[76]) );
  DFF_X1 sram_wdata_c_reg_75_ ( .D(N434), .CK(clk), .Q(sram_wdata_c[75]) );
  DFF_X1 sram_wdata_c_reg_74_ ( .D(N433), .CK(clk), .Q(sram_wdata_c[74]) );
  DFF_X1 sram_wdata_c_reg_73_ ( .D(N432), .CK(clk), .Q(sram_wdata_c[73]) );
  DFF_X1 sram_wdata_c_reg_72_ ( .D(N431), .CK(clk), .Q(sram_wdata_c[72]) );
  DFF_X1 sram_wdata_c_reg_71_ ( .D(N430), .CK(clk), .Q(sram_wdata_c[71]) );
  DFF_X1 sram_wdata_c_reg_70_ ( .D(N429), .CK(clk), .Q(sram_wdata_c[70]) );
  DFF_X1 sram_wdata_c_reg_69_ ( .D(N428), .CK(clk), .Q(sram_wdata_c[69]) );
  DFF_X1 sram_wdata_c_reg_68_ ( .D(N427), .CK(clk), .Q(sram_wdata_c[68]) );
  DFF_X1 sram_wdata_c_reg_67_ ( .D(N426), .CK(clk), .Q(sram_wdata_c[67]) );
  DFF_X1 sram_wdata_c_reg_66_ ( .D(N425), .CK(clk), .Q(sram_wdata_c[66]) );
  DFF_X1 sram_wdata_c_reg_65_ ( .D(N424), .CK(clk), .Q(sram_wdata_c[65]) );
  DFF_X1 sram_wdata_c_reg_64_ ( .D(N423), .CK(clk), .Q(sram_wdata_c[64]) );
  DFF_X1 sram_wdata_c_reg_63_ ( .D(N422), .CK(clk), .Q(sram_wdata_c[63]) );
  DFF_X1 sram_wdata_c_reg_62_ ( .D(N421), .CK(clk), .Q(sram_wdata_c[62]) );
  DFF_X1 sram_wdata_c_reg_61_ ( .D(N420), .CK(clk), .Q(sram_wdata_c[61]) );
  DFF_X1 sram_wdata_c_reg_60_ ( .D(N419), .CK(clk), .Q(sram_wdata_c[60]) );
  DFF_X1 sram_wdata_c_reg_59_ ( .D(N418), .CK(clk), .Q(sram_wdata_c[59]) );
  DFF_X1 sram_wdata_c_reg_58_ ( .D(N417), .CK(clk), .Q(sram_wdata_c[58]) );
  DFF_X1 sram_wdata_c_reg_57_ ( .D(N416), .CK(clk), .Q(sram_wdata_c[57]) );
  DFF_X1 sram_wdata_c_reg_56_ ( .D(N415), .CK(clk), .Q(sram_wdata_c[56]) );
  DFF_X1 sram_wdata_c_reg_55_ ( .D(N414), .CK(clk), .Q(sram_wdata_c[55]) );
  DFF_X1 sram_wdata_c_reg_54_ ( .D(N413), .CK(clk), .Q(sram_wdata_c[54]) );
  DFF_X1 sram_wdata_c_reg_53_ ( .D(N412), .CK(clk), .Q(sram_wdata_c[53]) );
  DFF_X1 sram_wdata_c_reg_52_ ( .D(N411), .CK(clk), .Q(sram_wdata_c[52]) );
  DFF_X1 sram_wdata_c_reg_51_ ( .D(N410), .CK(clk), .Q(sram_wdata_c[51]) );
  DFF_X1 sram_wdata_c_reg_50_ ( .D(N409), .CK(clk), .Q(sram_wdata_c[50]) );
  DFF_X1 sram_wdata_c_reg_49_ ( .D(N408), .CK(clk), .Q(sram_wdata_c[49]) );
  DFF_X1 sram_wdata_c_reg_48_ ( .D(N407), .CK(clk), .Q(sram_wdata_c[48]) );
  DFF_X1 sram_wdata_c_reg_47_ ( .D(N406), .CK(clk), .Q(sram_wdata_c[47]) );
  DFF_X1 sram_wdata_c_reg_46_ ( .D(N405), .CK(clk), .Q(sram_wdata_c[46]) );
  DFF_X1 sram_wdata_c_reg_45_ ( .D(N404), .CK(clk), .Q(sram_wdata_c[45]) );
  DFF_X1 sram_wdata_c_reg_44_ ( .D(N403), .CK(clk), .Q(sram_wdata_c[44]) );
  DFF_X1 sram_wdata_c_reg_43_ ( .D(N402), .CK(clk), .Q(sram_wdata_c[43]) );
  DFF_X1 sram_wdata_c_reg_42_ ( .D(N401), .CK(clk), .Q(sram_wdata_c[42]) );
  DFF_X1 sram_wdata_c_reg_41_ ( .D(N400), .CK(clk), .Q(sram_wdata_c[41]) );
  DFF_X1 sram_wdata_c_reg_40_ ( .D(N399), .CK(clk), .Q(sram_wdata_c[40]) );
  DFF_X1 sram_wdata_c_reg_39_ ( .D(N398), .CK(clk), .Q(sram_wdata_c[39]) );
  DFF_X1 sram_wdata_c_reg_38_ ( .D(N397), .CK(clk), .Q(sram_wdata_c[38]) );
  DFF_X1 sram_wdata_c_reg_37_ ( .D(N396), .CK(clk), .Q(sram_wdata_c[37]) );
  DFF_X1 sram_wdata_c_reg_36_ ( .D(N395), .CK(clk), .Q(sram_wdata_c[36]) );
  DFF_X1 sram_wdata_c_reg_35_ ( .D(N394), .CK(clk), .Q(sram_wdata_c[35]) );
  DFF_X1 sram_wdata_c_reg_34_ ( .D(N393), .CK(clk), .Q(sram_wdata_c[34]) );
  DFF_X1 sram_wdata_c_reg_33_ ( .D(N392), .CK(clk), .Q(sram_wdata_c[33]) );
  DFF_X1 sram_wdata_c_reg_32_ ( .D(N391), .CK(clk), .Q(sram_wdata_c[32]) );
  DFF_X1 sram_wdata_c_reg_31_ ( .D(N390), .CK(clk), .Q(sram_wdata_c[31]) );
  DFF_X1 sram_wdata_c_reg_30_ ( .D(N389), .CK(clk), .Q(sram_wdata_c[30]) );
  DFF_X1 sram_wdata_c_reg_29_ ( .D(N388), .CK(clk), .Q(sram_wdata_c[29]) );
  DFF_X1 sram_wdata_c_reg_28_ ( .D(N387), .CK(clk), .Q(sram_wdata_c[28]) );
  DFF_X1 sram_wdata_c_reg_27_ ( .D(N386), .CK(clk), .Q(sram_wdata_c[27]) );
  DFF_X1 sram_wdata_c_reg_26_ ( .D(N385), .CK(clk), .Q(sram_wdata_c[26]) );
  DFF_X1 sram_wdata_c_reg_25_ ( .D(N384), .CK(clk), .Q(sram_wdata_c[25]) );
  DFF_X1 sram_wdata_c_reg_24_ ( .D(N383), .CK(clk), .Q(sram_wdata_c[24]) );
  DFF_X1 sram_wdata_c_reg_23_ ( .D(N382), .CK(clk), .Q(sram_wdata_c[23]) );
  DFF_X1 sram_wdata_c_reg_22_ ( .D(N381), .CK(clk), .Q(sram_wdata_c[22]) );
  DFF_X1 sram_wdata_c_reg_21_ ( .D(N380), .CK(clk), .Q(sram_wdata_c[21]) );
  DFF_X1 sram_wdata_c_reg_20_ ( .D(N379), .CK(clk), .Q(sram_wdata_c[20]) );
  DFF_X1 sram_wdata_c_reg_19_ ( .D(N378), .CK(clk), .Q(sram_wdata_c[19]) );
  DFF_X1 sram_wdata_c_reg_18_ ( .D(N377), .CK(clk), .Q(sram_wdata_c[18]) );
  DFF_X1 sram_wdata_c_reg_17_ ( .D(N376), .CK(clk), .Q(sram_wdata_c[17]) );
  DFF_X1 sram_wdata_c_reg_16_ ( .D(N375), .CK(clk), .Q(sram_wdata_c[16]) );
  DFF_X1 sram_wdata_c_reg_15_ ( .D(N374), .CK(clk), .Q(sram_wdata_c[15]) );
  DFF_X1 sram_wdata_c_reg_14_ ( .D(N373), .CK(clk), .Q(sram_wdata_c[14]) );
  DFF_X1 sram_wdata_c_reg_13_ ( .D(N372), .CK(clk), .Q(sram_wdata_c[13]) );
  DFF_X1 sram_wdata_c_reg_12_ ( .D(N371), .CK(clk), .Q(sram_wdata_c[12]) );
  DFF_X1 sram_wdata_c_reg_11_ ( .D(N370), .CK(clk), .Q(sram_wdata_c[11]) );
  DFF_X1 sram_wdata_c_reg_10_ ( .D(N369), .CK(clk), .Q(sram_wdata_c[10]) );
  DFF_X1 sram_wdata_c_reg_9_ ( .D(N368), .CK(clk), .Q(sram_wdata_c[9]) );
  DFF_X1 sram_wdata_c_reg_8_ ( .D(N367), .CK(clk), .Q(sram_wdata_c[8]) );
  DFF_X1 sram_wdata_c_reg_7_ ( .D(N366), .CK(clk), .Q(sram_wdata_c[7]) );
  DFF_X1 sram_wdata_c_reg_6_ ( .D(N365), .CK(clk), .Q(sram_wdata_c[6]) );
  DFF_X1 sram_wdata_c_reg_5_ ( .D(N364), .CK(clk), .Q(sram_wdata_c[5]) );
  DFF_X1 sram_wdata_c_reg_4_ ( .D(N363), .CK(clk), .Q(sram_wdata_c[4]) );
  DFF_X1 sram_wdata_c_reg_3_ ( .D(N362), .CK(clk), .Q(sram_wdata_c[3]) );
  DFF_X1 sram_wdata_c_reg_2_ ( .D(N361), .CK(clk), .Q(sram_wdata_c[2]) );
  DFF_X1 sram_wdata_c_reg_1_ ( .D(N360), .CK(clk), .Q(sram_wdata_c[1]) );
  DFF_X1 sram_wdata_c_reg_0_ ( .D(N359), .CK(clk), .Q(sram_wdata_c[0]) );
  DFF_X1 sram_waddr_a_reg_5_ ( .D(N492), .CK(clk), .Q(sram_waddr_a[5]) );
  DFF_X1 sram_waddr_a_reg_4_ ( .D(N491), .CK(clk), .Q(sram_waddr_a[4]) );
  DFF_X1 sram_waddr_a_reg_3_ ( .D(N490), .CK(clk), .Q(sram_waddr_a[3]) );
  DFF_X1 sram_waddr_a_reg_2_ ( .D(N489), .CK(clk), .Q(sram_waddr_a[2]) );
  DFF_X1 sram_waddr_a_reg_1_ ( .D(N488), .CK(clk), .Q(sram_waddr_a[1]) );
  DFF_X1 sram_waddr_a_reg_0_ ( .D(N487), .CK(clk), .Q(sram_waddr_a[0]) );
  XOR2_X1 U3 ( .A(n2701), .B(n3007), .Z(n1) );
  NAND2_X1 U4 ( .A1(n1466), .A2(n1192), .ZN(n2) );
  BUF_X1 U5 ( .A(quantized_data[0]), .Z(n3) );
  BUF_X1 U6 ( .A(quantized_data[1]), .Z(n4) );
  BUF_X1 U7 ( .A(quantized_data[2]), .Z(n5) );
  BUF_X1 U8 ( .A(quantized_data[3]), .Z(n6) );
  BUF_X1 U9 ( .A(quantized_data[4]), .Z(n7) );
  BUF_X1 U10 ( .A(quantized_data[5]), .Z(n8) );
  BUF_X1 U11 ( .A(quantized_data[6]), .Z(n9) );
  BUF_X1 U12 ( .A(quantized_data[7]), .Z(n10) );
  BUF_X1 U13 ( .A(quantized_data[8]), .Z(n11) );
  BUF_X1 U14 ( .A(quantized_data[9]), .Z(n12) );
  BUF_X1 U15 ( .A(quantized_data[10]), .Z(n13) );
  BUF_X1 U16 ( .A(quantized_data[11]), .Z(n14) );
  BUF_X1 U17 ( .A(quantized_data[12]), .Z(n15) );
  BUF_X1 U18 ( .A(quantized_data[13]), .Z(n16) );
  BUF_X1 U19 ( .A(quantized_data[14]), .Z(n17) );
  BUF_X1 U20 ( .A(quantized_data[15]), .Z(n18) );
  BUF_X1 U21 ( .A(quantized_data[32]), .Z(n19) );
  BUF_X1 U22 ( .A(quantized_data[33]), .Z(n20) );
  BUF_X1 U23 ( .A(quantized_data[34]), .Z(n21) );
  BUF_X1 U24 ( .A(quantized_data[35]), .Z(n22) );
  BUF_X1 U25 ( .A(quantized_data[36]), .Z(n23) );
  BUF_X1 U26 ( .A(quantized_data[37]), .Z(n24) );
  BUF_X1 U27 ( .A(quantized_data[38]), .Z(n25) );
  BUF_X1 U28 ( .A(quantized_data[39]), .Z(n26) );
  BUF_X1 U29 ( .A(quantized_data[40]), .Z(n27) );
  BUF_X1 U30 ( .A(quantized_data[41]), .Z(n28) );
  BUF_X1 U31 ( .A(quantized_data[42]), .Z(n29) );
  BUF_X1 U32 ( .A(quantized_data[43]), .Z(n30) );
  BUF_X1 U33 ( .A(quantized_data[44]), .Z(n31) );
  BUF_X1 U34 ( .A(quantized_data[45]), .Z(n32) );
  BUF_X1 U35 ( .A(quantized_data[46]), .Z(n33) );
  BUF_X1 U36 ( .A(quantized_data[47]), .Z(n34) );
  BUF_X1 U37 ( .A(n546), .Z(n35) );
  BUF_X1 U38 ( .A(n87), .Z(n36) );
  INV_X1 U39 ( .A(n36), .ZN(n37) );
  BUF_X1 U40 ( .A(n540), .Z(n38) );
  BUF_X1 U41 ( .A(n15100), .Z(n39) );
  BUF_X1 U42 ( .A(n14900), .Z(n40) );
  BUF_X1 U43 ( .A(n14700), .Z(n41) );
  BUF_X1 U44 ( .A(n14500), .Z(n42) );
  BUF_X1 U45 ( .A(n14300), .Z(n43) );
  BUF_X1 U46 ( .A(n14100), .Z(n44) );
  BUF_X1 U47 ( .A(n13900), .Z(n45) );
  BUF_X1 U48 ( .A(n13700), .Z(n46) );
  BUF_X1 U49 ( .A(n13500), .Z(n47) );
  BUF_X1 U50 ( .A(n13300), .Z(n48) );
  BUF_X1 U51 ( .A(n13100), .Z(n49) );
  BUF_X1 U52 ( .A(n12900), .Z(n50) );
  BUF_X1 U53 ( .A(n12700), .Z(n51) );
  BUF_X1 U54 ( .A(n12500), .Z(n52) );
  BUF_X1 U55 ( .A(n12300), .Z(n53) );
  BUF_X1 U56 ( .A(n12100), .Z(n54) );
  BUF_X1 U57 ( .A(quantized_data[95]), .Z(n55) );
  BUF_X1 U58 ( .A(quantized_data[95]), .Z(n56) );
  BUF_X1 U59 ( .A(quantized_data[94]), .Z(n57) );
  BUF_X1 U60 ( .A(quantized_data[94]), .Z(n58) );
  BUF_X1 U61 ( .A(quantized_data[93]), .Z(n59) );
  BUF_X1 U62 ( .A(quantized_data[93]), .Z(n60) );
  BUF_X1 U63 ( .A(quantized_data[92]), .Z(n61) );
  BUF_X1 U64 ( .A(quantized_data[92]), .Z(n62) );
  BUF_X1 U65 ( .A(quantized_data[91]), .Z(n63) );
  BUF_X1 U66 ( .A(quantized_data[91]), .Z(n64) );
  BUF_X1 U67 ( .A(quantized_data[90]), .Z(n65) );
  BUF_X1 U68 ( .A(quantized_data[90]), .Z(n66) );
  BUF_X1 U69 ( .A(quantized_data[89]), .Z(n67) );
  BUF_X1 U70 ( .A(quantized_data[89]), .Z(n68) );
  BUF_X1 U71 ( .A(quantized_data[88]), .Z(n69) );
  BUF_X1 U72 ( .A(quantized_data[88]), .Z(n70) );
  BUF_X1 U73 ( .A(quantized_data[87]), .Z(n71) );
  BUF_X1 U74 ( .A(quantized_data[87]), .Z(n72) );
  BUF_X1 U75 ( .A(quantized_data[86]), .Z(n73) );
  BUF_X1 U76 ( .A(quantized_data[86]), .Z(n74) );
  BUF_X1 U77 ( .A(quantized_data[85]), .Z(n75) );
  BUF_X1 U78 ( .A(quantized_data[85]), .Z(n76) );
  BUF_X1 U79 ( .A(quantized_data[84]), .Z(n77) );
  BUF_X1 U80 ( .A(quantized_data[84]), .Z(n78) );
  BUF_X1 U81 ( .A(quantized_data[83]), .Z(n79) );
  BUF_X1 U82 ( .A(quantized_data[83]), .Z(n80) );
  BUF_X1 U83 ( .A(quantized_data[82]), .Z(n81) );
  BUF_X1 U84 ( .A(quantized_data[82]), .Z(n82) );
  BUF_X1 U85 ( .A(quantized_data[81]), .Z(n83) );
  BUF_X1 U86 ( .A(quantized_data[81]), .Z(n84) );
  BUF_X1 U87 ( .A(quantized_data[80]), .Z(n85) );
  BUF_X1 U88 ( .A(quantized_data[80]), .Z(n86) );
  BUF_X1 U89 ( .A(matrix_index[3]), .Z(n544) );
  INV_X1 U90 ( .A(n544), .ZN(n87) );
  INV_X1 U91 ( .A(n544), .ZN(n88) );
  INV_X1 U92 ( .A(quantized_data[96]), .ZN(n89) );
  INV_X1 U93 ( .A(quantized_data[97]), .ZN(n90) );
  INV_X1 U94 ( .A(quantized_data[98]), .ZN(n91) );
  INV_X1 U95 ( .A(quantized_data[99]), .ZN(n92) );
  INV_X1 U96 ( .A(quantized_data[100]), .ZN(n93) );
  INV_X1 U97 ( .A(quantized_data[101]), .ZN(n94) );
  INV_X1 U98 ( .A(quantized_data[102]), .ZN(n95) );
  INV_X1 U99 ( .A(quantized_data[103]), .ZN(n96) );
  INV_X1 U100 ( .A(quantized_data[104]), .ZN(n97) );
  INV_X1 U101 ( .A(quantized_data[105]), .ZN(n98) );
  INV_X1 U102 ( .A(quantized_data[106]), .ZN(n99) );
  INV_X1 U103 ( .A(quantized_data[107]), .ZN(n10000) );
  INV_X1 U104 ( .A(quantized_data[108]), .ZN(n10100) );
  INV_X1 U105 ( .A(quantized_data[109]), .ZN(n10200) );
  INV_X1 U106 ( .A(quantized_data[110]), .ZN(n10300) );
  INV_X1 U107 ( .A(quantized_data[111]), .ZN(n10400) );
  INV_X1 U108 ( .A(quantized_data[112]), .ZN(n10500) );
  INV_X1 U109 ( .A(quantized_data[113]), .ZN(n10600) );
  INV_X1 U110 ( .A(quantized_data[114]), .ZN(n10700) );
  INV_X1 U111 ( .A(quantized_data[115]), .ZN(n10800) );
  INV_X1 U112 ( .A(quantized_data[116]), .ZN(n10900) );
  INV_X1 U113 ( .A(quantized_data[117]), .ZN(n11000) );
  INV_X1 U114 ( .A(quantized_data[118]), .ZN(n11100) );
  INV_X1 U115 ( .A(quantized_data[119]), .ZN(n11200) );
  INV_X1 U116 ( .A(quantized_data[120]), .ZN(n11300) );
  INV_X1 U117 ( .A(quantized_data[121]), .ZN(n11400) );
  INV_X1 U118 ( .A(quantized_data[122]), .ZN(n11500) );
  INV_X1 U119 ( .A(quantized_data[123]), .ZN(n11600) );
  INV_X1 U120 ( .A(quantized_data[124]), .ZN(n11700) );
  INV_X1 U121 ( .A(quantized_data[125]), .ZN(n11800) );
  INV_X1 U122 ( .A(quantized_data[126]), .ZN(n11900) );
  INV_X1 U123 ( .A(quantized_data[127]), .ZN(n12000) );
  BUF_X1 U124 ( .A(quantized_data[31]), .Z(n12100) );
  BUF_X1 U125 ( .A(quantized_data[31]), .Z(n12200) );
  BUF_X1 U126 ( .A(quantized_data[30]), .Z(n12300) );
  BUF_X1 U127 ( .A(quantized_data[30]), .Z(n12400) );
  BUF_X1 U128 ( .A(quantized_data[29]), .Z(n12500) );
  BUF_X1 U129 ( .A(quantized_data[29]), .Z(n12600) );
  BUF_X1 U130 ( .A(quantized_data[28]), .Z(n12700) );
  BUF_X1 U131 ( .A(quantized_data[28]), .Z(n12800) );
  BUF_X1 U132 ( .A(quantized_data[27]), .Z(n12900) );
  BUF_X1 U133 ( .A(quantized_data[27]), .Z(n13000) );
  BUF_X1 U134 ( .A(quantized_data[26]), .Z(n13100) );
  BUF_X1 U135 ( .A(quantized_data[26]), .Z(n13200) );
  BUF_X1 U136 ( .A(quantized_data[25]), .Z(n13300) );
  BUF_X1 U137 ( .A(quantized_data[25]), .Z(n13400) );
  BUF_X1 U138 ( .A(quantized_data[24]), .Z(n13500) );
  BUF_X1 U139 ( .A(quantized_data[24]), .Z(n13600) );
  BUF_X1 U140 ( .A(quantized_data[23]), .Z(n13700) );
  BUF_X1 U141 ( .A(quantized_data[23]), .Z(n13800) );
  BUF_X1 U142 ( .A(quantized_data[22]), .Z(n13900) );
  BUF_X1 U143 ( .A(quantized_data[22]), .Z(n14000) );
  BUF_X1 U144 ( .A(quantized_data[21]), .Z(n14100) );
  BUF_X1 U145 ( .A(quantized_data[21]), .Z(n14200) );
  BUF_X1 U146 ( .A(quantized_data[20]), .Z(n14300) );
  BUF_X1 U147 ( .A(quantized_data[20]), .Z(n14400) );
  BUF_X1 U148 ( .A(quantized_data[19]), .Z(n14500) );
  BUF_X1 U149 ( .A(quantized_data[19]), .Z(n14600) );
  BUF_X1 U150 ( .A(quantized_data[18]), .Z(n14700) );
  BUF_X1 U151 ( .A(quantized_data[18]), .Z(n14800) );
  BUF_X1 U152 ( .A(quantized_data[17]), .Z(n14900) );
  BUF_X1 U153 ( .A(quantized_data[17]), .Z(n15000) );
  BUF_X1 U154 ( .A(quantized_data[16]), .Z(n15100) );
  BUF_X1 U155 ( .A(quantized_data[16]), .Z(n15200) );
  INV_X1 U156 ( .A(matrix_index[5]), .ZN(n15300) );
  INV_X1 U157 ( .A(n15300), .ZN(n15400) );
  INV_X1 U158 ( .A(n15300), .ZN(n15510) );
  INV_X1 U159 ( .A(quantized_data[79]), .ZN(n15630) );
  INV_X1 U160 ( .A(n15630), .ZN(n15700) );
  INV_X1 U161 ( .A(n15630), .ZN(n15800) );
  INV_X1 U162 ( .A(n1469), .ZN(n15970) );
  INV_X1 U163 ( .A(quantized_data[78]), .ZN(n16000) );
  INV_X1 U164 ( .A(n16000), .ZN(n16100) );
  INV_X1 U165 ( .A(n16000), .ZN(n16200) );
  INV_X1 U166 ( .A(n1462), .ZN(n16390) );
  INV_X1 U167 ( .A(quantized_data[77]), .ZN(n16400) );
  INV_X1 U168 ( .A(n16400), .ZN(n16500) );
  INV_X1 U169 ( .A(n16400), .ZN(n16600) );
  INV_X1 U170 ( .A(n1455), .ZN(n16700) );
  INV_X1 U171 ( .A(quantized_data[76]), .ZN(n16800) );
  INV_X1 U172 ( .A(n16800), .ZN(n16900) );
  INV_X1 U173 ( .A(n16800), .ZN(n17000) );
  INV_X1 U174 ( .A(n1448), .ZN(n17100) );
  INV_X1 U175 ( .A(quantized_data[75]), .ZN(n17200) );
  INV_X1 U176 ( .A(n17200), .ZN(n17300) );
  INV_X1 U177 ( .A(n17200), .ZN(n17400) );
  INV_X1 U178 ( .A(n1443), .ZN(n17500) );
  INV_X1 U179 ( .A(quantized_data[74]), .ZN(n17600) );
  INV_X1 U180 ( .A(n17600), .ZN(n17700) );
  INV_X1 U181 ( .A(n17600), .ZN(n17800) );
  INV_X1 U182 ( .A(n1436), .ZN(n17900) );
  INV_X1 U183 ( .A(quantized_data[73]), .ZN(n18000) );
  INV_X1 U184 ( .A(n18000), .ZN(n18100) );
  INV_X1 U185 ( .A(n18000), .ZN(n18200) );
  INV_X1 U186 ( .A(n1429), .ZN(n18300) );
  INV_X1 U187 ( .A(quantized_data[72]), .ZN(n18400) );
  INV_X1 U188 ( .A(n18400), .ZN(n18500) );
  INV_X1 U189 ( .A(n18400), .ZN(n18600) );
  INV_X1 U190 ( .A(n1422), .ZN(n18700) );
  INV_X1 U191 ( .A(quantized_data[71]), .ZN(n18800) );
  INV_X1 U192 ( .A(n18800), .ZN(n18900) );
  INV_X1 U193 ( .A(n18800), .ZN(n19000) );
  INV_X1 U194 ( .A(n1417), .ZN(n19100) );
  INV_X1 U195 ( .A(quantized_data[70]), .ZN(n19200) );
  INV_X1 U196 ( .A(n19200), .ZN(n19300) );
  INV_X1 U197 ( .A(n19200), .ZN(n19400) );
  INV_X1 U198 ( .A(n14101), .ZN(n19500) );
  INV_X1 U199 ( .A(quantized_data[69]), .ZN(n19600) );
  INV_X1 U200 ( .A(n19600), .ZN(n19700) );
  INV_X1 U201 ( .A(n19600), .ZN(n19800) );
  INV_X1 U202 ( .A(n1405), .ZN(n19900) );
  INV_X1 U203 ( .A(quantized_data[68]), .ZN(n20000) );
  INV_X1 U204 ( .A(n20000), .ZN(n20100) );
  INV_X1 U205 ( .A(n20000), .ZN(n20200) );
  INV_X1 U206 ( .A(n14001), .ZN(n20300) );
  INV_X1 U207 ( .A(quantized_data[67]), .ZN(n20400) );
  INV_X1 U208 ( .A(n20400), .ZN(n20500) );
  INV_X1 U209 ( .A(n20400), .ZN(n20600) );
  INV_X1 U210 ( .A(n1395), .ZN(n20700) );
  INV_X1 U211 ( .A(quantized_data[66]), .ZN(n20800) );
  INV_X1 U212 ( .A(n20800), .ZN(n20900) );
  INV_X1 U213 ( .A(n20800), .ZN(n21000) );
  INV_X1 U214 ( .A(n1388), .ZN(n21100) );
  INV_X1 U215 ( .A(quantized_data[65]), .ZN(n21200) );
  INV_X1 U216 ( .A(n21200), .ZN(n21300) );
  INV_X1 U217 ( .A(n21200), .ZN(n21400) );
  INV_X1 U218 ( .A(n1381), .ZN(n21500) );
  INV_X1 U219 ( .A(quantized_data[64]), .ZN(n21600) );
  INV_X1 U220 ( .A(n21600), .ZN(n21700) );
  INV_X1 U221 ( .A(n21600), .ZN(n21800) );
  INV_X1 U222 ( .A(n1374), .ZN(n21900) );
  INV_X1 U223 ( .A(quantized_data[47]), .ZN(n22000) );
  INV_X1 U224 ( .A(n22000), .ZN(n22100) );
  INV_X1 U225 ( .A(n22000), .ZN(n22200) );
  INV_X1 U226 ( .A(quantized_data[46]), .ZN(n22300) );
  INV_X1 U227 ( .A(n22300), .ZN(n22400) );
  INV_X1 U228 ( .A(n22300), .ZN(n22500) );
  INV_X1 U229 ( .A(quantized_data[45]), .ZN(n22600) );
  INV_X1 U230 ( .A(n22600), .ZN(n22700) );
  INV_X1 U231 ( .A(n22600), .ZN(n22800) );
  INV_X1 U232 ( .A(quantized_data[44]), .ZN(n22900) );
  INV_X1 U233 ( .A(n22900), .ZN(n23000) );
  INV_X1 U234 ( .A(n22900), .ZN(n23100) );
  INV_X1 U235 ( .A(quantized_data[43]), .ZN(n23200) );
  INV_X1 U236 ( .A(n23200), .ZN(n23300) );
  INV_X1 U237 ( .A(n23200), .ZN(n23400) );
  INV_X1 U238 ( .A(quantized_data[42]), .ZN(n23500) );
  INV_X1 U239 ( .A(n23500), .ZN(n23600) );
  INV_X1 U240 ( .A(n23500), .ZN(n23700) );
  INV_X1 U241 ( .A(quantized_data[41]), .ZN(n23800) );
  INV_X1 U242 ( .A(n23800), .ZN(n23900) );
  INV_X1 U243 ( .A(n23800), .ZN(n24000) );
  INV_X1 U244 ( .A(quantized_data[40]), .ZN(n24100) );
  INV_X1 U245 ( .A(n24100), .ZN(n24200) );
  INV_X1 U246 ( .A(n24100), .ZN(n24300) );
  INV_X1 U247 ( .A(quantized_data[39]), .ZN(n24400) );
  INV_X1 U248 ( .A(n24400), .ZN(n24500) );
  INV_X1 U249 ( .A(n24400), .ZN(n24600) );
  INV_X1 U250 ( .A(quantized_data[38]), .ZN(n24700) );
  INV_X1 U251 ( .A(n24700), .ZN(n24800) );
  INV_X1 U252 ( .A(n24700), .ZN(n24900) );
  INV_X1 U253 ( .A(quantized_data[37]), .ZN(n25000) );
  INV_X1 U254 ( .A(n25000), .ZN(n25100) );
  INV_X1 U255 ( .A(n25000), .ZN(n25200) );
  INV_X1 U256 ( .A(quantized_data[36]), .ZN(n25300) );
  INV_X1 U257 ( .A(n25300), .ZN(n25400) );
  INV_X1 U258 ( .A(n25300), .ZN(n25500) );
  INV_X1 U259 ( .A(quantized_data[35]), .ZN(n25600) );
  INV_X1 U260 ( .A(n25600), .ZN(n25700) );
  INV_X1 U261 ( .A(n25600), .ZN(n25800) );
  INV_X1 U262 ( .A(quantized_data[34]), .ZN(n25900) );
  INV_X1 U263 ( .A(n25900), .ZN(n26000) );
  INV_X1 U264 ( .A(n25900), .ZN(n26100) );
  INV_X1 U265 ( .A(quantized_data[33]), .ZN(n26200) );
  INV_X1 U266 ( .A(n26200), .ZN(n26300) );
  INV_X1 U267 ( .A(n26200), .ZN(n26400) );
  INV_X1 U268 ( .A(quantized_data[32]), .ZN(n26500) );
  INV_X1 U269 ( .A(n26500), .ZN(n26600) );
  INV_X1 U270 ( .A(n26500), .ZN(n26700) );
  INV_X1 U271 ( .A(quantized_data[15]), .ZN(n26800) );
  INV_X1 U272 ( .A(n26800), .ZN(n26900) );
  INV_X1 U273 ( .A(n26800), .ZN(n27000) );
  INV_X1 U274 ( .A(quantized_data[14]), .ZN(n27100) );
  INV_X1 U275 ( .A(n27100), .ZN(n27200) );
  INV_X1 U276 ( .A(n27100), .ZN(n27300) );
  INV_X1 U277 ( .A(quantized_data[13]), .ZN(n27400) );
  INV_X1 U278 ( .A(n27400), .ZN(n27500) );
  INV_X1 U279 ( .A(n27400), .ZN(n27600) );
  INV_X1 U280 ( .A(quantized_data[12]), .ZN(n27700) );
  INV_X1 U281 ( .A(n27700), .ZN(n27800) );
  INV_X1 U282 ( .A(n27700), .ZN(n27900) );
  INV_X1 U283 ( .A(quantized_data[11]), .ZN(n28000) );
  INV_X1 U284 ( .A(n28000), .ZN(n28100) );
  INV_X1 U285 ( .A(n28000), .ZN(n28200) );
  INV_X1 U286 ( .A(quantized_data[10]), .ZN(n28300) );
  INV_X1 U287 ( .A(n28300), .ZN(n28400) );
  INV_X1 U288 ( .A(n28300), .ZN(n28500) );
  INV_X1 U289 ( .A(quantized_data[9]), .ZN(n28600) );
  INV_X1 U290 ( .A(n28600), .ZN(n28700) );
  INV_X1 U291 ( .A(n28600), .ZN(n28800) );
  INV_X1 U292 ( .A(quantized_data[8]), .ZN(n28900) );
  INV_X1 U293 ( .A(n28900), .ZN(n29000) );
  INV_X1 U294 ( .A(n28900), .ZN(n29100) );
  INV_X1 U295 ( .A(quantized_data[7]), .ZN(n29200) );
  INV_X1 U296 ( .A(n29200), .ZN(n29300) );
  INV_X1 U297 ( .A(n29200), .ZN(n29400) );
  INV_X1 U298 ( .A(quantized_data[6]), .ZN(n29500) );
  INV_X1 U299 ( .A(n29500), .ZN(n29600) );
  INV_X1 U300 ( .A(n29500), .ZN(n29700) );
  INV_X1 U301 ( .A(quantized_data[5]), .ZN(n29800) );
  INV_X1 U302 ( .A(n29800), .ZN(n29900) );
  INV_X1 U303 ( .A(n29800), .ZN(n30000) );
  INV_X1 U304 ( .A(quantized_data[4]), .ZN(n30100) );
  INV_X1 U305 ( .A(n30100), .ZN(n30200) );
  INV_X1 U306 ( .A(n30100), .ZN(n30300) );
  INV_X1 U307 ( .A(quantized_data[3]), .ZN(n30400) );
  INV_X1 U308 ( .A(n30400), .ZN(n30500) );
  INV_X1 U309 ( .A(n30400), .ZN(n30600) );
  INV_X1 U310 ( .A(quantized_data[2]), .ZN(n30700) );
  INV_X1 U311 ( .A(n30700), .ZN(n30800) );
  INV_X1 U312 ( .A(n30700), .ZN(n30900) );
  INV_X1 U313 ( .A(quantized_data[1]), .ZN(n31000) );
  INV_X1 U314 ( .A(n31000), .ZN(n31100) );
  INV_X1 U315 ( .A(n31000), .ZN(n31200) );
  INV_X1 U316 ( .A(quantized_data[0]), .ZN(n31300) );
  INV_X1 U317 ( .A(n31300), .ZN(n31400) );
  INV_X1 U318 ( .A(n31300), .ZN(n31500) );
  INV_X1 U319 ( .A(quantized_data[63]), .ZN(n31600) );
  INV_X1 U320 ( .A(n31600), .ZN(n31700) );
  INV_X1 U321 ( .A(n31600), .ZN(n31800) );
  INV_X1 U322 ( .A(n1182), .ZN(n31900) );
  INV_X1 U323 ( .A(quantized_data[62]), .ZN(n32000) );
  INV_X1 U324 ( .A(n32000), .ZN(n32100) );
  INV_X1 U325 ( .A(n32000), .ZN(n32200) );
  INV_X1 U326 ( .A(n1185), .ZN(n32300) );
  INV_X1 U327 ( .A(quantized_data[61]), .ZN(n32400) );
  INV_X1 U328 ( .A(n32400), .ZN(n32500) );
  INV_X1 U329 ( .A(n32400), .ZN(n32600) );
  INV_X1 U330 ( .A(n1176), .ZN(n32700) );
  INV_X1 U331 ( .A(quantized_data[60]), .ZN(n32800) );
  INV_X1 U332 ( .A(n32800), .ZN(n32900) );
  INV_X1 U333 ( .A(n32800), .ZN(n33000) );
  INV_X1 U334 ( .A(n1179), .ZN(n33100) );
  INV_X1 U335 ( .A(quantized_data[59]), .ZN(n33200) );
  INV_X1 U336 ( .A(n33200), .ZN(n33300) );
  INV_X1 U337 ( .A(n33200), .ZN(n33400) );
  INV_X1 U338 ( .A(n11701), .ZN(n33500) );
  INV_X1 U339 ( .A(quantized_data[58]), .ZN(n33600) );
  INV_X1 U340 ( .A(n33600), .ZN(n33700) );
  INV_X1 U341 ( .A(n33600), .ZN(n33800) );
  INV_X1 U342 ( .A(n1173), .ZN(n33900) );
  INV_X1 U343 ( .A(quantized_data[57]), .ZN(n34000) );
  INV_X1 U344 ( .A(n34000), .ZN(n34100) );
  INV_X1 U345 ( .A(n34000), .ZN(n34200) );
  INV_X1 U346 ( .A(n1164), .ZN(n34300) );
  INV_X1 U347 ( .A(quantized_data[56]), .ZN(n34400) );
  INV_X1 U348 ( .A(n34400), .ZN(n34500) );
  INV_X1 U349 ( .A(n34400), .ZN(n34600) );
  INV_X1 U350 ( .A(n1167), .ZN(n34700) );
  INV_X1 U351 ( .A(quantized_data[55]), .ZN(n34800) );
  INV_X1 U352 ( .A(n34800), .ZN(n34900) );
  INV_X1 U353 ( .A(n34800), .ZN(n35000) );
  INV_X1 U354 ( .A(n1158), .ZN(n35100) );
  INV_X1 U355 ( .A(quantized_data[54]), .ZN(n35200) );
  INV_X1 U356 ( .A(n35200), .ZN(n35300) );
  INV_X1 U357 ( .A(n35200), .ZN(n35400) );
  INV_X1 U358 ( .A(n1161), .ZN(n35500) );
  INV_X1 U359 ( .A(quantized_data[53]), .ZN(n35600) );
  INV_X1 U360 ( .A(n35600), .ZN(n35700) );
  INV_X1 U361 ( .A(n35600), .ZN(n35800) );
  INV_X1 U362 ( .A(n1152), .ZN(n35900) );
  INV_X1 U363 ( .A(quantized_data[52]), .ZN(n36000) );
  INV_X1 U364 ( .A(n36000), .ZN(n36100) );
  INV_X1 U365 ( .A(n36000), .ZN(n36200) );
  INV_X1 U366 ( .A(n1155), .ZN(n36300) );
  INV_X1 U367 ( .A(quantized_data[51]), .ZN(n36400) );
  INV_X1 U368 ( .A(n36400), .ZN(n36500) );
  INV_X1 U369 ( .A(n36400), .ZN(n36600) );
  INV_X1 U370 ( .A(n1146), .ZN(n36700) );
  INV_X1 U371 ( .A(quantized_data[50]), .ZN(n36800) );
  INV_X1 U372 ( .A(n36800), .ZN(n36900) );
  INV_X1 U373 ( .A(n36800), .ZN(n37000) );
  INV_X1 U374 ( .A(n1149), .ZN(n37100) );
  INV_X1 U375 ( .A(quantized_data[49]), .ZN(n37200) );
  INV_X1 U376 ( .A(n37200), .ZN(n37300) );
  INV_X1 U377 ( .A(n37200), .ZN(n37400) );
  INV_X1 U378 ( .A(n11401), .ZN(n37500) );
  INV_X1 U379 ( .A(quantized_data[48]), .ZN(n37600) );
  INV_X1 U380 ( .A(n37600), .ZN(n37700) );
  INV_X1 U381 ( .A(n37600), .ZN(n37800) );
  INV_X1 U382 ( .A(n1143), .ZN(n37900) );
  INV_X1 U383 ( .A(quantized_data[127]), .ZN(n38000) );
  INV_X1 U384 ( .A(n38000), .ZN(n38100) );
  INV_X1 U385 ( .A(n12000), .ZN(n38200) );
  INV_X1 U386 ( .A(n38000), .ZN(n38300) );
  INV_X1 U387 ( .A(n12000), .ZN(n38400) );
  INV_X1 U388 ( .A(quantized_data[126]), .ZN(n38500) );
  INV_X1 U389 ( .A(n38500), .ZN(n38600) );
  INV_X1 U390 ( .A(n11900), .ZN(n38700) );
  INV_X1 U391 ( .A(n38500), .ZN(n38800) );
  INV_X1 U392 ( .A(n11900), .ZN(n38900) );
  INV_X1 U393 ( .A(quantized_data[125]), .ZN(n39000) );
  INV_X1 U394 ( .A(n39000), .ZN(n39100) );
  INV_X1 U395 ( .A(n11800), .ZN(n39200) );
  INV_X1 U396 ( .A(n39000), .ZN(n39300) );
  INV_X1 U397 ( .A(n11800), .ZN(n39400) );
  INV_X1 U398 ( .A(quantized_data[124]), .ZN(n39500) );
  INV_X1 U399 ( .A(n39500), .ZN(n39600) );
  INV_X1 U400 ( .A(n11700), .ZN(n39700) );
  INV_X1 U401 ( .A(n39500), .ZN(n39800) );
  INV_X1 U402 ( .A(n11700), .ZN(n39900) );
  INV_X1 U403 ( .A(quantized_data[123]), .ZN(n40000) );
  INV_X1 U404 ( .A(n40000), .ZN(n40100) );
  INV_X1 U405 ( .A(n11600), .ZN(n40200) );
  INV_X1 U406 ( .A(n40000), .ZN(n40300) );
  INV_X1 U407 ( .A(n11600), .ZN(n40400) );
  INV_X1 U408 ( .A(quantized_data[122]), .ZN(n40500) );
  INV_X1 U409 ( .A(n40500), .ZN(n40600) );
  INV_X1 U410 ( .A(n11500), .ZN(n40700) );
  INV_X1 U411 ( .A(n40500), .ZN(n40800) );
  INV_X1 U412 ( .A(n11500), .ZN(n40900) );
  INV_X1 U413 ( .A(quantized_data[121]), .ZN(n41000) );
  INV_X1 U414 ( .A(n41000), .ZN(n41100) );
  INV_X1 U415 ( .A(n11400), .ZN(n41200) );
  INV_X1 U416 ( .A(n41000), .ZN(n41300) );
  INV_X1 U417 ( .A(n11400), .ZN(n41400) );
  INV_X1 U418 ( .A(quantized_data[120]), .ZN(n41500) );
  INV_X1 U419 ( .A(n41500), .ZN(n41600) );
  INV_X1 U420 ( .A(n11300), .ZN(n41700) );
  INV_X1 U421 ( .A(n41500), .ZN(n41800) );
  INV_X1 U422 ( .A(n11300), .ZN(n41900) );
  INV_X1 U423 ( .A(quantized_data[119]), .ZN(n42000) );
  INV_X1 U424 ( .A(n42000), .ZN(n42100) );
  INV_X1 U425 ( .A(n11200), .ZN(n42200) );
  INV_X1 U426 ( .A(n42000), .ZN(n42300) );
  INV_X1 U427 ( .A(n11200), .ZN(n42400) );
  INV_X1 U428 ( .A(quantized_data[118]), .ZN(n42500) );
  INV_X1 U429 ( .A(n42500), .ZN(n42600) );
  INV_X1 U430 ( .A(n11100), .ZN(n42700) );
  INV_X1 U431 ( .A(n42500), .ZN(n42800) );
  INV_X1 U432 ( .A(n11100), .ZN(n42900) );
  INV_X1 U433 ( .A(quantized_data[117]), .ZN(n43000) );
  INV_X1 U434 ( .A(n43000), .ZN(n43100) );
  INV_X1 U435 ( .A(n11000), .ZN(n43200) );
  INV_X1 U436 ( .A(n43000), .ZN(n43300) );
  INV_X1 U437 ( .A(n11000), .ZN(n43400) );
  INV_X1 U438 ( .A(quantized_data[116]), .ZN(n43500) );
  INV_X1 U439 ( .A(n43500), .ZN(n43600) );
  INV_X1 U440 ( .A(n10900), .ZN(n43700) );
  INV_X1 U441 ( .A(n43500), .ZN(n43800) );
  INV_X1 U442 ( .A(n10900), .ZN(n43900) );
  INV_X1 U443 ( .A(quantized_data[115]), .ZN(n44000) );
  INV_X1 U444 ( .A(n44000), .ZN(n44100) );
  INV_X1 U445 ( .A(n10800), .ZN(n44200) );
  INV_X1 U446 ( .A(n44000), .ZN(n44300) );
  INV_X1 U447 ( .A(n10800), .ZN(n44400) );
  INV_X1 U448 ( .A(quantized_data[114]), .ZN(n44500) );
  INV_X1 U449 ( .A(n44500), .ZN(n44600) );
  INV_X1 U450 ( .A(n10700), .ZN(n44700) );
  INV_X1 U451 ( .A(n44500), .ZN(n44800) );
  INV_X1 U452 ( .A(n10700), .ZN(n44900) );
  INV_X1 U453 ( .A(quantized_data[113]), .ZN(n45000) );
  INV_X1 U454 ( .A(n45000), .ZN(n45100) );
  INV_X1 U455 ( .A(n10600), .ZN(n45200) );
  INV_X1 U456 ( .A(n45000), .ZN(n45300) );
  INV_X1 U457 ( .A(n10600), .ZN(n45400) );
  INV_X1 U458 ( .A(quantized_data[112]), .ZN(n45500) );
  INV_X1 U459 ( .A(n45500), .ZN(n45600) );
  INV_X1 U460 ( .A(n10500), .ZN(n45700) );
  INV_X1 U461 ( .A(n45500), .ZN(n45800) );
  INV_X1 U462 ( .A(n10500), .ZN(n45900) );
  INV_X1 U463 ( .A(quantized_data[111]), .ZN(n46000) );
  INV_X1 U464 ( .A(n46000), .ZN(n46100) );
  INV_X1 U465 ( .A(n10400), .ZN(n46200) );
  INV_X1 U466 ( .A(n10400), .ZN(n46300) );
  INV_X1 U467 ( .A(n46000), .ZN(n46400) );
  INV_X1 U468 ( .A(quantized_data[110]), .ZN(n46500) );
  INV_X1 U469 ( .A(n46500), .ZN(n46600) );
  INV_X1 U470 ( .A(n10300), .ZN(n46700) );
  INV_X1 U471 ( .A(n46500), .ZN(n46800) );
  INV_X1 U472 ( .A(n10300), .ZN(n46900) );
  INV_X1 U473 ( .A(quantized_data[109]), .ZN(n4700) );
  INV_X1 U474 ( .A(n4700), .ZN(n4710) );
  INV_X1 U475 ( .A(n10200), .ZN(n4720) );
  INV_X1 U476 ( .A(n4700), .ZN(n4730) );
  INV_X1 U477 ( .A(n10200), .ZN(n4740) );
  INV_X1 U478 ( .A(quantized_data[108]), .ZN(n4750) );
  INV_X1 U479 ( .A(n4750), .ZN(n4760) );
  INV_X1 U480 ( .A(n10100), .ZN(n4770) );
  INV_X1 U481 ( .A(n4750), .ZN(n4780) );
  INV_X1 U482 ( .A(n10100), .ZN(n4790) );
  INV_X1 U483 ( .A(quantized_data[107]), .ZN(n4800) );
  INV_X1 U484 ( .A(n4800), .ZN(n4810) );
  INV_X1 U485 ( .A(n10000), .ZN(n4820) );
  INV_X1 U486 ( .A(n4800), .ZN(n4830) );
  INV_X1 U487 ( .A(n10000), .ZN(n4840) );
  INV_X1 U488 ( .A(quantized_data[106]), .ZN(n4850) );
  INV_X1 U489 ( .A(n4850), .ZN(n4860) );
  INV_X1 U490 ( .A(n99), .ZN(n4870) );
  INV_X1 U491 ( .A(n4850), .ZN(n4880) );
  INV_X1 U492 ( .A(n99), .ZN(n4890) );
  INV_X1 U493 ( .A(quantized_data[105]), .ZN(n4900) );
  INV_X1 U494 ( .A(n4900), .ZN(n4910) );
  INV_X1 U495 ( .A(n98), .ZN(n4920) );
  INV_X1 U496 ( .A(n4900), .ZN(n493) );
  INV_X1 U497 ( .A(n98), .ZN(n494) );
  INV_X1 U498 ( .A(quantized_data[104]), .ZN(n495) );
  INV_X1 U499 ( .A(n495), .ZN(n496) );
  INV_X1 U500 ( .A(n97), .ZN(n497) );
  INV_X1 U501 ( .A(n495), .ZN(n498) );
  INV_X1 U502 ( .A(n97), .ZN(n4990) );
  INV_X1 U503 ( .A(quantized_data[103]), .ZN(n5000) );
  INV_X1 U504 ( .A(n5000), .ZN(n5010) );
  INV_X1 U505 ( .A(n96), .ZN(n5020) );
  INV_X1 U506 ( .A(n5000), .ZN(n5030) );
  INV_X1 U507 ( .A(n96), .ZN(n5040) );
  INV_X1 U508 ( .A(quantized_data[102]), .ZN(n505) );
  INV_X1 U509 ( .A(n505), .ZN(n506) );
  INV_X1 U510 ( .A(n95), .ZN(n507) );
  INV_X1 U511 ( .A(n505), .ZN(n508) );
  INV_X1 U512 ( .A(n95), .ZN(n509) );
  INV_X1 U513 ( .A(quantized_data[101]), .ZN(n510) );
  INV_X1 U514 ( .A(n510), .ZN(n511) );
  INV_X1 U515 ( .A(n94), .ZN(n512) );
  INV_X1 U516 ( .A(n510), .ZN(n513) );
  INV_X1 U517 ( .A(n94), .ZN(n514) );
  INV_X1 U518 ( .A(quantized_data[100]), .ZN(n515) );
  INV_X1 U519 ( .A(n515), .ZN(n516) );
  INV_X1 U520 ( .A(n93), .ZN(n517) );
  INV_X1 U521 ( .A(n515), .ZN(n518) );
  INV_X1 U522 ( .A(n93), .ZN(n519) );
  INV_X1 U523 ( .A(quantized_data[99]), .ZN(n520) );
  INV_X1 U524 ( .A(n520), .ZN(n521) );
  INV_X1 U525 ( .A(n92), .ZN(n522) );
  INV_X1 U526 ( .A(n520), .ZN(n523) );
  INV_X1 U527 ( .A(n92), .ZN(n524) );
  INV_X1 U528 ( .A(quantized_data[98]), .ZN(n525) );
  INV_X1 U529 ( .A(n525), .ZN(n526) );
  INV_X1 U530 ( .A(n91), .ZN(n527) );
  INV_X1 U531 ( .A(n525), .ZN(n528) );
  INV_X1 U532 ( .A(n91), .ZN(n529) );
  INV_X1 U533 ( .A(quantized_data[97]), .ZN(n530) );
  INV_X1 U534 ( .A(n530), .ZN(n531) );
  INV_X1 U535 ( .A(n90), .ZN(n532) );
  INV_X1 U536 ( .A(n530), .ZN(n533) );
  INV_X1 U537 ( .A(n90), .ZN(n534) );
  INV_X1 U538 ( .A(quantized_data[96]), .ZN(n535) );
  INV_X1 U539 ( .A(n535), .ZN(n536) );
  INV_X1 U540 ( .A(n89), .ZN(n537) );
  INV_X1 U541 ( .A(n535), .ZN(n538) );
  INV_X1 U542 ( .A(n89), .ZN(n539) );
  INV_X1 U543 ( .A(matrix_index[4]), .ZN(n540) );
  INV_X1 U544 ( .A(n540), .ZN(n541) );
  INV_X1 U545 ( .A(n38), .ZN(n542) );
  INV_X1 U546 ( .A(n38), .ZN(n543) );
  INV_X1 U547 ( .A(n87), .ZN(n545) );
  INV_X1 U548 ( .A(n88), .ZN(n546) );
  INV_X1 U549 ( .A(n36), .ZN(n547) );
  INV_X1 U550 ( .A(n88), .ZN(n548) );
  CLKBUF_X1 U551 ( .A(n3167), .Z(n549) );
  CLKBUF_X1 U552 ( .A(n3426), .Z(n550) );
  CLKBUF_X1 U553 ( .A(n37101), .Z(n551) );
  CLKBUF_X1 U554 ( .A(n37101), .Z(n552) );
  CLKBUF_X1 U555 ( .A(n4188), .Z(n553) );
  CLKBUF_X1 U556 ( .A(n4187), .Z(n554) );
  CLKBUF_X1 U557 ( .A(n4673), .Z(n555) );
  CLKBUF_X1 U558 ( .A(n1745), .Z(n556) );
  CLKBUF_X1 U559 ( .A(n3402), .Z(n557) );
  CLKBUF_X1 U560 ( .A(n909), .Z(n558) );
  CLKBUF_X1 U561 ( .A(n1196), .Z(n559) );
  CLKBUF_X1 U562 ( .A(n3836), .Z(n560) );
  CLKBUF_X1 U563 ( .A(n3838), .Z(n561) );
  CLKBUF_X1 U564 ( .A(n38401), .Z(n562) );
  CLKBUF_X1 U565 ( .A(n3833), .Z(n563) );
  CLKBUF_X1 U566 ( .A(n3844), .Z(n564) );
  CLKBUF_X1 U567 ( .A(n3846), .Z(n565) );
  CLKBUF_X1 U568 ( .A(n3848), .Z(n566) );
  CLKBUF_X1 U569 ( .A(n3842), .Z(n567) );
  CLKBUF_X1 U570 ( .A(n3852), .Z(n568) );
  CLKBUF_X1 U571 ( .A(n3854), .Z(n569) );
  CLKBUF_X1 U572 ( .A(n3856), .Z(n570) );
  CLKBUF_X1 U573 ( .A(n38501), .Z(n571) );
  CLKBUF_X1 U574 ( .A(n38601), .Z(n572) );
  CLKBUF_X1 U575 ( .A(n3862), .Z(n573) );
  CLKBUF_X1 U576 ( .A(n3864), .Z(n574) );
  CLKBUF_X1 U577 ( .A(n3858), .Z(n575) );
  CLKBUF_X1 U578 ( .A(n3431), .Z(n576) );
  CLKBUF_X1 U579 ( .A(n3721), .Z(n577) );
  AND2_X1 U580 ( .A1(n555), .A2(n1802), .ZN(n578) );
  CLKBUF_X1 U581 ( .A(n2785), .Z(n579) );
  CLKBUF_X1 U582 ( .A(n2696), .Z(n580) );
  CLKBUF_X1 U583 ( .A(n4121), .Z(n581) );
  CLKBUF_X1 U584 ( .A(n4117), .Z(n582) );
  CLKBUF_X1 U585 ( .A(n3796), .Z(n583) );
  AND2_X1 U586 ( .A1(n555), .A2(n2075), .ZN(n584) );
  CLKBUF_X1 U587 ( .A(n4189), .Z(n585) );
  CLKBUF_X1 U588 ( .A(n3965), .Z(n586) );
  AND2_X1 U589 ( .A1(n1115), .A2(n2536), .ZN(n587) );
  CLKBUF_X1 U590 ( .A(n4681), .Z(n588) );
  CLKBUF_X1 U591 ( .A(n964), .Z(n589) );
  CLKBUF_X1 U592 ( .A(n3299), .Z(n590) );
  CLKBUF_X1 U593 ( .A(n2703), .Z(n591) );
  CLKBUF_X1 U594 ( .A(n2705), .Z(n592) );
  CLKBUF_X1 U595 ( .A(n2707), .Z(n593) );
  CLKBUF_X1 U596 ( .A(n2709), .Z(n594) );
  CLKBUF_X1 U597 ( .A(n968), .Z(n595) );
  CLKBUF_X1 U598 ( .A(n3432), .Z(n596) );
  CLKBUF_X1 U599 ( .A(n2718), .Z(n597) );
  CLKBUF_X1 U600 ( .A(n27201), .Z(n598) );
  CLKBUF_X1 U601 ( .A(n970), .Z(n599) );
  CLKBUF_X1 U602 ( .A(n2743), .Z(n600) );
  CLKBUF_X1 U603 ( .A(n2745), .Z(n601) );
  CLKBUF_X1 U604 ( .A(n2747), .Z(n602) );
  CLKBUF_X1 U605 ( .A(n2751), .Z(n603) );
  CLKBUF_X1 U606 ( .A(n3373), .Z(n604) );
  CLKBUF_X1 U607 ( .A(n2754), .Z(n605) );
  CLKBUF_X1 U608 ( .A(n27601), .Z(n606) );
  CLKBUF_X1 U609 ( .A(n2762), .Z(n607) );
  CLKBUF_X1 U610 ( .A(n2764), .Z(n608) );
  CLKBUF_X1 U611 ( .A(n2766), .Z(n609) );
  CLKBUF_X1 U612 ( .A(n2768), .Z(n610) );
  CLKBUF_X1 U613 ( .A(n27701), .Z(n611) );
  CLKBUF_X1 U614 ( .A(n2772), .Z(n612) );
  CLKBUF_X1 U615 ( .A(n2774), .Z(n613) );
  CLKBUF_X1 U616 ( .A(n2776), .Z(n614) );
  CLKBUF_X1 U617 ( .A(n2778), .Z(n615) );
  CLKBUF_X1 U618 ( .A(n27801), .Z(n616) );
  CLKBUF_X1 U619 ( .A(n2782), .Z(n617) );
  CLKBUF_X1 U620 ( .A(n2787), .Z(n618) );
  CLKBUF_X1 U621 ( .A(n2789), .Z(n619) );
  CLKBUF_X1 U622 ( .A(n2791), .Z(n620) );
  CLKBUF_X1 U623 ( .A(n2793), .Z(n621) );
  CLKBUF_X1 U624 ( .A(n2795), .Z(n622) );
  CLKBUF_X1 U625 ( .A(n2797), .Z(n623) );
  CLKBUF_X1 U626 ( .A(n2799), .Z(n624) );
  CLKBUF_X1 U627 ( .A(n2801), .Z(n625) );
  CLKBUF_X1 U628 ( .A(n2803), .Z(n626) );
  CLKBUF_X1 U629 ( .A(n2805), .Z(n627) );
  CLKBUF_X1 U630 ( .A(n2807), .Z(n628) );
  CLKBUF_X1 U631 ( .A(n2809), .Z(n629) );
  CLKBUF_X1 U632 ( .A(n2811), .Z(n630) );
  CLKBUF_X1 U633 ( .A(n2813), .Z(n631) );
  OR2_X1 U634 ( .A1(n1236), .A2(n2124), .ZN(n632) );
  CLKBUF_X1 U635 ( .A(n3791), .Z(n633) );
  CLKBUF_X1 U636 ( .A(n3793), .Z(n634) );
  CLKBUF_X1 U637 ( .A(n3787), .Z(n635) );
  CLKBUF_X1 U638 ( .A(n3789), .Z(n636) );
  CLKBUF_X1 U639 ( .A(n3783), .Z(n637) );
  CLKBUF_X1 U640 ( .A(n3785), .Z(n638) );
  CLKBUF_X1 U641 ( .A(n3779), .Z(n639) );
  CLKBUF_X1 U642 ( .A(n3781), .Z(n640) );
  CLKBUF_X1 U643 ( .A(n3775), .Z(n641) );
  CLKBUF_X1 U644 ( .A(n3777), .Z(n642) );
  CLKBUF_X1 U645 ( .A(n3771), .Z(n643) );
  CLKBUF_X1 U646 ( .A(n3773), .Z(n644) );
  CLKBUF_X1 U647 ( .A(n3767), .Z(n645) );
  CLKBUF_X1 U648 ( .A(n3769), .Z(n646) );
  CLKBUF_X1 U649 ( .A(n3762), .Z(n647) );
  CLKBUF_X1 U650 ( .A(n3765), .Z(n648) );
  CLKBUF_X1 U651 ( .A(n3428), .Z(n649) );
  CLKBUF_X1 U652 ( .A(n2112), .Z(n650) );
  CLKBUF_X1 U653 ( .A(n2915), .Z(n651) );
  CLKBUF_X1 U654 ( .A(n2107), .Z(n652) );
  CLKBUF_X1 U655 ( .A(n2925), .Z(n653) );
  CLKBUF_X1 U656 ( .A(n2728), .Z(n654) );
  CLKBUF_X1 U657 ( .A(n1767), .Z(n655) );
  CLKBUF_X1 U658 ( .A(n3708), .Z(n656) );
  INV_X1 U659 ( .A(n966), .ZN(n657) );
  INV_X1 U660 ( .A(n657), .ZN(n658) );
  INV_X1 U661 ( .A(n657), .ZN(n659) );
  CLKBUF_X1 U662 ( .A(n536), .Z(n660) );
  CLKBUF_X1 U663 ( .A(n4675), .Z(n661) );
  CLKBUF_X1 U664 ( .A(n3961), .Z(n662) );
  CLKBUF_X1 U665 ( .A(n662), .Z(n663) );
  CLKBUF_X1 U666 ( .A(n526), .Z(n664) );
  CLKBUF_X1 U667 ( .A(n521), .Z(n665) );
  CLKBUF_X1 U668 ( .A(n516), .Z(n666) );
  CLKBUF_X1 U669 ( .A(n3956), .Z(n667) );
  CLKBUF_X1 U670 ( .A(n3954), .Z(n668) );
  CLKBUF_X1 U671 ( .A(n3952), .Z(n669) );
  CLKBUF_X1 U672 ( .A(n496), .Z(n670) );
  CLKBUF_X1 U673 ( .A(n3949), .Z(n671) );
  CLKBUF_X1 U674 ( .A(n4860), .Z(n672) );
  CLKBUF_X1 U675 ( .A(n4810), .Z(n673) );
  CLKBUF_X1 U676 ( .A(n4760), .Z(n674) );
  CLKBUF_X1 U677 ( .A(n3944), .Z(n675) );
  CLKBUF_X1 U678 ( .A(n675), .Z(n676) );
  CLKBUF_X1 U679 ( .A(n46600), .Z(n677) );
  CLKBUF_X1 U680 ( .A(n46100), .Z(n678) );
  CLKBUF_X1 U681 ( .A(n541), .Z(n679) );
  CLKBUF_X1 U682 ( .A(n3869), .Z(n680) );
  CLKBUF_X1 U683 ( .A(n1467), .Z(n681) );
  CLKBUF_X1 U684 ( .A(n3711), .Z(n682) );
  CLKBUF_X1 U685 ( .A(n2942), .Z(n683) );
  CLKBUF_X1 U686 ( .A(n1189), .Z(n684) );
  CLKBUF_X1 U687 ( .A(n1477), .Z(n685) );
  CLKBUF_X1 U688 ( .A(n1472), .Z(n686) );
  CLKBUF_X1 U689 ( .A(n14801), .Z(n687) );
  CLKBUF_X1 U690 ( .A(n1195), .Z(n688) );
  CLKBUF_X1 U691 ( .A(n1483), .Z(n689) );
  CLKBUF_X1 U692 ( .A(n14701), .Z(n690) );
  CLKBUF_X1 U693 ( .A(n1486), .Z(n691) );
  CLKBUF_X1 U694 ( .A(n3425), .Z(n692) );
  CLKBUF_X1 U695 ( .A(n3016), .Z(n693) );
  CLKBUF_X1 U696 ( .A(n1497), .Z(n694) );
  CLKBUF_X1 U697 ( .A(n1489), .Z(n695) );
  CLKBUF_X1 U698 ( .A(n15001), .Z(n696) );
  CLKBUF_X1 U699 ( .A(n12201), .Z(n697) );
  CLKBUF_X1 U700 ( .A(n1503), .Z(n698) );
  CLKBUF_X1 U701 ( .A(n2582), .Z(n699) );
  CLKBUF_X1 U702 ( .A(n2578), .Z(n700) );
  CLKBUF_X1 U703 ( .A(n2574), .Z(n701) );
  CLKBUF_X1 U704 ( .A(n2573), .Z(n702) );
  CLKBUF_X1 U705 ( .A(n2566), .Z(n703) );
  CLKBUF_X1 U706 ( .A(n2565), .Z(n704) );
  CLKBUF_X1 U707 ( .A(n2562), .Z(n705) );
  CLKBUF_X1 U708 ( .A(n2561), .Z(n706) );
  CLKBUF_X1 U709 ( .A(n2564), .Z(n707) );
  CLKBUF_X1 U710 ( .A(n2563), .Z(n708) );
  CLKBUF_X1 U711 ( .A(n2559), .Z(n709) );
  CLKBUF_X1 U712 ( .A(n25601), .Z(n710) );
  CLKBUF_X1 U713 ( .A(n1205), .Z(n711) );
  CLKBUF_X1 U714 ( .A(n2557), .Z(n712) );
  CLKBUF_X1 U715 ( .A(n2558), .Z(n713) );
  CLKBUF_X1 U716 ( .A(n2552), .Z(n714) );
  CLKBUF_X1 U717 ( .A(n2553), .Z(n715) );
  CLKBUF_X1 U718 ( .A(n2549), .Z(n716) );
  CLKBUF_X1 U719 ( .A(n2548), .Z(n717) );
  CLKBUF_X1 U720 ( .A(n2545), .Z(n718) );
  CLKBUF_X1 U721 ( .A(n4101), .Z(n719) );
  CLKBUF_X1 U722 ( .A(n1619), .Z(n720) );
  CLKBUF_X1 U723 ( .A(n39701), .Z(n721) );
  CLKBUF_X1 U724 ( .A(n1622), .Z(n722) );
  CLKBUF_X1 U725 ( .A(n4002), .Z(n723) );
  CLKBUF_X1 U726 ( .A(n16250), .Z(n724) );
  CLKBUF_X1 U727 ( .A(n4136), .Z(n725) );
  CLKBUF_X1 U728 ( .A(n16280), .Z(n726) );
  CLKBUF_X1 U729 ( .A(n4611), .Z(n727) );
  CLKBUF_X1 U730 ( .A(n16310), .Z(n728) );
  CLKBUF_X1 U731 ( .A(n4134), .Z(n729) );
  CLKBUF_X1 U732 ( .A(n16340), .Z(n730) );
  CLKBUF_X1 U733 ( .A(n4135), .Z(n731) );
  CLKBUF_X1 U734 ( .A(n16370), .Z(n732) );
  CLKBUF_X1 U735 ( .A(n41001), .Z(n733) );
  CLKBUF_X1 U736 ( .A(n16401), .Z(n734) );
  CLKBUF_X1 U737 ( .A(n3967), .Z(n735) );
  CLKBUF_X1 U738 ( .A(n1643), .Z(n736) );
  CLKBUF_X1 U739 ( .A(n4098), .Z(n737) );
  CLKBUF_X1 U740 ( .A(n1646), .Z(n738) );
  CLKBUF_X1 U741 ( .A(n4137), .Z(n739) );
  CLKBUF_X1 U742 ( .A(n1649), .Z(n740) );
  CLKBUF_X1 U743 ( .A(n4679), .Z(n741) );
  CLKBUF_X1 U744 ( .A(n1652), .Z(n742) );
  CLKBUF_X1 U745 ( .A(n4127), .Z(n743) );
  CLKBUF_X1 U746 ( .A(n1655), .Z(n744) );
  CLKBUF_X1 U747 ( .A(n4124), .Z(n745) );
  CLKBUF_X1 U748 ( .A(n1658), .Z(n746) );
  CLKBUF_X1 U749 ( .A(n4123), .Z(n747) );
  CLKBUF_X1 U750 ( .A(n1661), .Z(n748) );
  CLKBUF_X1 U751 ( .A(n4126), .Z(n749) );
  CLKBUF_X1 U752 ( .A(n1664), .Z(n750) );
  CLKBUF_X1 U753 ( .A(n4041), .Z(n751) );
  CLKBUF_X1 U754 ( .A(n1667), .Z(n752) );
  CLKBUF_X1 U755 ( .A(n4122), .Z(n753) );
  CLKBUF_X1 U756 ( .A(n16701), .Z(n754) );
  CLKBUF_X1 U757 ( .A(n1673), .Z(n755) );
  CLKBUF_X1 U758 ( .A(n4194), .Z(n756) );
  CLKBUF_X1 U759 ( .A(n1676), .Z(n757) );
  CLKBUF_X1 U760 ( .A(n4607), .Z(n758) );
  CLKBUF_X1 U761 ( .A(n1679), .Z(n759) );
  CLKBUF_X1 U762 ( .A(n44701), .Z(n760) );
  CLKBUF_X1 U763 ( .A(n1682), .Z(n761) );
  CLKBUF_X1 U764 ( .A(n4539), .Z(n762) );
  CLKBUF_X1 U765 ( .A(n1685), .Z(n763) );
  CLKBUF_X1 U766 ( .A(n4334), .Z(n764) );
  CLKBUF_X1 U767 ( .A(n1688), .Z(n765) );
  CLKBUF_X1 U768 ( .A(n4404), .Z(n766) );
  CLKBUF_X1 U769 ( .A(n1691), .Z(n767) );
  CLKBUF_X1 U770 ( .A(n4192), .Z(n768) );
  CLKBUF_X1 U771 ( .A(n1694), .Z(n769) );
  CLKBUF_X1 U772 ( .A(n4265), .Z(n770) );
  CLKBUF_X1 U773 ( .A(n1697), .Z(n771) );
  CLKBUF_X1 U774 ( .A(n3799), .Z(n772) );
  CLKBUF_X1 U775 ( .A(n17001), .Z(n773) );
  CLKBUF_X1 U776 ( .A(n3835), .Z(n774) );
  CLKBUF_X1 U777 ( .A(n1703), .Z(n775) );
  CLKBUF_X1 U778 ( .A(n3726), .Z(n776) );
  CLKBUF_X1 U779 ( .A(n1706), .Z(n777) );
  CLKBUF_X1 U780 ( .A(n3764), .Z(n778) );
  CLKBUF_X1 U781 ( .A(n1709), .Z(n779) );
  CLKBUF_X1 U782 ( .A(n3871), .Z(n780) );
  CLKBUF_X1 U783 ( .A(n1721), .Z(n781) );
  CLKBUF_X1 U784 ( .A(n3942), .Z(n782) );
  CLKBUF_X1 U785 ( .A(n1724), .Z(n783) );
  CLKBUF_X1 U786 ( .A(n3907), .Z(n784) );
  CLKBUF_X1 U787 ( .A(n1727), .Z(n785) );
  CLKBUF_X1 U788 ( .A(n4023), .Z(n786) );
  CLKBUF_X1 U789 ( .A(n17301), .Z(n787) );
  CLKBUF_X1 U790 ( .A(n1733), .Z(n788) );
  CLKBUF_X1 U791 ( .A(n4043), .Z(n789) );
  CLKBUF_X1 U792 ( .A(n1736), .Z(n790) );
  CLKBUF_X1 U793 ( .A(n4097), .Z(n791) );
  CLKBUF_X1 U794 ( .A(n1739), .Z(n792) );
  CLKBUF_X1 U795 ( .A(n4139), .Z(n793) );
  CLKBUF_X1 U796 ( .A(n41401), .Z(n794) );
  CLKBUF_X1 U797 ( .A(n3707), .Z(n795) );
  CLKBUF_X1 U798 ( .A(n1135), .Z(n796) );
  CLKBUF_X1 U799 ( .A(n1766), .Z(n797) );
  CLKBUF_X1 U800 ( .A(n1285), .Z(n798) );
  CLKBUF_X1 U801 ( .A(n2104), .Z(n799) );
  CLKBUF_X1 U802 ( .A(n3424), .Z(n800) );
  CLKBUF_X1 U803 ( .A(n3421), .Z(n801) );
  CLKBUF_X1 U804 ( .A(n1219), .Z(n802) );
  CLKBUF_X1 U805 ( .A(n1213), .Z(n803) );
  CLKBUF_X1 U806 ( .A(n4474), .Z(n804) );
  CLKBUF_X1 U807 ( .A(n12101), .Z(n805) );
  CLKBUF_X1 U808 ( .A(n1212), .Z(n806) );
  CLKBUF_X1 U809 ( .A(n3213), .Z(n807) );
  CLKBUF_X1 U810 ( .A(n2131), .Z(n808) );
  CLKBUF_X1 U811 ( .A(n4095), .Z(n809) );
  CLKBUF_X1 U812 ( .A(n3905), .Z(n810) );
  CLKBUF_X1 U813 ( .A(n3908), .Z(n811) );
  CLKBUF_X1 U814 ( .A(n39101), .Z(n812) );
  CLKBUF_X1 U815 ( .A(n3912), .Z(n813) );
  CLKBUF_X1 U816 ( .A(n3914), .Z(n814) );
  CLKBUF_X1 U817 ( .A(n3916), .Z(n815) );
  CLKBUF_X1 U818 ( .A(n3918), .Z(n816) );
  CLKBUF_X1 U819 ( .A(n39201), .Z(n817) );
  CLKBUF_X1 U820 ( .A(n3922), .Z(n818) );
  CLKBUF_X1 U821 ( .A(n3924), .Z(n819) );
  CLKBUF_X1 U822 ( .A(n3926), .Z(n820) );
  CLKBUF_X1 U823 ( .A(n3928), .Z(n821) );
  CLKBUF_X1 U824 ( .A(n39301), .Z(n822) );
  CLKBUF_X1 U825 ( .A(n3932), .Z(n823) );
  CLKBUF_X1 U826 ( .A(n3934), .Z(n824) );
  CLKBUF_X1 U827 ( .A(n3936), .Z(n825) );
  CLKBUF_X1 U828 ( .A(n1757), .Z(n826) );
  CLKBUF_X1 U829 ( .A(n26901), .Z(n827) );
  CLKBUF_X1 U830 ( .A(n1123), .Z(n828) );
  CLKBUF_X1 U831 ( .A(n1134), .Z(n829) );
  CLKBUF_X1 U832 ( .A(n1492), .Z(n830) );
  CLKBUF_X1 U833 ( .A(n2587), .Z(n831) );
  CLKBUF_X1 U834 ( .A(n1524), .Z(n832) );
  CLKBUF_X1 U835 ( .A(n1529), .Z(n833) );
  CLKBUF_X1 U836 ( .A(n2911), .Z(n834) );
  CLKBUF_X1 U837 ( .A(n2911), .Z(n835) );
  CLKBUF_X1 U838 ( .A(n2689), .Z(n836) );
  CLKBUF_X1 U839 ( .A(n15610), .Z(n837) );
  CLKBUF_X1 U840 ( .A(n2118), .Z(n838) );
  CLKBUF_X1 U841 ( .A(n4676), .Z(n839) );
  CLKBUF_X1 U842 ( .A(n4021), .Z(n840) );
  CLKBUF_X1 U843 ( .A(n840), .Z(n841) );
  CLKBUF_X1 U844 ( .A(n2226), .Z(n842) );
  CLKBUF_X1 U845 ( .A(n4678), .Z(n843) );
  CLKBUF_X1 U846 ( .A(n2226), .Z(n844) );
  CLKBUF_X1 U847 ( .A(n2242), .Z(n845) );
  CLKBUF_X1 U848 ( .A(n2242), .Z(n846) );
  CLKBUF_X1 U849 ( .A(n4138), .Z(n847) );
  CLKBUF_X1 U850 ( .A(n2249), .Z(n848) );
  CLKBUF_X1 U851 ( .A(n2248), .Z(n849) );
  CLKBUF_X1 U852 ( .A(n3318), .Z(n850) );
  CLKBUF_X1 U853 ( .A(n2273), .Z(n851) );
  CLKBUF_X1 U854 ( .A(n2272), .Z(n852) );
  CLKBUF_X1 U855 ( .A(n3317), .Z(n853) );
  CLKBUF_X1 U856 ( .A(n3795), .Z(n854) );
  CLKBUF_X1 U857 ( .A(n3761), .Z(n855) );
  CLKBUF_X1 U858 ( .A(n2295), .Z(n856) );
  CLKBUF_X1 U859 ( .A(n2294), .Z(n857) );
  CLKBUF_X1 U860 ( .A(n23201), .Z(n858) );
  CLKBUF_X1 U861 ( .A(n2319), .Z(n859) );
  CLKBUF_X1 U862 ( .A(n3316), .Z(n860) );
  CLKBUF_X1 U863 ( .A(n4469), .Z(n861) );
  CLKBUF_X1 U864 ( .A(n4403), .Z(n862) );
  CLKBUF_X1 U865 ( .A(n2342), .Z(n863) );
  CLKBUF_X1 U866 ( .A(n2341), .Z(n864) );
  CLKBUF_X1 U867 ( .A(n2367), .Z(n865) );
  CLKBUF_X1 U868 ( .A(n2366), .Z(n866) );
  CLKBUF_X1 U869 ( .A(n3315), .Z(n867) );
  CLKBUF_X1 U870 ( .A(n3902), .Z(n868) );
  CLKBUF_X1 U871 ( .A(n3868), .Z(n869) );
  CLKBUF_X1 U872 ( .A(n2389), .Z(n870) );
  CLKBUF_X1 U873 ( .A(n2388), .Z(n871) );
  CLKBUF_X1 U874 ( .A(n3314), .Z(n872) );
  CLKBUF_X1 U875 ( .A(n3938), .Z(n873) );
  CLKBUF_X1 U876 ( .A(n2408), .Z(n874) );
  CLKBUF_X1 U877 ( .A(n3904), .Z(n875) );
  CLKBUF_X1 U878 ( .A(n2408), .Z(n876) );
  CLKBUF_X1 U879 ( .A(n2409), .Z(n877) );
  CLKBUF_X1 U880 ( .A(n2409), .Z(n878) );
  CLKBUF_X1 U881 ( .A(n2433), .Z(n879) );
  CLKBUF_X1 U882 ( .A(n2432), .Z(n880) );
  CLKBUF_X1 U883 ( .A(n2432), .Z(n881) );
  CLKBUF_X1 U884 ( .A(n2433), .Z(n882) );
  CLKBUF_X1 U885 ( .A(n2454), .Z(n883) );
  CLKBUF_X1 U886 ( .A(n3698), .Z(n884) );
  CLKBUF_X1 U887 ( .A(n884), .Z(n885) );
  CLKBUF_X1 U888 ( .A(n2454), .Z(n886) );
  CLKBUF_X1 U889 ( .A(n2455), .Z(n887) );
  CLKBUF_X1 U890 ( .A(n3699), .Z(n888) );
  CLKBUF_X1 U891 ( .A(n2455), .Z(n889) );
  CLKBUF_X1 U892 ( .A(n2477), .Z(n890) );
  CLKBUF_X1 U893 ( .A(n3704), .Z(n891) );
  CLKBUF_X1 U894 ( .A(n891), .Z(n892) );
  CLKBUF_X1 U895 ( .A(n2477), .Z(n893) );
  CLKBUF_X1 U896 ( .A(n2476), .Z(n894) );
  CLKBUF_X1 U897 ( .A(n2685), .Z(n895) );
  CLKBUF_X1 U898 ( .A(n2476), .Z(n896) );
  CLKBUF_X1 U899 ( .A(n24901), .Z(n897) );
  CLKBUF_X1 U900 ( .A(n2491), .Z(n898) );
  CLKBUF_X1 U901 ( .A(n24901), .Z(n899) );
  CLKBUF_X1 U902 ( .A(n2491), .Z(n900) );
  CLKBUF_X1 U903 ( .A(n2497), .Z(n901) );
  CLKBUF_X1 U904 ( .A(n2684), .Z(n902) );
  CLKBUF_X1 U905 ( .A(n2497), .Z(n903) );
  CLKBUF_X1 U906 ( .A(n2498), .Z(n904) );
  CLKBUF_X1 U907 ( .A(n2498), .Z(n905) );
  CLKBUF_X1 U908 ( .A(n2515), .Z(n906) );
  CLKBUF_X1 U909 ( .A(n2514), .Z(n907) );
  CLKBUF_X1 U910 ( .A(n2514), .Z(n908) );
  CLKBUF_X1 U911 ( .A(n2684), .Z(n909) );
  CLKBUF_X1 U912 ( .A(matrix_index[1]), .Z(n910) );
  CLKBUF_X1 U913 ( .A(n912), .Z(n911) );
  AND2_X1 U914 ( .A1(n553), .A2(n2914), .ZN(n912) );
  CLKBUF_X1 U915 ( .A(n3715), .Z(n913) );
  CLKBUF_X1 U916 ( .A(n3706), .Z(n914) );
  CLKBUF_X1 U917 ( .A(n3278), .Z(n915) );
  CLKBUF_X1 U918 ( .A(n2121), .Z(n916) );
  CLKBUF_X1 U919 ( .A(n2555), .Z(n917) );
  CLKBUF_X1 U920 ( .A(n2127), .Z(n918) );
  CLKBUF_X1 U921 ( .A(n21301), .Z(n919) );
  CLKBUF_X1 U922 ( .A(n3265), .Z(n920) );
  CLKBUF_X1 U923 ( .A(n2136), .Z(n921) );
  CLKBUF_X1 U924 ( .A(n2568), .Z(n922) );
  CLKBUF_X1 U925 ( .A(n2571), .Z(n923) );
  CLKBUF_X1 U926 ( .A(n2142), .Z(n9240) );
  CLKBUF_X1 U927 ( .A(N100), .Z(n9250) );
  CLKBUF_X1 U928 ( .A(N102), .Z(n9260) );
  CLKBUF_X1 U929 ( .A(n17701), .Z(n9270) );
  CLKBUF_X1 U930 ( .A(n2152), .Z(n9280) );
  CLKBUF_X1 U931 ( .A(n1217), .Z(n9290) );
  CLKBUF_X1 U932 ( .A(n3423), .Z(n9300) );
  CLKBUF_X1 U933 ( .A(n1778), .Z(n9310) );
  CLKBUF_X1 U934 ( .A(n1519), .Z(n9320) );
  CLKBUF_X1 U935 ( .A(n1783), .Z(n9330) );
  CLKBUF_X1 U936 ( .A(n1516), .Z(n9340) );
  CLKBUF_X1 U937 ( .A(n1214), .Z(n9350) );
  CLKBUF_X1 U938 ( .A(n1513), .Z(n9360) );
  CLKBUF_X1 U939 ( .A(n1789), .Z(n9370) );
  CLKBUF_X1 U940 ( .A(n15101), .Z(n9380) );
  CLKBUF_X1 U941 ( .A(n1199), .Z(n9390) );
  CLKBUF_X1 U942 ( .A(n1507), .Z(n940) );
  CLKBUF_X1 U943 ( .A(n3905), .Z(n941) );
  CLKBUF_X1 U944 ( .A(n3908), .Z(n942) );
  CLKBUF_X1 U945 ( .A(n39101), .Z(n943) );
  CLKBUF_X1 U946 ( .A(n3912), .Z(n944) );
  CLKBUF_X1 U947 ( .A(n3914), .Z(n945) );
  CLKBUF_X1 U948 ( .A(n3916), .Z(n946) );
  CLKBUF_X1 U949 ( .A(n3918), .Z(n947) );
  CLKBUF_X1 U950 ( .A(n39201), .Z(n948) );
  CLKBUF_X1 U951 ( .A(n3922), .Z(n949) );
  CLKBUF_X1 U952 ( .A(n3924), .Z(n950) );
  CLKBUF_X1 U953 ( .A(n3926), .Z(n951) );
  CLKBUF_X1 U954 ( .A(n3928), .Z(n952) );
  CLKBUF_X1 U955 ( .A(n39301), .Z(n953) );
  CLKBUF_X1 U956 ( .A(n3932), .Z(n954) );
  CLKBUF_X1 U957 ( .A(n3934), .Z(n955) );
  CLKBUF_X1 U958 ( .A(n3936), .Z(n956) );
  AND2_X1 U959 ( .A1(n4189), .A2(n548), .ZN(n957) );
  NAND2_X1 U960 ( .A1(n12260), .A2(n1535), .ZN(n958) );
  NOR2_X1 U961 ( .A1(n2216), .A2(n2209), .ZN(n959) );
  XNOR2_X1 U962 ( .A(n3454), .B(n3221), .ZN(n960) );
  CLKBUF_X1 U963 ( .A(n2688), .Z(n961) );
  AND3_X1 U964 ( .A1(n1466), .A2(n2702), .A3(n1361), .ZN(n962) );
  NAND3_X1 U965 ( .A1(n3471), .A2(n34701), .A3(n3446), .ZN(n963) );
  CLKBUF_X1 U966 ( .A(n850), .Z(n964) );
  INV_X1 U967 ( .A(r290_B_3_), .ZN(n965) );
  INV_X1 U968 ( .A(r290_B_3_), .ZN(n966) );
  CLKBUF_X1 U969 ( .A(n3708), .Z(n967) );
  CLKBUF_X1 U970 ( .A(n43401), .Z(n968) );
  CLKBUF_X1 U971 ( .A(n2158), .Z(n969) );
  CLKBUF_X1 U972 ( .A(n4202), .Z(n970) );
  CLKBUF_X1 U973 ( .A(n3826), .Z(n971) );
  CLKBUF_X1 U974 ( .A(n3828), .Z(n972) );
  CLKBUF_X1 U975 ( .A(n3822), .Z(n973) );
  CLKBUF_X1 U976 ( .A(n3824), .Z(n974) );
  CLKBUF_X1 U977 ( .A(n3818), .Z(n975) );
  CLKBUF_X1 U978 ( .A(n38201), .Z(n976) );
  CLKBUF_X1 U979 ( .A(n3814), .Z(n977) );
  CLKBUF_X1 U980 ( .A(n3816), .Z(n978) );
  CLKBUF_X1 U981 ( .A(n38101), .Z(n979) );
  CLKBUF_X1 U982 ( .A(n3812), .Z(n980) );
  CLKBUF_X1 U983 ( .A(n3806), .Z(n981) );
  CLKBUF_X1 U984 ( .A(n3808), .Z(n982) );
  CLKBUF_X1 U985 ( .A(n3802), .Z(n983) );
  CLKBUF_X1 U986 ( .A(n3804), .Z(n984) );
  CLKBUF_X1 U987 ( .A(n3797), .Z(n985) );
  CLKBUF_X1 U988 ( .A(n38001), .Z(n986) );
  CLKBUF_X1 U989 ( .A(n633), .Z(n987) );
  CLKBUF_X1 U990 ( .A(n634), .Z(n988) );
  CLKBUF_X1 U991 ( .A(n635), .Z(n989) );
  CLKBUF_X1 U992 ( .A(n636), .Z(n990) );
  CLKBUF_X1 U993 ( .A(n637), .Z(n991) );
  CLKBUF_X1 U994 ( .A(n638), .Z(n992) );
  CLKBUF_X1 U995 ( .A(n639), .Z(n993) );
  CLKBUF_X1 U996 ( .A(n640), .Z(n994) );
  CLKBUF_X1 U997 ( .A(n641), .Z(n995) );
  CLKBUF_X1 U998 ( .A(n642), .Z(n996) );
  CLKBUF_X1 U999 ( .A(n643), .Z(n997) );
  CLKBUF_X1 U1000 ( .A(n644), .Z(n998) );
  CLKBUF_X1 U1001 ( .A(n645), .Z(n999) );
  CLKBUF_X1 U1002 ( .A(n646), .Z(n10001) );
  CLKBUF_X1 U1003 ( .A(n647), .Z(n1001) );
  CLKBUF_X1 U1004 ( .A(n648), .Z(n1002) );
  CLKBUF_X1 U1005 ( .A(n3753), .Z(n1003) );
  CLKBUF_X1 U1006 ( .A(n3755), .Z(n1004) );
  CLKBUF_X1 U1007 ( .A(n3749), .Z(n1005) );
  CLKBUF_X1 U1008 ( .A(n3751), .Z(n1006) );
  CLKBUF_X1 U1009 ( .A(n3745), .Z(n1007) );
  CLKBUF_X1 U1010 ( .A(n3747), .Z(n1008) );
  CLKBUF_X1 U1011 ( .A(n3741), .Z(n1009) );
  CLKBUF_X1 U1012 ( .A(n3743), .Z(n10101) );
  CLKBUF_X1 U1013 ( .A(n3737), .Z(n1011) );
  CLKBUF_X1 U1014 ( .A(n3739), .Z(n1012) );
  CLKBUF_X1 U1015 ( .A(n3733), .Z(n1013) );
  CLKBUF_X1 U1016 ( .A(n3735), .Z(n1014) );
  CLKBUF_X1 U1017 ( .A(n3729), .Z(n1015) );
  CLKBUF_X1 U1018 ( .A(n3731), .Z(n1016) );
  CLKBUF_X1 U1019 ( .A(n3724), .Z(n1017) );
  CLKBUF_X1 U1020 ( .A(n3727), .Z(n1018) );
  CLKBUF_X1 U1021 ( .A(n649), .Z(n1019) );
  CLKBUF_X1 U1022 ( .A(n1347), .Z(n10201) );
  CLKBUF_X1 U1023 ( .A(n2109), .Z(n1021) );
  CLKBUF_X1 U1024 ( .A(n650), .Z(n1022) );
  CLKBUF_X1 U1025 ( .A(n651), .Z(n1023) );
  CLKBUF_X1 U1026 ( .A(n652), .Z(n1024) );
  CLKBUF_X1 U1027 ( .A(n1351), .Z(n1025) );
  CLKBUF_X1 U1028 ( .A(n653), .Z(n1026) );
  CLKBUF_X1 U1029 ( .A(n654), .Z(n1027) );
  CLKBUF_X1 U1030 ( .A(n655), .Z(n1028) );
  CLKBUF_X1 U1031 ( .A(n1356), .Z(n1029) );
  CLKBUF_X1 U1032 ( .A(n656), .Z(n10301) );
  CLKBUF_X1 U1033 ( .A(n1359), .Z(n1031) );
  CLKBUF_X1 U1034 ( .A(n1366), .Z(n1032) );
  CLKBUF_X1 U1035 ( .A(n1371), .Z(n1033) );
  CLKBUF_X1 U1036 ( .A(n1378), .Z(n1034) );
  CLKBUF_X1 U1037 ( .A(n1385), .Z(n1035) );
  CLKBUF_X1 U1038 ( .A(n1392), .Z(n1036) );
  CLKBUF_X1 U1039 ( .A(n667), .Z(n1037) );
  CLKBUF_X1 U1040 ( .A(n1397), .Z(n1038) );
  CLKBUF_X1 U1041 ( .A(n668), .Z(n1039) );
  CLKBUF_X1 U1042 ( .A(n1402), .Z(n10401) );
  CLKBUF_X1 U1043 ( .A(n669), .Z(n1041) );
  CLKBUF_X1 U1044 ( .A(n1407), .Z(n1042) );
  CLKBUF_X1 U1045 ( .A(n1414), .Z(n1043) );
  CLKBUF_X1 U1046 ( .A(n671), .Z(n1044) );
  CLKBUF_X1 U1047 ( .A(n1419), .Z(n1045) );
  CLKBUF_X1 U1048 ( .A(n1426), .Z(n1046) );
  CLKBUF_X1 U1049 ( .A(n1433), .Z(n1047) );
  CLKBUF_X1 U1050 ( .A(n14401), .Z(n1048) );
  CLKBUF_X1 U1051 ( .A(n1445), .Z(n1049) );
  CLKBUF_X1 U1052 ( .A(n1452), .Z(n10501) );
  CLKBUF_X1 U1053 ( .A(n1459), .Z(n1051) );
  CLKBUF_X1 U1054 ( .A(n680), .Z(n1052) );
  CLKBUF_X1 U1055 ( .A(n684), .Z(n1053) );
  CLKBUF_X1 U1056 ( .A(n686), .Z(n1054) );
  CLKBUF_X1 U1057 ( .A(n688), .Z(n1055) );
  CLKBUF_X1 U1058 ( .A(n690), .Z(n1056) );
  CLKBUF_X1 U1059 ( .A(n693), .Z(n1057) );
  CLKBUF_X1 U1060 ( .A(n695), .Z(n1058) );
  CLKBUF_X1 U1061 ( .A(n697), .Z(n1059) );
  CLKBUF_X1 U1062 ( .A(n1209), .Z(n10601) );
  CLKBUF_X1 U1063 ( .A(n597), .Z(n1061) );
  CLKBUF_X1 U1064 ( .A(n599), .Z(n1062) );
  INV_X1 U1065 ( .A(n2145), .ZN(n3424) );
  AND2_X1 U1066 ( .A1(n553), .A2(n10201), .ZN(n1063) );
  CLKBUF_X1 U1067 ( .A(n2544), .Z(n1064) );
  CLKBUF_X1 U1068 ( .A(n719), .Z(n1065) );
  CLKBUF_X1 U1069 ( .A(n721), .Z(n1066) );
  CLKBUF_X1 U1070 ( .A(n723), .Z(n1067) );
  CLKBUF_X1 U1071 ( .A(n725), .Z(n1068) );
  CLKBUF_X1 U1072 ( .A(n727), .Z(n1069) );
  CLKBUF_X1 U1073 ( .A(n729), .Z(n10701) );
  CLKBUF_X1 U1074 ( .A(n731), .Z(n1071) );
  CLKBUF_X1 U1075 ( .A(n733), .Z(n1072) );
  CLKBUF_X1 U1076 ( .A(n735), .Z(n1073) );
  CLKBUF_X1 U1077 ( .A(n737), .Z(n1074) );
  CLKBUF_X1 U1078 ( .A(n739), .Z(n1075) );
  CLKBUF_X1 U1079 ( .A(n741), .Z(n1076) );
  CLKBUF_X1 U1080 ( .A(n743), .Z(n1077) );
  CLKBUF_X1 U1081 ( .A(n745), .Z(n1078) );
  CLKBUF_X1 U1082 ( .A(n747), .Z(n1079) );
  CLKBUF_X1 U1083 ( .A(n749), .Z(n10801) );
  CLKBUF_X1 U1084 ( .A(n751), .Z(n1081) );
  CLKBUF_X1 U1085 ( .A(n753), .Z(n1082) );
  CLKBUF_X1 U1086 ( .A(n1124), .Z(n1083) );
  CLKBUF_X1 U1087 ( .A(n756), .Z(n1084) );
  CLKBUF_X1 U1088 ( .A(n758), .Z(n1085) );
  CLKBUF_X1 U1089 ( .A(n760), .Z(n1086) );
  CLKBUF_X1 U1090 ( .A(n762), .Z(n1087) );
  CLKBUF_X1 U1091 ( .A(n764), .Z(n1088) );
  CLKBUF_X1 U1092 ( .A(n766), .Z(n1089) );
  CLKBUF_X1 U1093 ( .A(n768), .Z(n10901) );
  CLKBUF_X1 U1094 ( .A(n770), .Z(n1091) );
  CLKBUF_X1 U1095 ( .A(n772), .Z(n1092) );
  CLKBUF_X1 U1096 ( .A(n774), .Z(n1093) );
  CLKBUF_X1 U1097 ( .A(n776), .Z(n1094) );
  CLKBUF_X1 U1098 ( .A(n778), .Z(n1095) );
  CLKBUF_X1 U1099 ( .A(n1717), .Z(n1096) );
  CLKBUF_X1 U1100 ( .A(n780), .Z(n1097) );
  CLKBUF_X1 U1101 ( .A(n782), .Z(n1098) );
  CLKBUF_X1 U1102 ( .A(n784), .Z(n1099) );
  CLKBUF_X1 U1103 ( .A(n786), .Z(n11001) );
  CLKBUF_X1 U1104 ( .A(n1126), .Z(n1101) );
  CLKBUF_X1 U1105 ( .A(n789), .Z(n1102) );
  CLKBUF_X1 U1106 ( .A(n791), .Z(n1103) );
  CLKBUF_X1 U1107 ( .A(n1742), .Z(n1104) );
  CLKBUF_X1 U1108 ( .A(n1747), .Z(n1105) );
  CLKBUF_X1 U1109 ( .A(n793), .Z(n1106) );
  CLKBUF_X1 U1110 ( .A(n794), .Z(n1107) );
  CLKBUF_X1 U1111 ( .A(n795), .Z(n1108) );
  CLKBUF_X1 U1112 ( .A(n595), .Z(n1109) );
  CLKBUF_X1 U1113 ( .A(n796), .Z(n11101) );
  CLKBUF_X1 U1114 ( .A(n1761), .Z(n1111) );
  CLKBUF_X1 U1115 ( .A(n1763), .Z(n1112) );
  CLKBUF_X1 U1116 ( .A(n1765), .Z(n1113) );
  CLKBUF_X1 U1117 ( .A(n800), .Z(n1114) );
  CLKBUF_X1 U1118 ( .A(n801), .Z(n1115) );
  CLKBUF_X1 U1119 ( .A(n804), .Z(n1116) );
  CLKBUF_X1 U1120 ( .A(n1211), .Z(n1117) );
  CLKBUF_X1 U1121 ( .A(n1207), .Z(n1118) );
  CLKBUF_X1 U1122 ( .A(n594), .Z(n1119) );
  CLKBUF_X1 U1123 ( .A(n1793), .Z(n11201) );
  CLKBUF_X1 U1124 ( .A(n2159), .Z(n1121) );
  CLKBUF_X1 U1125 ( .A(n807), .Z(n1122) );
  INV_X1 U1126 ( .A(n4131), .ZN(n1123) );
  INV_X1 U1127 ( .A(n1123), .ZN(n1124) );
  INV_X1 U1128 ( .A(n4201), .ZN(n1125) );
  INV_X1 U1129 ( .A(n1125), .ZN(n1126) );
  INV_X1 U1130 ( .A(n1125), .ZN(n1127) );
  INV_X1 U1131 ( .A(n584), .ZN(n1128) );
  INV_X1 U1132 ( .A(n584), .ZN(n1129) );
  INV_X1 U1133 ( .A(n587), .ZN(n11301) );
  INV_X1 U1134 ( .A(n587), .ZN(n1131) );
  INV_X1 U1135 ( .A(n4683), .ZN(n1132) );
  INV_X1 U1136 ( .A(n1132), .ZN(n1133) );
  INV_X1 U1137 ( .A(n2029), .ZN(n1134) );
  INV_X1 U1138 ( .A(n1134), .ZN(n1135) );
  INV_X1 U1139 ( .A(n589), .ZN(n1136) );
  INV_X1 U1140 ( .A(n589), .ZN(n1137) );
  INV_X1 U1141 ( .A(n3862), .ZN(n1138) );
  INV_X1 U1142 ( .A(n1138), .ZN(n1139) );
  INV_X1 U1143 ( .A(n1138), .ZN(n11401) );
  INV_X1 U1144 ( .A(n3864), .ZN(n1141) );
  INV_X1 U1145 ( .A(n1141), .ZN(n1142) );
  INV_X1 U1146 ( .A(n1141), .ZN(n1143) );
  INV_X1 U1147 ( .A(n3858), .ZN(n1144) );
  INV_X1 U1148 ( .A(n1144), .ZN(n1145) );
  INV_X1 U1149 ( .A(n1144), .ZN(n1146) );
  INV_X1 U1150 ( .A(n38601), .ZN(n1147) );
  INV_X1 U1151 ( .A(n1147), .ZN(n1148) );
  INV_X1 U1152 ( .A(n1147), .ZN(n1149) );
  INV_X1 U1153 ( .A(n3854), .ZN(n11501) );
  INV_X1 U1154 ( .A(n11501), .ZN(n1151) );
  INV_X1 U1155 ( .A(n11501), .ZN(n1152) );
  INV_X1 U1156 ( .A(n3856), .ZN(n1153) );
  INV_X1 U1157 ( .A(n1153), .ZN(n1154) );
  INV_X1 U1158 ( .A(n1153), .ZN(n1155) );
  INV_X1 U1159 ( .A(n38501), .ZN(n1156) );
  INV_X1 U1160 ( .A(n1156), .ZN(n1157) );
  INV_X1 U1161 ( .A(n1156), .ZN(n1158) );
  INV_X1 U1162 ( .A(n3852), .ZN(n1159) );
  INV_X1 U1163 ( .A(n1159), .ZN(n11601) );
  INV_X1 U1164 ( .A(n1159), .ZN(n1161) );
  INV_X1 U1165 ( .A(n3846), .ZN(n1162) );
  INV_X1 U1166 ( .A(n1162), .ZN(n1163) );
  INV_X1 U1167 ( .A(n1162), .ZN(n1164) );
  INV_X1 U1168 ( .A(n3848), .ZN(n1165) );
  INV_X1 U1169 ( .A(n1165), .ZN(n1166) );
  INV_X1 U1170 ( .A(n1165), .ZN(n1167) );
  INV_X1 U1171 ( .A(n3842), .ZN(n1168) );
  INV_X1 U1172 ( .A(n1168), .ZN(n1169) );
  INV_X1 U1173 ( .A(n1168), .ZN(n11701) );
  INV_X1 U1174 ( .A(n3844), .ZN(n1171) );
  INV_X1 U1175 ( .A(n1171), .ZN(n1172) );
  INV_X1 U1176 ( .A(n1171), .ZN(n1173) );
  INV_X1 U1177 ( .A(n3838), .ZN(n1174) );
  INV_X1 U1178 ( .A(n1174), .ZN(n1175) );
  INV_X1 U1179 ( .A(n1174), .ZN(n1176) );
  INV_X1 U1180 ( .A(n38401), .ZN(n1177) );
  INV_X1 U1181 ( .A(n1177), .ZN(n1178) );
  INV_X1 U1182 ( .A(n1177), .ZN(n1179) );
  INV_X1 U1183 ( .A(n3833), .ZN(n11801) );
  INV_X1 U1184 ( .A(n11801), .ZN(n1181) );
  INV_X1 U1185 ( .A(n11801), .ZN(n1182) );
  INV_X1 U1186 ( .A(n3836), .ZN(n1183) );
  INV_X1 U1187 ( .A(n1183), .ZN(n1184) );
  INV_X1 U1188 ( .A(n1183), .ZN(n1185) );
  INV_X1 U1189 ( .A(n590), .ZN(n1186) );
  INV_X1 U1190 ( .A(n590), .ZN(n1187) );
  INV_X1 U1191 ( .A(n967), .ZN(n1188) );
  INV_X1 U1192 ( .A(n1188), .ZN(n1189) );
  INV_X1 U1193 ( .A(n1188), .ZN(n11901) );
  INV_X1 U1194 ( .A(n2701), .ZN(n1191) );
  INV_X1 U1195 ( .A(n1191), .ZN(n1192) );
  INV_X1 U1196 ( .A(n1191), .ZN(n1193) );
  INV_X1 U1197 ( .A(n967), .ZN(n1194) );
  INV_X1 U1198 ( .A(n1194), .ZN(n1195) );
  INV_X1 U1199 ( .A(n1194), .ZN(n1196) );
  INV_X1 U1200 ( .A(n591), .ZN(n1197) );
  INV_X1 U1201 ( .A(n591), .ZN(n1198) );
  INV_X1 U1202 ( .A(n592), .ZN(n1199) );
  INV_X1 U1203 ( .A(n592), .ZN(n12001) );
  INV_X1 U1204 ( .A(n593), .ZN(n1201) );
  INV_X1 U1205 ( .A(n593), .ZN(n1202) );
  INV_X1 U1206 ( .A(n594), .ZN(n1203) );
  INV_X1 U1207 ( .A(n595), .ZN(n1204) );
  INV_X1 U1208 ( .A(n596), .ZN(n1205) );
  INV_X1 U1209 ( .A(n596), .ZN(n1206) );
  INV_X1 U1210 ( .A(n2714), .ZN(n1207) );
  INV_X1 U1211 ( .A(n1207), .ZN(n1208) );
  INV_X1 U1212 ( .A(n4272), .ZN(n1209) );
  INV_X1 U1213 ( .A(n1209), .ZN(n12101) );
  INV_X1 U1214 ( .A(n969), .ZN(n1211) );
  INV_X1 U1215 ( .A(n1211), .ZN(n1212) );
  INV_X1 U1216 ( .A(n597), .ZN(n1213) );
  INV_X1 U1217 ( .A(n598), .ZN(n1214) );
  INV_X1 U1218 ( .A(n598), .ZN(n1215) );
  INV_X1 U1219 ( .A(n33201), .ZN(n1216) );
  INV_X1 U1220 ( .A(n1216), .ZN(n1217) );
  INV_X1 U1221 ( .A(n1216), .ZN(n1218) );
  INV_X1 U1222 ( .A(n599), .ZN(n1219) );
  INV_X1 U1223 ( .A(n600), .ZN(n12201) );
  INV_X1 U1224 ( .A(n600), .ZN(n1221) );
  INV_X1 U1225 ( .A(n601), .ZN(n1222) );
  INV_X1 U1226 ( .A(n601), .ZN(n1223) );
  INV_X1 U1227 ( .A(n602), .ZN(n1224) );
  INV_X1 U1228 ( .A(n602), .ZN(n12250) );
  INV_X1 U1229 ( .A(n603), .ZN(n12260) );
  INV_X1 U1230 ( .A(n603), .ZN(n1227) );
  INV_X1 U1231 ( .A(n604), .ZN(n12280) );
  INV_X1 U1232 ( .A(n604), .ZN(n12290) );
  INV_X1 U1233 ( .A(n605), .ZN(n12301) );
  INV_X1 U1234 ( .A(n605), .ZN(n1231) );
  INV_X1 U1235 ( .A(n606), .ZN(n1232) );
  INV_X1 U1236 ( .A(n606), .ZN(n1233) );
  INV_X1 U1237 ( .A(n607), .ZN(n1234) );
  INV_X1 U1238 ( .A(n607), .ZN(n1235) );
  INV_X1 U1239 ( .A(n608), .ZN(n1236) );
  INV_X1 U1240 ( .A(n608), .ZN(n1237) );
  INV_X1 U1241 ( .A(n609), .ZN(n1238) );
  INV_X1 U1242 ( .A(n609), .ZN(n1239) );
  INV_X1 U1243 ( .A(n610), .ZN(n12401) );
  INV_X1 U1244 ( .A(n610), .ZN(n1241) );
  INV_X1 U1245 ( .A(n611), .ZN(n1242) );
  INV_X1 U1246 ( .A(n611), .ZN(n1243) );
  INV_X1 U1247 ( .A(n4142), .ZN(n1244) );
  INV_X1 U1248 ( .A(n1244), .ZN(n1245) );
  INV_X1 U1249 ( .A(n1244), .ZN(n1246) );
  INV_X1 U1250 ( .A(n612), .ZN(n1247) );
  INV_X1 U1251 ( .A(n612), .ZN(n1248) );
  INV_X1 U1252 ( .A(n613), .ZN(n1249) );
  INV_X1 U1253 ( .A(n613), .ZN(n12501) );
  INV_X1 U1254 ( .A(n614), .ZN(n1251) );
  INV_X1 U1255 ( .A(n614), .ZN(n1252) );
  INV_X1 U1256 ( .A(n615), .ZN(n1253) );
  INV_X1 U1257 ( .A(n615), .ZN(n1254) );
  INV_X1 U1258 ( .A(n616), .ZN(n1255) );
  INV_X1 U1259 ( .A(n616), .ZN(n1256) );
  INV_X1 U1260 ( .A(n617), .ZN(n1257) );
  INV_X1 U1261 ( .A(n617), .ZN(n1258) );
  INV_X1 U1262 ( .A(n618), .ZN(n1259) );
  INV_X1 U1263 ( .A(n618), .ZN(n12601) );
  INV_X1 U1264 ( .A(n619), .ZN(n1261) );
  INV_X1 U1265 ( .A(n619), .ZN(n1262) );
  INV_X1 U1266 ( .A(n620), .ZN(n1263) );
  INV_X1 U1267 ( .A(n620), .ZN(n1264) );
  INV_X1 U1268 ( .A(n621), .ZN(n1265) );
  INV_X1 U1269 ( .A(n621), .ZN(n1266) );
  INV_X1 U1270 ( .A(n622), .ZN(n1267) );
  INV_X1 U1271 ( .A(n622), .ZN(n1268) );
  INV_X1 U1272 ( .A(n623), .ZN(n1269) );
  INV_X1 U1273 ( .A(n623), .ZN(n12701) );
  INV_X1 U1274 ( .A(n624), .ZN(n1271) );
  INV_X1 U1275 ( .A(n624), .ZN(n1272) );
  INV_X1 U1276 ( .A(n625), .ZN(n1273) );
  INV_X1 U1277 ( .A(n625), .ZN(n1274) );
  INV_X1 U1278 ( .A(n626), .ZN(n1275) );
  INV_X1 U1279 ( .A(n626), .ZN(n1276) );
  INV_X1 U1280 ( .A(n627), .ZN(n1277) );
  INV_X1 U1281 ( .A(n627), .ZN(n1278) );
  INV_X1 U1282 ( .A(n628), .ZN(n1279) );
  INV_X1 U1283 ( .A(n628), .ZN(n12801) );
  INV_X1 U1284 ( .A(n629), .ZN(n1281) );
  INV_X1 U1285 ( .A(n629), .ZN(n1282) );
  INV_X1 U1286 ( .A(n630), .ZN(n1283) );
  INV_X1 U1287 ( .A(n630), .ZN(n1284) );
  INV_X1 U1288 ( .A(n631), .ZN(n1285) );
  INV_X1 U1289 ( .A(n631), .ZN(n1286) );
  INV_X1 U1290 ( .A(n4673), .ZN(n1287) );
  INV_X1 U1291 ( .A(n1287), .ZN(n1288) );
  INV_X1 U1292 ( .A(n1287), .ZN(n1289) );
  INV_X1 U1293 ( .A(n4188), .ZN(n12901) );
  INV_X1 U1294 ( .A(n12901), .ZN(n1291) );
  INV_X1 U1295 ( .A(n12901), .ZN(n1292) );
  INV_X1 U1296 ( .A(n632), .ZN(n1293) );
  INV_X1 U1297 ( .A(n632), .ZN(n1294) );
  INV_X1 U1298 ( .A(n4187), .ZN(n1295) );
  INV_X1 U1299 ( .A(n1295), .ZN(n1296) );
  INV_X1 U1300 ( .A(n1295), .ZN(n1297) );
  INV_X1 U1301 ( .A(n3826), .ZN(n1298) );
  INV_X1 U1302 ( .A(n3828), .ZN(n1299) );
  INV_X1 U1303 ( .A(n3822), .ZN(n13001) );
  INV_X1 U1304 ( .A(n3824), .ZN(n1301) );
  INV_X1 U1305 ( .A(n3818), .ZN(n1302) );
  INV_X1 U1306 ( .A(n38201), .ZN(n1303) );
  INV_X1 U1307 ( .A(n3814), .ZN(n1304) );
  INV_X1 U1308 ( .A(n3816), .ZN(n1305) );
  INV_X1 U1309 ( .A(n38101), .ZN(n1306) );
  INV_X1 U1310 ( .A(n3812), .ZN(n1307) );
  INV_X1 U1311 ( .A(n3806), .ZN(n1308) );
  INV_X1 U1312 ( .A(n3808), .ZN(n1309) );
  INV_X1 U1313 ( .A(n3802), .ZN(n13101) );
  INV_X1 U1314 ( .A(n3804), .ZN(n1311) );
  INV_X1 U1315 ( .A(n3797), .ZN(n1312) );
  INV_X1 U1316 ( .A(n38001), .ZN(n1313) );
  INV_X1 U1317 ( .A(n633), .ZN(n1314) );
  INV_X1 U1318 ( .A(n634), .ZN(n1315) );
  INV_X1 U1319 ( .A(n635), .ZN(n1316) );
  INV_X1 U1320 ( .A(n636), .ZN(n1317) );
  INV_X1 U1321 ( .A(n637), .ZN(n1318) );
  INV_X1 U1322 ( .A(n638), .ZN(n1319) );
  INV_X1 U1323 ( .A(n639), .ZN(n13201) );
  INV_X1 U1324 ( .A(n640), .ZN(n1321) );
  INV_X1 U1325 ( .A(n641), .ZN(n1322) );
  INV_X1 U1326 ( .A(n642), .ZN(n1323) );
  INV_X1 U1327 ( .A(n643), .ZN(n1324) );
  INV_X1 U1328 ( .A(n644), .ZN(n1325) );
  INV_X1 U1329 ( .A(n645), .ZN(n1326) );
  INV_X1 U1330 ( .A(n646), .ZN(n1327) );
  INV_X1 U1331 ( .A(n647), .ZN(n1328) );
  INV_X1 U1332 ( .A(n648), .ZN(n1329) );
  INV_X1 U1333 ( .A(n3753), .ZN(n13301) );
  INV_X1 U1334 ( .A(n3755), .ZN(n1331) );
  INV_X1 U1335 ( .A(n3749), .ZN(n1332) );
  INV_X1 U1336 ( .A(n3751), .ZN(n1333) );
  INV_X1 U1337 ( .A(n3745), .ZN(n1334) );
  INV_X1 U1338 ( .A(n3747), .ZN(n1335) );
  INV_X1 U1339 ( .A(n3741), .ZN(n1336) );
  INV_X1 U1340 ( .A(n3743), .ZN(n1337) );
  INV_X1 U1341 ( .A(n3737), .ZN(n1338) );
  INV_X1 U1342 ( .A(n3739), .ZN(n1339) );
  INV_X1 U1343 ( .A(n3733), .ZN(n13401) );
  INV_X1 U1344 ( .A(n3735), .ZN(n1341) );
  INV_X1 U1345 ( .A(n3729), .ZN(n1342) );
  INV_X1 U1346 ( .A(n3731), .ZN(n1343) );
  INV_X1 U1347 ( .A(n3724), .ZN(n1344) );
  INV_X1 U1348 ( .A(n3727), .ZN(n1345) );
  INV_X1 U1349 ( .A(n649), .ZN(n1346) );
  INV_X1 U1350 ( .A(n965), .ZN(n1347) );
  INV_X1 U1351 ( .A(n650), .ZN(n1348) );
  INV_X1 U1352 ( .A(n651), .ZN(n1349) );
  INV_X1 U1353 ( .A(n652), .ZN(n13501) );
  INV_X1 U1354 ( .A(n2927), .ZN(n1351) );
  INV_X1 U1355 ( .A(n1351), .ZN(n1352) );
  INV_X1 U1356 ( .A(n653), .ZN(n1353) );
  INV_X1 U1357 ( .A(n654), .ZN(n1354) );
  INV_X1 U1358 ( .A(n655), .ZN(n1355) );
  INV_X1 U1359 ( .A(n2936), .ZN(n1356) );
  INV_X1 U1360 ( .A(n1356), .ZN(n1357) );
  INV_X1 U1361 ( .A(n656), .ZN(n1358) );
  INV_X1 U1362 ( .A(n658), .ZN(n1359) );
  INV_X1 U1363 ( .A(n1359), .ZN(n13601) );
  INV_X1 U1364 ( .A(n658), .ZN(n1361) );
  INV_X1 U1365 ( .A(n13601), .ZN(n1362) );
  INV_X1 U1366 ( .A(n1365), .ZN(n1363) );
  INV_X1 U1367 ( .A(n660), .ZN(n1364) );
  INV_X1 U1368 ( .A(n660), .ZN(n1365) );
  INV_X1 U1369 ( .A(n661), .ZN(n1366) );
  INV_X1 U1370 ( .A(n1366), .ZN(n1367) );
  INV_X1 U1371 ( .A(n1367), .ZN(n1368) );
  INV_X1 U1372 ( .A(n661), .ZN(n1369) );
  INV_X1 U1373 ( .A(n662), .ZN(n13701) );
  INV_X1 U1374 ( .A(n2949), .ZN(n1371) );
  INV_X1 U1375 ( .A(n1371), .ZN(n1372) );
  INV_X1 U1376 ( .A(n1372), .ZN(n1373) );
  INV_X1 U1377 ( .A(n2949), .ZN(n1374) );
  INV_X1 U1378 ( .A(n1377), .ZN(n1375) );
  INV_X1 U1379 ( .A(n664), .ZN(n1376) );
  INV_X1 U1380 ( .A(n664), .ZN(n1377) );
  INV_X1 U1381 ( .A(n2953), .ZN(n1378) );
  INV_X1 U1382 ( .A(n1378), .ZN(n1379) );
  INV_X1 U1383 ( .A(n1379), .ZN(n13801) );
  INV_X1 U1384 ( .A(n2953), .ZN(n1381) );
  INV_X1 U1385 ( .A(n1384), .ZN(n1382) );
  INV_X1 U1386 ( .A(n665), .ZN(n1383) );
  INV_X1 U1387 ( .A(n665), .ZN(n1384) );
  INV_X1 U1388 ( .A(n2957), .ZN(n1385) );
  INV_X1 U1389 ( .A(n1385), .ZN(n1386) );
  INV_X1 U1390 ( .A(n1386), .ZN(n1387) );
  INV_X1 U1391 ( .A(n2957), .ZN(n1388) );
  INV_X1 U1392 ( .A(n1391), .ZN(n1389) );
  INV_X1 U1393 ( .A(n666), .ZN(n13901) );
  INV_X1 U1394 ( .A(n666), .ZN(n1391) );
  INV_X1 U1395 ( .A(n2961), .ZN(n1392) );
  INV_X1 U1396 ( .A(n1392), .ZN(n1393) );
  INV_X1 U1397 ( .A(n1393), .ZN(n1394) );
  INV_X1 U1398 ( .A(n2961), .ZN(n1395) );
  INV_X1 U1399 ( .A(n667), .ZN(n1396) );
  INV_X1 U1400 ( .A(n2965), .ZN(n1397) );
  INV_X1 U1401 ( .A(n1397), .ZN(n1398) );
  INV_X1 U1402 ( .A(n1398), .ZN(n1399) );
  INV_X1 U1403 ( .A(n2965), .ZN(n14001) );
  INV_X1 U1404 ( .A(n668), .ZN(n1401) );
  INV_X1 U1405 ( .A(n2969), .ZN(n1402) );
  INV_X1 U1406 ( .A(n1402), .ZN(n1403) );
  INV_X1 U1407 ( .A(n1403), .ZN(n1404) );
  INV_X1 U1408 ( .A(n2969), .ZN(n1405) );
  INV_X1 U1409 ( .A(n669), .ZN(n1406) );
  INV_X1 U1410 ( .A(n2973), .ZN(n1407) );
  INV_X1 U1411 ( .A(n1407), .ZN(n1408) );
  INV_X1 U1412 ( .A(n1408), .ZN(n1409) );
  INV_X1 U1413 ( .A(n2973), .ZN(n14101) );
  INV_X1 U1414 ( .A(n1413), .ZN(n1411) );
  INV_X1 U1415 ( .A(n670), .ZN(n1412) );
  INV_X1 U1416 ( .A(n670), .ZN(n1413) );
  INV_X1 U1417 ( .A(n2977), .ZN(n1414) );
  INV_X1 U1418 ( .A(n1414), .ZN(n1415) );
  INV_X1 U1419 ( .A(n1415), .ZN(n1416) );
  INV_X1 U1420 ( .A(n2977), .ZN(n1417) );
  INV_X1 U1421 ( .A(n671), .ZN(n1418) );
  INV_X1 U1422 ( .A(n2981), .ZN(n1419) );
  INV_X1 U1423 ( .A(n1419), .ZN(n14201) );
  INV_X1 U1424 ( .A(n14201), .ZN(n1421) );
  INV_X1 U1425 ( .A(n2981), .ZN(n1422) );
  INV_X1 U1426 ( .A(n1425), .ZN(n1423) );
  INV_X1 U1427 ( .A(n672), .ZN(n1424) );
  INV_X1 U1428 ( .A(n672), .ZN(n1425) );
  INV_X1 U1429 ( .A(n2985), .ZN(n1426) );
  INV_X1 U1430 ( .A(n1426), .ZN(n1427) );
  INV_X1 U1431 ( .A(n1427), .ZN(n1428) );
  INV_X1 U1432 ( .A(n2985), .ZN(n1429) );
  INV_X1 U1433 ( .A(n1432), .ZN(n14301) );
  INV_X1 U1434 ( .A(n673), .ZN(n1431) );
  INV_X1 U1435 ( .A(n673), .ZN(n1432) );
  INV_X1 U1436 ( .A(n2989), .ZN(n1433) );
  INV_X1 U1437 ( .A(n1433), .ZN(n1434) );
  INV_X1 U1438 ( .A(n1434), .ZN(n1435) );
  INV_X1 U1439 ( .A(n2989), .ZN(n1436) );
  INV_X1 U1440 ( .A(n1439), .ZN(n1437) );
  INV_X1 U1441 ( .A(n674), .ZN(n1438) );
  INV_X1 U1442 ( .A(n674), .ZN(n1439) );
  INV_X1 U1443 ( .A(n2993), .ZN(n14401) );
  INV_X1 U1444 ( .A(n14401), .ZN(n1441) );
  INV_X1 U1445 ( .A(n1441), .ZN(n1442) );
  INV_X1 U1446 ( .A(n2993), .ZN(n1443) );
  INV_X1 U1447 ( .A(n675), .ZN(n1444) );
  INV_X1 U1448 ( .A(n2997), .ZN(n1445) );
  INV_X1 U1449 ( .A(n1445), .ZN(n1446) );
  INV_X1 U1450 ( .A(n1446), .ZN(n1447) );
  INV_X1 U1451 ( .A(n2997), .ZN(n1448) );
  INV_X1 U1452 ( .A(n1451), .ZN(n1449) );
  INV_X1 U1453 ( .A(n677), .ZN(n14501) );
  INV_X1 U1454 ( .A(n677), .ZN(n1451) );
  INV_X1 U1455 ( .A(n3001), .ZN(n1452) );
  INV_X1 U1456 ( .A(n1452), .ZN(n1453) );
  INV_X1 U1457 ( .A(n1453), .ZN(n1454) );
  INV_X1 U1458 ( .A(n3001), .ZN(n1455) );
  INV_X1 U1459 ( .A(n1458), .ZN(n1456) );
  INV_X1 U1460 ( .A(n678), .ZN(n1457) );
  INV_X1 U1461 ( .A(n678), .ZN(n1458) );
  INV_X1 U1462 ( .A(n3005), .ZN(n1459) );
  INV_X1 U1463 ( .A(n1459), .ZN(n14601) );
  INV_X1 U1464 ( .A(n14601), .ZN(n1461) );
  INV_X1 U1465 ( .A(n3005), .ZN(n1462) );
  INV_X1 U1466 ( .A(n679), .ZN(n1463) );
  INV_X1 U1467 ( .A(n1463), .ZN(n1464) );
  INV_X1 U1468 ( .A(n679), .ZN(n1465) );
  INV_X1 U1469 ( .A(n1464), .ZN(n1466) );
  INV_X1 U1470 ( .A(n680), .ZN(n1467) );
  INV_X1 U1471 ( .A(n681), .ZN(n1468) );
  INV_X1 U1472 ( .A(n681), .ZN(n1469) );
  INV_X1 U1473 ( .A(n682), .ZN(n14701) );
  INV_X1 U1474 ( .A(n682), .ZN(n1471) );
  INV_X1 U1475 ( .A(n2698), .ZN(n1472) );
  INV_X1 U1476 ( .A(n3709), .ZN(n1473) );
  INV_X1 U1477 ( .A(n3445), .ZN(n1474) );
  INV_X1 U1478 ( .A(n1474), .ZN(n1475) );
  INV_X1 U1479 ( .A(n1474), .ZN(n1476) );
  INV_X1 U1480 ( .A(n684), .ZN(n1477) );
  INV_X1 U1481 ( .A(n685), .ZN(n1478) );
  INV_X1 U1482 ( .A(n685), .ZN(n1479) );
  INV_X1 U1483 ( .A(n686), .ZN(n14801) );
  INV_X1 U1484 ( .A(n687), .ZN(n1481) );
  INV_X1 U1485 ( .A(n687), .ZN(n1482) );
  INV_X1 U1486 ( .A(n688), .ZN(n1483) );
  INV_X1 U1487 ( .A(n689), .ZN(n1484) );
  INV_X1 U1488 ( .A(n689), .ZN(n1485) );
  INV_X1 U1489 ( .A(n690), .ZN(n1486) );
  INV_X1 U1490 ( .A(n691), .ZN(n1487) );
  INV_X1 U1491 ( .A(n691), .ZN(n1488) );
  INV_X1 U1492 ( .A(n692), .ZN(n1489) );
  INV_X1 U1493 ( .A(n692), .ZN(n14901) );
  INV_X1 U1494 ( .A(n2029), .ZN(n1491) );
  INV_X1 U1495 ( .A(n1491), .ZN(n1492) );
  INV_X1 U1496 ( .A(n1491), .ZN(n1493) );
  INV_X1 U1497 ( .A(n3022), .ZN(n1494) );
  INV_X1 U1498 ( .A(n1494), .ZN(n1495) );
  INV_X1 U1499 ( .A(n1494), .ZN(n1496) );
  INV_X1 U1500 ( .A(n693), .ZN(n1497) );
  INV_X1 U1501 ( .A(n694), .ZN(n1498) );
  INV_X1 U1502 ( .A(n694), .ZN(n1499) );
  INV_X1 U1503 ( .A(n695), .ZN(n15001) );
  INV_X1 U1504 ( .A(n696), .ZN(n1501) );
  INV_X1 U1505 ( .A(n696), .ZN(n1502) );
  INV_X1 U1506 ( .A(n697), .ZN(n1503) );
  INV_X1 U1507 ( .A(n698), .ZN(n1504) );
  INV_X1 U1508 ( .A(n698), .ZN(n1505) );
  INV_X1 U1509 ( .A(n42701), .ZN(n1506) );
  INV_X1 U1510 ( .A(n1506), .ZN(n1507) );
  INV_X1 U1511 ( .A(n1506), .ZN(n1508) );
  INV_X1 U1512 ( .A(n3311), .ZN(n1509) );
  INV_X1 U1513 ( .A(n1509), .ZN(n15101) );
  INV_X1 U1514 ( .A(n1509), .ZN(n1511) );
  INV_X1 U1515 ( .A(n3313), .ZN(n1512) );
  INV_X1 U1516 ( .A(n1512), .ZN(n1513) );
  INV_X1 U1517 ( .A(n1512), .ZN(n1514) );
  INV_X1 U1518 ( .A(n4338), .ZN(n1515) );
  INV_X1 U1519 ( .A(n1515), .ZN(n1516) );
  INV_X1 U1520 ( .A(n1515), .ZN(n1517) );
  INV_X1 U1521 ( .A(n2927), .ZN(n1518) );
  INV_X1 U1522 ( .A(n1518), .ZN(n1519) );
  INV_X1 U1523 ( .A(n1518), .ZN(n15201) );
  INV_X1 U1524 ( .A(n3321), .ZN(n1521) );
  INV_X1 U1525 ( .A(n1521), .ZN(n1522) );
  INV_X1 U1526 ( .A(n1521), .ZN(n1523) );
  INV_X1 U1527 ( .A(n699), .ZN(n1524) );
  INV_X1 U1528 ( .A(n699), .ZN(n1525) );
  INV_X1 U1529 ( .A(N102), .ZN(n1526) );
  INV_X1 U1530 ( .A(n1526), .ZN(n1527) );
  INV_X1 U1531 ( .A(n1526), .ZN(n1528) );
  INV_X1 U1532 ( .A(n700), .ZN(n1529) );
  INV_X1 U1533 ( .A(n700), .ZN(n15301) );
  INV_X1 U1534 ( .A(N100), .ZN(n1531) );
  INV_X1 U1535 ( .A(n1531), .ZN(n1532) );
  INV_X1 U1536 ( .A(n1531), .ZN(n1533) );
  INV_X1 U1537 ( .A(n34301), .ZN(n1534) );
  INV_X1 U1538 ( .A(n1534), .ZN(n1535) );
  INV_X1 U1539 ( .A(n1534), .ZN(n1536) );
  INV_X1 U1540 ( .A(n3431), .ZN(n1537) );
  INV_X1 U1541 ( .A(n576), .ZN(n1538) );
  INV_X1 U1542 ( .A(n701), .ZN(n15390) );
  INV_X1 U1543 ( .A(n701), .ZN(n15401) );
  INV_X1 U1544 ( .A(n702), .ZN(n1541) );
  INV_X1 U1545 ( .A(n702), .ZN(n1542) );
  INV_X1 U1546 ( .A(n703), .ZN(n1543) );
  INV_X1 U1547 ( .A(n703), .ZN(n1544) );
  INV_X1 U1548 ( .A(n704), .ZN(n1545) );
  INV_X1 U1549 ( .A(n704), .ZN(n1546) );
  INV_X1 U1550 ( .A(n705), .ZN(n15470) );
  INV_X1 U1551 ( .A(n705), .ZN(n15480) );
  INV_X1 U1552 ( .A(n706), .ZN(n15490) );
  INV_X1 U1553 ( .A(n706), .ZN(n15500) );
  INV_X1 U1554 ( .A(n707), .ZN(n15511) );
  INV_X1 U1555 ( .A(n707), .ZN(n15520) );
  INV_X1 U1556 ( .A(n708), .ZN(n15530) );
  INV_X1 U1557 ( .A(n708), .ZN(n15540) );
  INV_X1 U1558 ( .A(n709), .ZN(n15550) );
  INV_X1 U1559 ( .A(n709), .ZN(n15560) );
  INV_X1 U1560 ( .A(n710), .ZN(n15570) );
  INV_X1 U1561 ( .A(n710), .ZN(n15580) );
  INV_X1 U1562 ( .A(n711), .ZN(n15590) );
  INV_X1 U1563 ( .A(n711), .ZN(n15600) );
  INV_X1 U1564 ( .A(n712), .ZN(n15610) );
  INV_X1 U1565 ( .A(n712), .ZN(n15620) );
  INV_X1 U1566 ( .A(n713), .ZN(n15631) );
  INV_X1 U1567 ( .A(n713), .ZN(n1564) );
  INV_X1 U1568 ( .A(n3719), .ZN(n1565) );
  INV_X1 U1569 ( .A(n1206), .ZN(n1566) );
  INV_X1 U1570 ( .A(n714), .ZN(n1567) );
  INV_X1 U1571 ( .A(n714), .ZN(n1568) );
  INV_X1 U1572 ( .A(n715), .ZN(n1569) );
  INV_X1 U1573 ( .A(n715), .ZN(n15701) );
  INV_X1 U1574 ( .A(n716), .ZN(n1571) );
  INV_X1 U1575 ( .A(n716), .ZN(n1572) );
  INV_X1 U1576 ( .A(n717), .ZN(n1573) );
  INV_X1 U1577 ( .A(n717), .ZN(n1574) );
  INV_X1 U1578 ( .A(n3288), .ZN(n1575) );
  INV_X1 U1579 ( .A(n1575), .ZN(n1576) );
  INV_X1 U1580 ( .A(n1575), .ZN(n1577) );
  INV_X1 U1581 ( .A(n3279), .ZN(n1578) );
  INV_X1 U1582 ( .A(n1578), .ZN(n1579) );
  INV_X1 U1583 ( .A(n1578), .ZN(n15801) );
  INV_X1 U1584 ( .A(n3312), .ZN(n15810) );
  INV_X1 U1585 ( .A(n15810), .ZN(n15820) );
  INV_X1 U1586 ( .A(n15810), .ZN(n15830) );
  INV_X1 U1587 ( .A(n718), .ZN(n15840) );
  INV_X1 U1588 ( .A(n718), .ZN(n15850) );
  INV_X1 U1589 ( .A(n3284), .ZN(n15860) );
  INV_X1 U1590 ( .A(n15860), .ZN(n15870) );
  INV_X1 U1591 ( .A(n15860), .ZN(n15880) );
  INV_X1 U1592 ( .A(n3285), .ZN(n15890) );
  INV_X1 U1593 ( .A(n15890), .ZN(n15900) );
  INV_X1 U1594 ( .A(n15890), .ZN(n15910) );
  INV_X1 U1595 ( .A(n3288), .ZN(n15920) );
  INV_X1 U1596 ( .A(n15920), .ZN(n15930) );
  INV_X1 U1597 ( .A(n15920), .ZN(n15940) );
  INV_X1 U1598 ( .A(n3287), .ZN(n15950) );
  INV_X1 U1599 ( .A(n15950), .ZN(n15960) );
  INV_X1 U1600 ( .A(n15950), .ZN(n15971) );
  INV_X1 U1601 ( .A(n2539), .ZN(n1598) );
  INV_X1 U1602 ( .A(n1598), .ZN(n1599) );
  INV_X1 U1603 ( .A(n1598), .ZN(n16001) );
  INV_X1 U1604 ( .A(n3292), .ZN(n1601) );
  INV_X1 U1605 ( .A(n1601), .ZN(n1602) );
  INV_X1 U1606 ( .A(n1601), .ZN(n1603) );
  INV_X1 U1607 ( .A(n3294), .ZN(n1604) );
  INV_X1 U1608 ( .A(n1604), .ZN(n1605) );
  INV_X1 U1609 ( .A(n1604), .ZN(n1606) );
  INV_X1 U1610 ( .A(n3285), .ZN(n1607) );
  INV_X1 U1611 ( .A(n1607), .ZN(n1608) );
  INV_X1 U1612 ( .A(n1607), .ZN(n1609) );
  INV_X1 U1613 ( .A(n3297), .ZN(n16101) );
  INV_X1 U1614 ( .A(n16101), .ZN(n1611) );
  INV_X1 U1615 ( .A(n16101), .ZN(n1612) );
  INV_X1 U1616 ( .A(n3298), .ZN(n1613) );
  INV_X1 U1617 ( .A(n1613), .ZN(n1614) );
  INV_X1 U1618 ( .A(n1613), .ZN(n1615) );
  INV_X1 U1619 ( .A(n33001), .ZN(n1616) );
  INV_X1 U1620 ( .A(n1616), .ZN(n1617) );
  INV_X1 U1621 ( .A(n1616), .ZN(n1618) );
  INV_X1 U1622 ( .A(n719), .ZN(n1619) );
  INV_X1 U1623 ( .A(n720), .ZN(n16201) );
  INV_X1 U1624 ( .A(n720), .ZN(n1621) );
  INV_X1 U1625 ( .A(n721), .ZN(n1622) );
  INV_X1 U1626 ( .A(n722), .ZN(n16230) );
  INV_X1 U1627 ( .A(n722), .ZN(n16240) );
  INV_X1 U1628 ( .A(n723), .ZN(n16250) );
  INV_X1 U1629 ( .A(n724), .ZN(n16260) );
  INV_X1 U1630 ( .A(n724), .ZN(n16270) );
  INV_X1 U1631 ( .A(n725), .ZN(n16280) );
  INV_X1 U1632 ( .A(n726), .ZN(n16290) );
  INV_X1 U1633 ( .A(n726), .ZN(n16300) );
  INV_X1 U1634 ( .A(n727), .ZN(n16310) );
  INV_X1 U1635 ( .A(n728), .ZN(n16320) );
  INV_X1 U1636 ( .A(n728), .ZN(n16330) );
  INV_X1 U1637 ( .A(n729), .ZN(n16340) );
  INV_X1 U1638 ( .A(n730), .ZN(n16350) );
  INV_X1 U1639 ( .A(n730), .ZN(n16360) );
  INV_X1 U1640 ( .A(n731), .ZN(n16370) );
  INV_X1 U1641 ( .A(n732), .ZN(n16380) );
  INV_X1 U1642 ( .A(n732), .ZN(n16391) );
  INV_X1 U1643 ( .A(n733), .ZN(n16401) );
  INV_X1 U1644 ( .A(n734), .ZN(n1641) );
  INV_X1 U1645 ( .A(n734), .ZN(n1642) );
  INV_X1 U1646 ( .A(n735), .ZN(n1643) );
  INV_X1 U1647 ( .A(n736), .ZN(n1644) );
  INV_X1 U1648 ( .A(n736), .ZN(n1645) );
  INV_X1 U1649 ( .A(n737), .ZN(n1646) );
  INV_X1 U1650 ( .A(n738), .ZN(n1647) );
  INV_X1 U1651 ( .A(n738), .ZN(n1648) );
  INV_X1 U1652 ( .A(n739), .ZN(n1649) );
  INV_X1 U1653 ( .A(n740), .ZN(n16501) );
  INV_X1 U1654 ( .A(n740), .ZN(n1651) );
  INV_X1 U1655 ( .A(n741), .ZN(n1652) );
  INV_X1 U1656 ( .A(n742), .ZN(n1653) );
  INV_X1 U1657 ( .A(n742), .ZN(n1654) );
  INV_X1 U1658 ( .A(n743), .ZN(n1655) );
  INV_X1 U1659 ( .A(n744), .ZN(n1656) );
  INV_X1 U1660 ( .A(n744), .ZN(n1657) );
  INV_X1 U1661 ( .A(n745), .ZN(n1658) );
  INV_X1 U1662 ( .A(n746), .ZN(n1659) );
  INV_X1 U1663 ( .A(n746), .ZN(n16601) );
  INV_X1 U1664 ( .A(n747), .ZN(n1661) );
  INV_X1 U1665 ( .A(n748), .ZN(n1662) );
  INV_X1 U1666 ( .A(n748), .ZN(n1663) );
  INV_X1 U1667 ( .A(n749), .ZN(n1664) );
  INV_X1 U1668 ( .A(n750), .ZN(n1665) );
  INV_X1 U1669 ( .A(n750), .ZN(n1666) );
  INV_X1 U1670 ( .A(n751), .ZN(n1667) );
  INV_X1 U1671 ( .A(n752), .ZN(n1668) );
  INV_X1 U1672 ( .A(n752), .ZN(n1669) );
  INV_X1 U1673 ( .A(n753), .ZN(n16701) );
  INV_X1 U1674 ( .A(n754), .ZN(n1671) );
  INV_X1 U1675 ( .A(n754), .ZN(n1672) );
  INV_X1 U1676 ( .A(n4131), .ZN(n1673) );
  INV_X1 U1677 ( .A(n755), .ZN(n1674) );
  INV_X1 U1678 ( .A(n755), .ZN(n1675) );
  INV_X1 U1679 ( .A(n756), .ZN(n1676) );
  INV_X1 U1680 ( .A(n757), .ZN(n1677) );
  INV_X1 U1681 ( .A(n757), .ZN(n1678) );
  INV_X1 U1682 ( .A(n758), .ZN(n1679) );
  INV_X1 U1683 ( .A(n759), .ZN(n16801) );
  INV_X1 U1684 ( .A(n759), .ZN(n1681) );
  INV_X1 U1685 ( .A(n760), .ZN(n1682) );
  INV_X1 U1686 ( .A(n761), .ZN(n1683) );
  INV_X1 U1687 ( .A(n761), .ZN(n1684) );
  INV_X1 U1688 ( .A(n762), .ZN(n1685) );
  INV_X1 U1689 ( .A(n763), .ZN(n1686) );
  INV_X1 U1690 ( .A(n763), .ZN(n1687) );
  INV_X1 U1691 ( .A(n764), .ZN(n1688) );
  INV_X1 U1692 ( .A(n765), .ZN(n1689) );
  INV_X1 U1693 ( .A(n765), .ZN(n16901) );
  INV_X1 U1694 ( .A(n766), .ZN(n1691) );
  INV_X1 U1695 ( .A(n767), .ZN(n1692) );
  INV_X1 U1696 ( .A(n767), .ZN(n1693) );
  INV_X1 U1697 ( .A(n768), .ZN(n1694) );
  INV_X1 U1698 ( .A(n769), .ZN(n1695) );
  INV_X1 U1699 ( .A(n769), .ZN(n1696) );
  INV_X1 U1700 ( .A(n770), .ZN(n1697) );
  INV_X1 U1701 ( .A(n771), .ZN(n1698) );
  INV_X1 U1702 ( .A(n771), .ZN(n1699) );
  INV_X1 U1703 ( .A(n772), .ZN(n17001) );
  INV_X1 U1704 ( .A(n773), .ZN(n1701) );
  INV_X1 U1705 ( .A(n773), .ZN(n1702) );
  INV_X1 U1706 ( .A(n774), .ZN(n1703) );
  INV_X1 U1707 ( .A(n775), .ZN(n1704) );
  INV_X1 U1708 ( .A(n775), .ZN(n1705) );
  INV_X1 U1709 ( .A(n776), .ZN(n1706) );
  INV_X1 U1710 ( .A(n777), .ZN(n1707) );
  INV_X1 U1711 ( .A(n777), .ZN(n1708) );
  INV_X1 U1712 ( .A(n778), .ZN(n1709) );
  INV_X1 U1713 ( .A(n779), .ZN(n17101) );
  INV_X1 U1714 ( .A(n779), .ZN(n1711) );
  INV_X1 U1715 ( .A(n3353), .ZN(n1712) );
  INV_X1 U1716 ( .A(n1712), .ZN(n1713) );
  INV_X1 U1717 ( .A(n1712), .ZN(n1714) );
  INV_X1 U1718 ( .A(n3353), .ZN(n1715) );
  INV_X1 U1719 ( .A(n1713), .ZN(n1716) );
  INV_X1 U1720 ( .A(n3356), .ZN(n1717) );
  INV_X1 U1721 ( .A(n1717), .ZN(n1718) );
  INV_X1 U1722 ( .A(n3356), .ZN(n1719) );
  INV_X1 U1723 ( .A(n1718), .ZN(n17201) );
  INV_X1 U1724 ( .A(n780), .ZN(n1721) );
  INV_X1 U1725 ( .A(n781), .ZN(n1722) );
  INV_X1 U1726 ( .A(n781), .ZN(n1723) );
  INV_X1 U1727 ( .A(n782), .ZN(n1724) );
  INV_X1 U1728 ( .A(n783), .ZN(n1725) );
  INV_X1 U1729 ( .A(n783), .ZN(n1726) );
  INV_X1 U1730 ( .A(n784), .ZN(n1727) );
  INV_X1 U1731 ( .A(n785), .ZN(n1728) );
  INV_X1 U1732 ( .A(n785), .ZN(n1729) );
  INV_X1 U1733 ( .A(n786), .ZN(n17301) );
  INV_X1 U1734 ( .A(n787), .ZN(n1731) );
  INV_X1 U1735 ( .A(n787), .ZN(n1732) );
  INV_X1 U1736 ( .A(n4201), .ZN(n1733) );
  INV_X1 U1737 ( .A(n788), .ZN(n1734) );
  INV_X1 U1738 ( .A(n788), .ZN(n1735) );
  INV_X1 U1739 ( .A(n789), .ZN(n1736) );
  INV_X1 U1740 ( .A(n790), .ZN(n1737) );
  INV_X1 U1741 ( .A(n790), .ZN(n1738) );
  INV_X1 U1742 ( .A(n791), .ZN(n1739) );
  INV_X1 U1743 ( .A(n792), .ZN(n17401) );
  INV_X1 U1744 ( .A(n792), .ZN(n1741) );
  INV_X1 U1745 ( .A(n1131), .ZN(n1742) );
  INV_X1 U1746 ( .A(n1742), .ZN(n1743) );
  INV_X1 U1747 ( .A(n1104), .ZN(n1744) );
  INV_X1 U1748 ( .A(n1744), .ZN(n1745) );
  INV_X1 U1749 ( .A(n1744), .ZN(n1746) );
  INV_X1 U1750 ( .A(n3367), .ZN(n1747) );
  INV_X1 U1751 ( .A(n1747), .ZN(n1748) );
  INV_X1 U1752 ( .A(n3367), .ZN(n1749) );
  INV_X1 U1753 ( .A(n1748), .ZN(n17501) );
  INV_X1 U1754 ( .A(n793), .ZN(n1751) );
  INV_X1 U1755 ( .A(n1106), .ZN(n1752) );
  INV_X1 U1756 ( .A(n1752), .ZN(n1753) );
  INV_X1 U1757 ( .A(n1752), .ZN(n1754) );
  INV_X1 U1758 ( .A(n794), .ZN(n1755) );
  INV_X1 U1759 ( .A(n1107), .ZN(n1756) );
  INV_X1 U1760 ( .A(n1756), .ZN(n1757) );
  INV_X1 U1761 ( .A(n1756), .ZN(n1758) );
  INV_X1 U1762 ( .A(n795), .ZN(n1759) );
  INV_X1 U1763 ( .A(n796), .ZN(n17601) );
  INV_X1 U1764 ( .A(n2936), .ZN(n1761) );
  INV_X1 U1765 ( .A(n1761), .ZN(n1762) );
  INV_X1 U1766 ( .A(n3387), .ZN(n1763) );
  INV_X1 U1767 ( .A(n1763), .ZN(n1764) );
  INV_X1 U1768 ( .A(n3387), .ZN(n1765) );
  INV_X1 U1769 ( .A(n1765), .ZN(n1766) );
  INV_X1 U1770 ( .A(n797), .ZN(n1767) );
  INV_X1 U1771 ( .A(n797), .ZN(n1768) );
  INV_X1 U1772 ( .A(n798), .ZN(n1769) );
  INV_X1 U1773 ( .A(n798), .ZN(n17701) );
  INV_X1 U1774 ( .A(n799), .ZN(n1771) );
  INV_X1 U1775 ( .A(n799), .ZN(n1772) );
  INV_X1 U1776 ( .A(n800), .ZN(n1773) );
  INV_X1 U1777 ( .A(n801), .ZN(n1774) );
  INV_X1 U1778 ( .A(n802), .ZN(n1775) );
  INV_X1 U1779 ( .A(n802), .ZN(n1776) );
  INV_X1 U1780 ( .A(n1775), .ZN(n1777) );
  INV_X1 U1781 ( .A(n1777), .ZN(n1778) );
  INV_X1 U1782 ( .A(n1777), .ZN(n1779) );
  INV_X1 U1783 ( .A(n803), .ZN(n17801) );
  INV_X1 U1784 ( .A(n803), .ZN(n1781) );
  INV_X1 U1785 ( .A(n17801), .ZN(n1782) );
  INV_X1 U1786 ( .A(n1782), .ZN(n1783) );
  INV_X1 U1787 ( .A(n1782), .ZN(n1784) );
  INV_X1 U1788 ( .A(n804), .ZN(n1785) );
  INV_X1 U1789 ( .A(n805), .ZN(n1786) );
  INV_X1 U1790 ( .A(n805), .ZN(n1787) );
  INV_X1 U1791 ( .A(n1786), .ZN(n1788) );
  INV_X1 U1792 ( .A(n1788), .ZN(n1789) );
  INV_X1 U1793 ( .A(n1788), .ZN(n17901) );
  INV_X1 U1794 ( .A(n806), .ZN(n1791) );
  INV_X1 U1795 ( .A(n806), .ZN(n1792) );
  INV_X1 U1796 ( .A(n1127), .ZN(n1793) );
  INV_X1 U1797 ( .A(n1793), .ZN(n1794) );
  INV_X1 U1798 ( .A(n3463), .ZN(n1795) );
  INV_X1 U1799 ( .A(n3463), .ZN(n1796) );
  INV_X1 U1800 ( .A(n807), .ZN(n1797) );
  INV_X1 U1801 ( .A(n808), .ZN(n1798) );
  INV_X1 U1802 ( .A(n808), .ZN(n1799) );
  INV_X1 U1803 ( .A(n4606), .ZN(n18001) );
  INV_X1 U1804 ( .A(n826), .ZN(n1801) );
  INV_X1 U1805 ( .A(n826), .ZN(n1802) );
  INV_X1 U1806 ( .A(n827), .ZN(n1803) );
  INV_X1 U1807 ( .A(n827), .ZN(n1804) );
  INV_X1 U1808 ( .A(n841), .ZN(n1805) );
  INV_X1 U1809 ( .A(n1805), .ZN(n1806) );
  INV_X1 U1810 ( .A(n1805), .ZN(n1807) );
  INV_X1 U1811 ( .A(n840), .ZN(n1808) );
  INV_X1 U1812 ( .A(n1808), .ZN(n1809) );
  INV_X1 U1813 ( .A(n1808), .ZN(n18101) );
  INV_X1 U1814 ( .A(n841), .ZN(n1811) );
  INV_X1 U1815 ( .A(n1811), .ZN(n1812) );
  INV_X1 U1816 ( .A(n1811), .ZN(n1813) );
  INV_X1 U1817 ( .A(n4021), .ZN(n1814) );
  INV_X1 U1818 ( .A(n1814), .ZN(n1815) );
  INV_X1 U1819 ( .A(n1814), .ZN(n1816) );
  CLKBUF_X1 U1820 ( .A(n1818), .Z(n1817) );
  CLKBUF_X1 U1821 ( .A(n4101), .Z(n1818) );
  INV_X1 U1822 ( .A(n16201), .ZN(n1819) );
  INV_X1 U1823 ( .A(n1819), .ZN(n18201) );
  INV_X1 U1824 ( .A(n1819), .ZN(n1821) );
  INV_X1 U1825 ( .A(n1818), .ZN(n1822) );
  INV_X1 U1826 ( .A(n1822), .ZN(n1823) );
  INV_X1 U1827 ( .A(n1822), .ZN(n1824) );
  CLKBUF_X1 U1828 ( .A(n1826), .Z(n1825) );
  CLKBUF_X1 U1829 ( .A(n39701), .Z(n1826) );
  INV_X1 U1830 ( .A(n16230), .ZN(n1827) );
  INV_X1 U1831 ( .A(n1827), .ZN(n1828) );
  INV_X1 U1832 ( .A(n1827), .ZN(n1829) );
  INV_X1 U1833 ( .A(n1826), .ZN(n18301) );
  INV_X1 U1834 ( .A(n18301), .ZN(n1831) );
  INV_X1 U1835 ( .A(n18301), .ZN(n1832) );
  CLKBUF_X1 U1836 ( .A(n1834), .Z(n1833) );
  CLKBUF_X1 U1837 ( .A(n4002), .Z(n1834) );
  INV_X1 U1838 ( .A(n16260), .ZN(n1835) );
  INV_X1 U1839 ( .A(n1835), .ZN(n1836) );
  INV_X1 U1840 ( .A(n1835), .ZN(n1837) );
  INV_X1 U1841 ( .A(n1834), .ZN(n1838) );
  INV_X1 U1842 ( .A(n1838), .ZN(n1839) );
  INV_X1 U1843 ( .A(n1838), .ZN(n18401) );
  CLKBUF_X1 U1844 ( .A(n1842), .Z(n1841) );
  CLKBUF_X1 U1845 ( .A(n4136), .Z(n1842) );
  INV_X1 U1846 ( .A(n16290), .ZN(n1843) );
  INV_X1 U1847 ( .A(n1843), .ZN(n1844) );
  INV_X1 U1848 ( .A(n1843), .ZN(n1845) );
  INV_X1 U1849 ( .A(n1842), .ZN(n1846) );
  INV_X1 U1850 ( .A(n1846), .ZN(n1847) );
  INV_X1 U1851 ( .A(n1846), .ZN(n1848) );
  CLKBUF_X1 U1852 ( .A(n18501), .Z(n1849) );
  CLKBUF_X1 U1853 ( .A(n4611), .Z(n18501) );
  INV_X1 U1854 ( .A(n16320), .ZN(n1851) );
  INV_X1 U1855 ( .A(n1851), .ZN(n1852) );
  INV_X1 U1856 ( .A(n1851), .ZN(n1853) );
  INV_X1 U1857 ( .A(n18501), .ZN(n1854) );
  INV_X1 U1858 ( .A(n1854), .ZN(n1855) );
  INV_X1 U1859 ( .A(n1854), .ZN(n1856) );
  CLKBUF_X1 U1860 ( .A(n1858), .Z(n1857) );
  CLKBUF_X1 U1861 ( .A(n4134), .Z(n1858) );
  INV_X1 U1862 ( .A(n16350), .ZN(n1859) );
  INV_X1 U1863 ( .A(n1859), .ZN(n18601) );
  INV_X1 U1864 ( .A(n1859), .ZN(n1861) );
  INV_X1 U1865 ( .A(n1858), .ZN(n1862) );
  INV_X1 U1866 ( .A(n1862), .ZN(n1863) );
  INV_X1 U1867 ( .A(n1862), .ZN(n1864) );
  CLKBUF_X1 U1868 ( .A(n1866), .Z(n1865) );
  CLKBUF_X1 U1869 ( .A(n4135), .Z(n1866) );
  INV_X1 U1870 ( .A(n16380), .ZN(n1867) );
  INV_X1 U1871 ( .A(n1867), .ZN(n1868) );
  INV_X1 U1872 ( .A(n1867), .ZN(n1869) );
  INV_X1 U1873 ( .A(n1866), .ZN(n18701) );
  INV_X1 U1874 ( .A(n18701), .ZN(n1871) );
  INV_X1 U1875 ( .A(n18701), .ZN(n1872) );
  CLKBUF_X1 U1876 ( .A(n1874), .Z(n1873) );
  CLKBUF_X1 U1877 ( .A(n41001), .Z(n1874) );
  INV_X1 U1878 ( .A(n1641), .ZN(n1875) );
  INV_X1 U1879 ( .A(n1875), .ZN(n1876) );
  INV_X1 U1880 ( .A(n1875), .ZN(n1877) );
  INV_X1 U1881 ( .A(n1874), .ZN(n1878) );
  INV_X1 U1882 ( .A(n1878), .ZN(n1879) );
  INV_X1 U1883 ( .A(n1878), .ZN(n18801) );
  CLKBUF_X1 U1884 ( .A(n1882), .Z(n1881) );
  CLKBUF_X1 U1885 ( .A(n3967), .Z(n1882) );
  INV_X1 U1886 ( .A(n1644), .ZN(n1883) );
  INV_X1 U1887 ( .A(n1883), .ZN(n1884) );
  INV_X1 U1888 ( .A(n1883), .ZN(n1885) );
  INV_X1 U1889 ( .A(n1882), .ZN(n1886) );
  INV_X1 U1890 ( .A(n1886), .ZN(n1887) );
  INV_X1 U1891 ( .A(n1886), .ZN(n1888) );
  CLKBUF_X1 U1892 ( .A(n18901), .Z(n1889) );
  CLKBUF_X1 U1893 ( .A(n4098), .Z(n18901) );
  INV_X1 U1894 ( .A(n18901), .ZN(n1891) );
  INV_X1 U1895 ( .A(n1891), .ZN(n1892) );
  INV_X1 U1896 ( .A(n1891), .ZN(n1893) );
  INV_X1 U1897 ( .A(n1647), .ZN(n1894) );
  INV_X1 U1898 ( .A(n1894), .ZN(n1895) );
  INV_X1 U1899 ( .A(n1894), .ZN(n1896) );
  CLKBUF_X1 U1900 ( .A(n1898), .Z(n1897) );
  CLKBUF_X1 U1901 ( .A(n4137), .Z(n1898) );
  INV_X1 U1902 ( .A(n16501), .ZN(n1899) );
  INV_X1 U1903 ( .A(n1899), .ZN(n19001) );
  INV_X1 U1904 ( .A(n1899), .ZN(n1901) );
  INV_X1 U1905 ( .A(n1898), .ZN(n1902) );
  INV_X1 U1906 ( .A(n1902), .ZN(n1903) );
  INV_X1 U1907 ( .A(n1902), .ZN(n1904) );
  CLKBUF_X1 U1908 ( .A(n1906), .Z(n1905) );
  CLKBUF_X1 U1909 ( .A(n4679), .Z(n1906) );
  INV_X1 U1910 ( .A(n1653), .ZN(n1907) );
  INV_X1 U1911 ( .A(n1907), .ZN(n1908) );
  INV_X1 U1912 ( .A(n1907), .ZN(n1909) );
  INV_X1 U1913 ( .A(n1906), .ZN(n19101) );
  INV_X1 U1914 ( .A(n19101), .ZN(n1911) );
  INV_X1 U1915 ( .A(n19101), .ZN(n1912) );
  CLKBUF_X1 U1916 ( .A(n1914), .Z(n1913) );
  CLKBUF_X1 U1917 ( .A(n4127), .Z(n1914) );
  INV_X1 U1918 ( .A(n1656), .ZN(n1915) );
  INV_X1 U1919 ( .A(n1915), .ZN(n1916) );
  INV_X1 U1920 ( .A(n1915), .ZN(n1917) );
  INV_X1 U1921 ( .A(n1914), .ZN(n1918) );
  INV_X1 U1922 ( .A(n1918), .ZN(n1919) );
  INV_X1 U1923 ( .A(n1918), .ZN(n19201) );
  CLKBUF_X1 U1924 ( .A(n1922), .Z(n1921) );
  CLKBUF_X1 U1925 ( .A(n4124), .Z(n1922) );
  INV_X1 U1926 ( .A(n1659), .ZN(n1923) );
  INV_X1 U1927 ( .A(n1923), .ZN(n1924) );
  INV_X1 U1928 ( .A(n1923), .ZN(n1925) );
  INV_X1 U1929 ( .A(n1922), .ZN(n1926) );
  INV_X1 U1930 ( .A(n1926), .ZN(n1927) );
  INV_X1 U1931 ( .A(n1926), .ZN(n1928) );
  CLKBUF_X1 U1932 ( .A(n19301), .Z(n1929) );
  CLKBUF_X1 U1933 ( .A(n4123), .Z(n19301) );
  INV_X1 U1934 ( .A(n1662), .ZN(n1931) );
  INV_X1 U1935 ( .A(n1931), .ZN(n1932) );
  INV_X1 U1936 ( .A(n1931), .ZN(n1933) );
  INV_X1 U1937 ( .A(n19301), .ZN(n1934) );
  INV_X1 U1938 ( .A(n1934), .ZN(n1935) );
  INV_X1 U1939 ( .A(n1934), .ZN(n1936) );
  CLKBUF_X1 U1940 ( .A(n1938), .Z(n1937) );
  CLKBUF_X1 U1941 ( .A(n4126), .Z(n1938) );
  OAI21_X1 U1942 ( .B1(n4129), .B2(n41301), .A(n16001), .ZN(n4126) );
  INV_X1 U1943 ( .A(n1665), .ZN(n1939) );
  INV_X1 U1944 ( .A(n1939), .ZN(n19401) );
  INV_X1 U1945 ( .A(n1939), .ZN(n1941) );
  INV_X1 U1946 ( .A(n1938), .ZN(n1942) );
  INV_X1 U1947 ( .A(n1942), .ZN(n1943) );
  INV_X1 U1948 ( .A(n1942), .ZN(n1944) );
  CLKBUF_X1 U1949 ( .A(n1946), .Z(n1945) );
  CLKBUF_X1 U1950 ( .A(n4041), .Z(n1946) );
  OAI21_X1 U1951 ( .B1(n1797), .B2(n3438), .A(n1251), .ZN(n4041) );
  INV_X1 U1952 ( .A(n1946), .ZN(n1947) );
  INV_X1 U1953 ( .A(n1947), .ZN(n1948) );
  INV_X1 U1954 ( .A(n1947), .ZN(n1949) );
  INV_X1 U1955 ( .A(n1668), .ZN(n19501) );
  INV_X1 U1956 ( .A(n19501), .ZN(n1951) );
  INV_X1 U1957 ( .A(n19501), .ZN(n1952) );
  CLKBUF_X1 U1958 ( .A(n1954), .Z(n1953) );
  CLKBUF_X1 U1959 ( .A(n4122), .Z(n1954) );
  OAI21_X1 U1960 ( .B1(n3214), .B2(n4094), .A(n4125), .ZN(n4122) );
  INV_X1 U1961 ( .A(n1671), .ZN(n1955) );
  INV_X1 U1962 ( .A(n1955), .ZN(n1956) );
  INV_X1 U1963 ( .A(n1955), .ZN(n1957) );
  INV_X1 U1964 ( .A(n1954), .ZN(n1958) );
  INV_X1 U1965 ( .A(n1958), .ZN(n1959) );
  INV_X1 U1966 ( .A(n1958), .ZN(n19601) );
  CLKBUF_X1 U1967 ( .A(n1124), .Z(n1961) );
  OAI21_X1 U1968 ( .B1(n4191), .B2(n3435), .A(n2034), .ZN(n4131) );
  INV_X1 U1969 ( .A(n1674), .ZN(n1962) );
  INV_X1 U1970 ( .A(n1962), .ZN(n1963) );
  INV_X1 U1971 ( .A(n1962), .ZN(n1964) );
  INV_X1 U1972 ( .A(n828), .ZN(n1965) );
  INV_X1 U1973 ( .A(n828), .ZN(n1966) );
  CLKBUF_X1 U1974 ( .A(n1968), .Z(n1967) );
  CLKBUF_X1 U1975 ( .A(n4194), .Z(n1968) );
  INV_X1 U1976 ( .A(n1968), .ZN(n1969) );
  INV_X1 U1977 ( .A(n1969), .ZN(n19701) );
  INV_X1 U1978 ( .A(n1969), .ZN(n1971) );
  CLKBUF_X1 U1979 ( .A(n1973), .Z(n1972) );
  CLKBUF_X1 U1980 ( .A(n4607), .Z(n1973) );
  INV_X1 U1981 ( .A(n1973), .ZN(n1974) );
  INV_X1 U1982 ( .A(n1974), .ZN(n1975) );
  INV_X1 U1983 ( .A(n1974), .ZN(n1976) );
  CLKBUF_X1 U1984 ( .A(n1978), .Z(n1977) );
  CLKBUF_X1 U1985 ( .A(n44701), .Z(n1978) );
  INV_X1 U1986 ( .A(n1978), .ZN(n1979) );
  INV_X1 U1987 ( .A(n1979), .ZN(n19801) );
  INV_X1 U1988 ( .A(n1979), .ZN(n1981) );
  CLKBUF_X1 U1989 ( .A(n1983), .Z(n1982) );
  CLKBUF_X1 U1990 ( .A(n4539), .Z(n1983) );
  INV_X1 U1991 ( .A(n1983), .ZN(n1984) );
  INV_X1 U1992 ( .A(n1984), .ZN(n1985) );
  INV_X1 U1993 ( .A(n1984), .ZN(n1986) );
  CLKBUF_X1 U1994 ( .A(n1988), .Z(n1987) );
  CLKBUF_X1 U1995 ( .A(n4334), .Z(n1988) );
  INV_X1 U1996 ( .A(n1988), .ZN(n1989) );
  INV_X1 U1997 ( .A(n1989), .ZN(n19901) );
  INV_X1 U1998 ( .A(n1989), .ZN(n1991) );
  CLKBUF_X1 U1999 ( .A(n1993), .Z(n1992) );
  CLKBUF_X1 U2000 ( .A(n4404), .Z(n1993) );
  INV_X1 U2001 ( .A(n1993), .ZN(n1994) );
  INV_X1 U2002 ( .A(n1994), .ZN(n1995) );
  INV_X1 U2003 ( .A(n1994), .ZN(n1996) );
  CLKBUF_X1 U2004 ( .A(n1998), .Z(n1997) );
  CLKBUF_X1 U2005 ( .A(n4192), .Z(n1998) );
  INV_X1 U2006 ( .A(n1998), .ZN(n1999) );
  INV_X1 U2007 ( .A(n1999), .ZN(n20001) );
  INV_X1 U2008 ( .A(n1999), .ZN(n2001) );
  CLKBUF_X1 U2009 ( .A(n2003), .Z(n2002) );
  CLKBUF_X1 U2010 ( .A(n4265), .Z(n2003) );
  INV_X1 U2011 ( .A(n2003), .ZN(n2004) );
  INV_X1 U2012 ( .A(n2004), .ZN(n2005) );
  INV_X1 U2013 ( .A(n2004), .ZN(n2006) );
  CLKBUF_X1 U2014 ( .A(n2008), .Z(n2007) );
  CLKBUF_X1 U2015 ( .A(n3799), .Z(n2008) );
  INV_X1 U2016 ( .A(n2008), .ZN(n2009) );
  INV_X1 U2017 ( .A(n2009), .ZN(n20101) );
  INV_X1 U2018 ( .A(n2009), .ZN(n2011) );
  CLKBUF_X1 U2019 ( .A(n2013), .Z(n2012) );
  CLKBUF_X1 U2020 ( .A(n3835), .Z(n2013) );
  INV_X1 U2021 ( .A(n2013), .ZN(n2014) );
  INV_X1 U2022 ( .A(n2014), .ZN(n2015) );
  INV_X1 U2023 ( .A(n2014), .ZN(n2016) );
  CLKBUF_X1 U2024 ( .A(n2018), .Z(n2017) );
  CLKBUF_X1 U2025 ( .A(n3726), .Z(n2018) );
  INV_X1 U2026 ( .A(n2018), .ZN(n2019) );
  INV_X1 U2027 ( .A(n2019), .ZN(n20201) );
  INV_X1 U2028 ( .A(n2019), .ZN(n2021) );
  CLKBUF_X1 U2029 ( .A(n2023), .Z(n2022) );
  CLKBUF_X1 U2030 ( .A(n3764), .Z(n2023) );
  INV_X1 U2031 ( .A(n2023), .ZN(n2024) );
  INV_X1 U2032 ( .A(n2024), .ZN(n2025) );
  INV_X1 U2033 ( .A(n2024), .ZN(n2026) );
  CLKBUF_X1 U2034 ( .A(n2028), .Z(n2027) );
  CLKBUF_X1 U2035 ( .A(n4267), .Z(n2028) );
  INV_X1 U2036 ( .A(n2028), .ZN(n2029) );
  INV_X1 U2037 ( .A(n1135), .ZN(n20301) );
  CLKBUF_X1 U2038 ( .A(n2032), .Z(n2031) );
  CLKBUF_X1 U2039 ( .A(n3714), .Z(n2032) );
  NOR2_X1 U2040 ( .A1(n1803), .A2(n1532), .ZN(n3714) );
  INV_X1 U2041 ( .A(n2032), .ZN(n2033) );
  INV_X1 U2042 ( .A(n2033), .ZN(n2034) );
  INV_X1 U2043 ( .A(n2033), .ZN(n2035) );
  CLKBUF_X1 U2044 ( .A(n2037), .Z(n2036) );
  CLKBUF_X1 U2045 ( .A(n3871), .Z(n2037) );
  INV_X1 U2046 ( .A(n2037), .ZN(n2038) );
  INV_X1 U2047 ( .A(n2038), .ZN(n2039) );
  INV_X1 U2048 ( .A(n2038), .ZN(n20401) );
  CLKBUF_X1 U2049 ( .A(n2042), .Z(n2041) );
  CLKBUF_X1 U2050 ( .A(n3942), .Z(n2042) );
  INV_X1 U2051 ( .A(n2042), .ZN(n2043) );
  INV_X1 U2052 ( .A(n2043), .ZN(n2044) );
  INV_X1 U2053 ( .A(n2043), .ZN(n2045) );
  CLKBUF_X1 U2054 ( .A(n2047), .Z(n2046) );
  CLKBUF_X1 U2055 ( .A(n3907), .Z(n2047) );
  INV_X1 U2056 ( .A(n2047), .ZN(n2048) );
  INV_X1 U2057 ( .A(n2048), .ZN(n2049) );
  INV_X1 U2058 ( .A(n2048), .ZN(n20501) );
  CLKBUF_X1 U2059 ( .A(n2052), .Z(n2051) );
  CLKBUF_X1 U2060 ( .A(n4023), .Z(n2052) );
  AOI21_X1 U2061 ( .B1(n2687), .B2(n40201), .A(n3296), .ZN(n4023) );
  INV_X1 U2062 ( .A(n2052), .ZN(n2053) );
  INV_X1 U2063 ( .A(n2053), .ZN(n2054) );
  INV_X1 U2064 ( .A(n2053), .ZN(n2055) );
  CLKBUF_X1 U2065 ( .A(n2057), .Z(n2056) );
  CLKBUF_X1 U2066 ( .A(n1127), .Z(n2057) );
  INV_X1 U2067 ( .A(n2057), .ZN(n2058) );
  INV_X1 U2068 ( .A(n2058), .ZN(n2059) );
  INV_X1 U2069 ( .A(n2058), .ZN(n20601) );
  CLKBUF_X1 U2070 ( .A(n2062), .Z(n2061) );
  CLKBUF_X1 U2071 ( .A(n4043), .Z(n2062) );
  OAI21_X1 U2072 ( .B1(n3273), .B2(n3439), .A(n17201), .ZN(n4043) );
  INV_X1 U2073 ( .A(n2062), .ZN(n2063) );
  INV_X1 U2074 ( .A(n2063), .ZN(n2064) );
  INV_X1 U2075 ( .A(n2063), .ZN(n2065) );
  CLKBUF_X1 U2076 ( .A(n2067), .Z(n2066) );
  CLKBUF_X1 U2077 ( .A(n4097), .Z(n2067) );
  OAI21_X1 U2078 ( .B1(n920), .B2(n3435), .A(n2786), .ZN(n4097) );
  INV_X1 U2079 ( .A(n2067), .ZN(n2068) );
  INV_X1 U2080 ( .A(n2068), .ZN(n2069) );
  INV_X1 U2081 ( .A(n2068), .ZN(n20701) );
  CLKBUF_X1 U2082 ( .A(n4142), .Z(n2071) );
  CLKBUF_X1 U2083 ( .A(n2073), .Z(n2072) );
  CLKBUF_X1 U2084 ( .A(n3718), .Z(n2073) );
  INV_X1 U2085 ( .A(n1108), .ZN(n2074) );
  INV_X1 U2086 ( .A(n2074), .ZN(n2075) );
  INV_X1 U2087 ( .A(n2074), .ZN(n2076) );
  INV_X1 U2088 ( .A(n3374), .ZN(n2077) );
  INV_X1 U2089 ( .A(n2077), .ZN(n2078) );
  INV_X1 U2090 ( .A(n2077), .ZN(n2079) );
  INV_X1 U2091 ( .A(n830), .ZN(n20801) );
  INV_X1 U2092 ( .A(n830), .ZN(n2081) );
  INV_X1 U2093 ( .A(n3377), .ZN(n2082) );
  INV_X1 U2094 ( .A(n2082), .ZN(n2083) );
  INV_X1 U2095 ( .A(n2082), .ZN(n2084) );
  INV_X1 U2096 ( .A(n3375), .ZN(n2085) );
  INV_X1 U2097 ( .A(n2085), .ZN(n2086) );
  INV_X1 U2098 ( .A(n2085), .ZN(n2087) );
  INV_X1 U2099 ( .A(n3427), .ZN(n2088) );
  INV_X1 U2100 ( .A(n2088), .ZN(n2089) );
  INV_X1 U2101 ( .A(n2088), .ZN(n20901) );
  CLKBUF_X1 U2102 ( .A(n3701), .Z(n2091) );
  INV_X1 U2103 ( .A(n3384), .ZN(n2092) );
  INV_X1 U2104 ( .A(n2092), .ZN(n2093) );
  INV_X1 U2105 ( .A(n2092), .ZN(n2094) );
  CLKBUF_X1 U2106 ( .A(n37001), .Z(n2095) );
  INV_X1 U2107 ( .A(n1112), .ZN(n2096) );
  INV_X1 U2108 ( .A(n2096), .ZN(n2097) );
  INV_X1 U2109 ( .A(n2096), .ZN(n2098) );
  INV_X1 U2110 ( .A(n3224), .ZN(n2099) );
  INV_X1 U2111 ( .A(n2099), .ZN(n21001) );
  INV_X1 U2112 ( .A(n2099), .ZN(n2101) );
  INV_X1 U2113 ( .A(n831), .ZN(n2102) );
  INV_X1 U2114 ( .A(n831), .ZN(n2103) );
  INV_X1 U2115 ( .A(n832), .ZN(n2104) );
  INV_X1 U2116 ( .A(n832), .ZN(n2105) );
  INV_X1 U2117 ( .A(n3394), .ZN(n2106) );
  INV_X1 U2118 ( .A(n2106), .ZN(n2107) );
  INV_X1 U2119 ( .A(n2106), .ZN(n2108) );
  INV_X1 U2120 ( .A(n833), .ZN(n2109) );
  INV_X1 U2121 ( .A(n833), .ZN(n21101) );
  INV_X1 U2122 ( .A(n3398), .ZN(n2111) );
  INV_X1 U2123 ( .A(n2111), .ZN(n2112) );
  INV_X1 U2124 ( .A(n2111), .ZN(n2113) );
  INV_X1 U2125 ( .A(n1114), .ZN(n2114) );
  INV_X1 U2126 ( .A(n2114), .ZN(n2115) );
  INV_X1 U2127 ( .A(n2114), .ZN(n2116) );
  INV_X1 U2128 ( .A(n3403), .ZN(n2117) );
  INV_X1 U2129 ( .A(n2117), .ZN(n2118) );
  INV_X1 U2130 ( .A(n2117), .ZN(n2119) );
  INV_X1 U2131 ( .A(n1791), .ZN(n21201) );
  INV_X1 U2132 ( .A(n21201), .ZN(n2121) );
  INV_X1 U2133 ( .A(n21201), .ZN(n2122) );
  INV_X1 U2134 ( .A(n3412), .ZN(n2123) );
  INV_X1 U2135 ( .A(n2123), .ZN(n2124) );
  INV_X1 U2136 ( .A(n2123), .ZN(n2125) );
  INV_X1 U2137 ( .A(n15590), .ZN(n2126) );
  INV_X1 U2138 ( .A(n2126), .ZN(n2127) );
  INV_X1 U2139 ( .A(n2126), .ZN(n2128) );
  INV_X1 U2140 ( .A(n3413), .ZN(n2129) );
  INV_X1 U2141 ( .A(n2129), .ZN(n21301) );
  INV_X1 U2142 ( .A(n2129), .ZN(n2131) );
  INV_X1 U2143 ( .A(n1118), .ZN(n2132) );
  INV_X1 U2144 ( .A(n2132), .ZN(n2133) );
  INV_X1 U2145 ( .A(n2132), .ZN(n2134) );
  INV_X1 U2146 ( .A(n3416), .ZN(n2135) );
  INV_X1 U2147 ( .A(n2135), .ZN(n2136) );
  INV_X1 U2148 ( .A(n2135), .ZN(n2137) );
  INV_X1 U2149 ( .A(n1119), .ZN(n2138) );
  INV_X1 U2150 ( .A(n2138), .ZN(n2139) );
  INV_X1 U2151 ( .A(n2138), .ZN(n21401) );
  INV_X1 U2152 ( .A(n3418), .ZN(n2141) );
  INV_X1 U2153 ( .A(n2141), .ZN(n2142) );
  INV_X1 U2154 ( .A(n2141), .ZN(n2143) );
  INV_X1 U2155 ( .A(n34201), .ZN(n2144) );
  INV_X1 U2156 ( .A(n2144), .ZN(n2145) );
  INV_X1 U2157 ( .A(n2144), .ZN(n2146) );
  INV_X1 U2158 ( .A(n3427), .ZN(n2147) );
  INV_X1 U2159 ( .A(n2147), .ZN(n2148) );
  INV_X1 U2160 ( .A(n2147), .ZN(n2149) );
  INV_X1 U2161 ( .A(n834), .ZN(n21501) );
  INV_X1 U2162 ( .A(n834), .ZN(n2151) );
  INV_X1 U2163 ( .A(n835), .ZN(n2152) );
  INV_X1 U2164 ( .A(n835), .ZN(n2153) );
  INV_X1 U2165 ( .A(n3429), .ZN(n2154) );
  INV_X1 U2166 ( .A(n2154), .ZN(n2155) );
  INV_X1 U2167 ( .A(n2154), .ZN(n2156) );
  INV_X1 U2168 ( .A(n34301), .ZN(n2157) );
  INV_X1 U2169 ( .A(n2157), .ZN(n2158) );
  INV_X1 U2170 ( .A(n2157), .ZN(n2159) );
  INV_X1 U2171 ( .A(n961), .ZN(n21601) );
  INV_X1 U2172 ( .A(n21601), .ZN(n2161) );
  INV_X1 U2173 ( .A(n21601), .ZN(n2162) );
  INV_X1 U2174 ( .A(n4061), .ZN(n2163) );
  INV_X1 U2175 ( .A(n2689), .ZN(n2164) );
  INV_X1 U2176 ( .A(n961), .ZN(n2165) );
  INV_X1 U2177 ( .A(n2165), .ZN(n2166) );
  INV_X1 U2178 ( .A(n2165), .ZN(n2167) );
  INV_X1 U2179 ( .A(n836), .ZN(n2168) );
  INV_X1 U2180 ( .A(n836), .ZN(n2169) );
  INV_X1 U2181 ( .A(n3437), .ZN(n21701) );
  INV_X1 U2182 ( .A(n21701), .ZN(n2171) );
  INV_X1 U2183 ( .A(n21701), .ZN(n2172) );
  INV_X1 U2184 ( .A(n3437), .ZN(n2173) );
  INV_X1 U2185 ( .A(n2173), .ZN(n2174) );
  INV_X1 U2186 ( .A(n2173), .ZN(n2175) );
  INV_X1 U2187 ( .A(n3307), .ZN(n2176) );
  INV_X1 U2188 ( .A(n2176), .ZN(n2177) );
  INV_X1 U2189 ( .A(n2176), .ZN(n2178) );
  INV_X1 U2190 ( .A(n34401), .ZN(n2179) );
  INV_X1 U2191 ( .A(n2179), .ZN(n21801) );
  INV_X1 U2192 ( .A(n2179), .ZN(n2181) );
  INV_X1 U2193 ( .A(n34401), .ZN(n2182) );
  INV_X1 U2194 ( .A(n2182), .ZN(n2183) );
  INV_X1 U2195 ( .A(n2182), .ZN(n2184) );
  INV_X1 U2196 ( .A(n3441), .ZN(n2185) );
  INV_X1 U2197 ( .A(n2185), .ZN(n2186) );
  INV_X1 U2198 ( .A(n2185), .ZN(n2187) );
  INV_X1 U2199 ( .A(n3441), .ZN(n2188) );
  INV_X1 U2200 ( .A(n2188), .ZN(n2189) );
  INV_X1 U2201 ( .A(n2188), .ZN(n21901) );
  INV_X1 U2202 ( .A(n3443), .ZN(n2191) );
  INV_X1 U2203 ( .A(n2191), .ZN(n2192) );
  INV_X1 U2204 ( .A(n2191), .ZN(n2193) );
  INV_X1 U2205 ( .A(n3442), .ZN(n2194) );
  INV_X1 U2206 ( .A(n2194), .ZN(n2195) );
  INV_X1 U2207 ( .A(n2194), .ZN(n2196) );
  INV_X1 U2208 ( .A(n3442), .ZN(n2197) );
  INV_X1 U2209 ( .A(n2197), .ZN(n2198) );
  INV_X1 U2210 ( .A(n2197), .ZN(n2199) );
  INV_X1 U2211 ( .A(n3443), .ZN(n22001) );
  INV_X1 U2212 ( .A(n22001), .ZN(n2201) );
  INV_X1 U2213 ( .A(n22001), .ZN(n2202) );
  INV_X1 U2214 ( .A(n29401), .ZN(n2203) );
  INV_X1 U2215 ( .A(n2203), .ZN(n2204) );
  INV_X1 U2216 ( .A(n2203), .ZN(n2205) );
  INV_X1 U2217 ( .A(n3445), .ZN(n2206) );
  INV_X1 U2218 ( .A(n2206), .ZN(n2207) );
  INV_X1 U2219 ( .A(n2206), .ZN(n2208) );
  INV_X1 U2220 ( .A(n837), .ZN(n2209) );
  INV_X1 U2221 ( .A(n837), .ZN(n22101) );
  INV_X1 U2222 ( .A(n838), .ZN(n2211) );
  INV_X1 U2223 ( .A(n838), .ZN(n2212) );
  INV_X1 U2224 ( .A(n3415), .ZN(n2213) );
  INV_X1 U2225 ( .A(n2213), .ZN(n2214) );
  INV_X1 U2226 ( .A(n2213), .ZN(n2215) );
  INV_X1 U2227 ( .A(n839), .ZN(n2216) );
  INV_X1 U2228 ( .A(n839), .ZN(n2217) );
  INV_X1 U2229 ( .A(n843), .ZN(n2218) );
  INV_X1 U2230 ( .A(n2218), .ZN(n2219) );
  INV_X1 U2231 ( .A(n2218), .ZN(n22201) );
  INV_X1 U2232 ( .A(n843), .ZN(n2221) );
  INV_X1 U2233 ( .A(n2221), .ZN(n2222) );
  INV_X1 U2234 ( .A(n2221), .ZN(n2223) );
  INV_X1 U2235 ( .A(n842), .ZN(n2224) );
  INV_X1 U2236 ( .A(n842), .ZN(n2225) );
  INV_X1 U2237 ( .A(n4678), .ZN(n2226) );
  INV_X1 U2238 ( .A(n844), .ZN(n2227) );
  INV_X1 U2239 ( .A(n844), .ZN(n2228) );
  INV_X1 U2240 ( .A(n845), .ZN(n2229) );
  INV_X1 U2241 ( .A(n845), .ZN(n22301) );
  INV_X1 U2242 ( .A(n847), .ZN(n2231) );
  INV_X1 U2243 ( .A(n2231), .ZN(n2232) );
  INV_X1 U2244 ( .A(n2231), .ZN(n2233) );
  INV_X1 U2245 ( .A(n846), .ZN(n2234) );
  INV_X1 U2246 ( .A(n846), .ZN(n2235) );
  INV_X1 U2247 ( .A(n4138), .ZN(n2236) );
  INV_X1 U2248 ( .A(n2236), .ZN(n2237) );
  INV_X1 U2249 ( .A(n2236), .ZN(n2238) );
  INV_X1 U2250 ( .A(n849), .ZN(n2239) );
  INV_X1 U2251 ( .A(n2239), .ZN(n22401) );
  INV_X1 U2252 ( .A(n2239), .ZN(n2241) );
  INV_X1 U2253 ( .A(n847), .ZN(n2242) );
  INV_X1 U2254 ( .A(n848), .ZN(n2243) );
  INV_X1 U2255 ( .A(n848), .ZN(n2244) );
  INV_X1 U2256 ( .A(n849), .ZN(n2245) );
  INV_X1 U2257 ( .A(n2245), .ZN(n2246) );
  INV_X1 U2258 ( .A(n2245), .ZN(n2247) );
  INV_X1 U2259 ( .A(n38301), .ZN(n2248) );
  INV_X1 U2260 ( .A(n2248), .ZN(n2249) );
  INV_X1 U2261 ( .A(n38301), .ZN(n22501) );
  INV_X1 U2262 ( .A(n2249), .ZN(n2251) );
  INV_X1 U2263 ( .A(n33201), .ZN(n2252) );
  INV_X1 U2264 ( .A(n2252), .ZN(n2253) );
  INV_X1 U2265 ( .A(n2252), .ZN(n2254) );
  INV_X1 U2266 ( .A(n3321), .ZN(n2255) );
  INV_X1 U2267 ( .A(n2255), .ZN(n2256) );
  INV_X1 U2268 ( .A(n2255), .ZN(n2257) );
  INV_X1 U2269 ( .A(n3319), .ZN(n2258) );
  INV_X1 U2270 ( .A(n2258), .ZN(n2259) );
  INV_X1 U2271 ( .A(n2258), .ZN(n22601) );
  INV_X1 U2272 ( .A(n852), .ZN(n2261) );
  INV_X1 U2273 ( .A(n2261), .ZN(n2262) );
  INV_X1 U2274 ( .A(n2261), .ZN(n2263) );
  INV_X1 U2275 ( .A(n34201), .ZN(n2264) );
  INV_X1 U2276 ( .A(n2264), .ZN(n2265) );
  INV_X1 U2277 ( .A(n2264), .ZN(n2266) );
  INV_X1 U2278 ( .A(n851), .ZN(n2267) );
  INV_X1 U2279 ( .A(n851), .ZN(n2268) );
  INV_X1 U2280 ( .A(n852), .ZN(n2269) );
  INV_X1 U2281 ( .A(n2269), .ZN(n22701) );
  INV_X1 U2282 ( .A(n2269), .ZN(n2271) );
  INV_X1 U2283 ( .A(n4674), .ZN(n2272) );
  INV_X1 U2284 ( .A(n2272), .ZN(n2273) );
  INV_X1 U2285 ( .A(n4674), .ZN(n2274) );
  INV_X1 U2286 ( .A(n2273), .ZN(n2275) );
  INV_X1 U2287 ( .A(n853), .ZN(n2276) );
  INV_X1 U2288 ( .A(n853), .ZN(n2277) );
  INV_X1 U2289 ( .A(n855), .ZN(n2278) );
  INV_X1 U2290 ( .A(n2278), .ZN(n2279) );
  INV_X1 U2291 ( .A(n2278), .ZN(n22801) );
  INV_X1 U2292 ( .A(n854), .ZN(n2281) );
  INV_X1 U2293 ( .A(n854), .ZN(n2282) );
  INV_X1 U2294 ( .A(n855), .ZN(n2283) );
  INV_X1 U2295 ( .A(n2283), .ZN(n2284) );
  INV_X1 U2296 ( .A(n2283), .ZN(n2285) );
  INV_X1 U2297 ( .A(n857), .ZN(n2286) );
  INV_X1 U2298 ( .A(n2286), .ZN(n2287) );
  INV_X1 U2299 ( .A(n2286), .ZN(n2288) );
  INV_X1 U2300 ( .A(n856), .ZN(n2289) );
  INV_X1 U2301 ( .A(n856), .ZN(n22901) );
  INV_X1 U2302 ( .A(n857), .ZN(n2291) );
  INV_X1 U2303 ( .A(n2291), .ZN(n2292) );
  INV_X1 U2304 ( .A(n2291), .ZN(n2293) );
  INV_X1 U2305 ( .A(n4536), .ZN(n2294) );
  INV_X1 U2306 ( .A(n2294), .ZN(n2295) );
  INV_X1 U2307 ( .A(n4536), .ZN(n2296) );
  INV_X1 U2308 ( .A(n2295), .ZN(n2297) );
  INV_X1 U2309 ( .A(n4538), .ZN(n2298) );
  INV_X1 U2310 ( .A(n2298), .ZN(n2299) );
  INV_X1 U2311 ( .A(n2298), .ZN(n23001) );
  INV_X1 U2312 ( .A(n2313), .ZN(n2301) );
  INV_X1 U2313 ( .A(n2301), .ZN(n2302) );
  INV_X1 U2314 ( .A(n2301), .ZN(n2303) );
  INV_X1 U2315 ( .A(n2313), .ZN(n2304) );
  INV_X1 U2316 ( .A(n2304), .ZN(n2305) );
  INV_X1 U2317 ( .A(n2304), .ZN(n2306) );
  INV_X1 U2318 ( .A(n4538), .ZN(n2307) );
  INV_X1 U2319 ( .A(n2307), .ZN(n2308) );
  INV_X1 U2320 ( .A(n2307), .ZN(n2309) );
  INV_X1 U2321 ( .A(n859), .ZN(n23101) );
  INV_X1 U2322 ( .A(n23101), .ZN(n2311) );
  INV_X1 U2323 ( .A(n23101), .ZN(n2312) );
  INV_X1 U2324 ( .A(n4604), .ZN(n2313) );
  INV_X1 U2325 ( .A(n858), .ZN(n2314) );
  INV_X1 U2326 ( .A(n858), .ZN(n2315) );
  INV_X1 U2327 ( .A(n859), .ZN(n2316) );
  INV_X1 U2328 ( .A(n2316), .ZN(n2317) );
  INV_X1 U2329 ( .A(n2316), .ZN(n2318) );
  INV_X1 U2330 ( .A(n4401), .ZN(n2319) );
  INV_X1 U2331 ( .A(n2319), .ZN(n23201) );
  INV_X1 U2332 ( .A(n4401), .ZN(n2321) );
  INV_X1 U2333 ( .A(n23201), .ZN(n2322) );
  INV_X1 U2334 ( .A(n860), .ZN(n2323) );
  INV_X1 U2335 ( .A(n860), .ZN(n2324) );
  INV_X1 U2336 ( .A(n862), .ZN(n2325) );
  INV_X1 U2337 ( .A(n2325), .ZN(n2326) );
  INV_X1 U2338 ( .A(n2325), .ZN(n2327) );
  INV_X1 U2339 ( .A(n861), .ZN(n2328) );
  INV_X1 U2340 ( .A(n861), .ZN(n2329) );
  INV_X1 U2341 ( .A(n862), .ZN(n23301) );
  INV_X1 U2342 ( .A(n23301), .ZN(n2331) );
  INV_X1 U2343 ( .A(n23301), .ZN(n2332) );
  INV_X1 U2344 ( .A(n864), .ZN(n2333) );
  INV_X1 U2345 ( .A(n2333), .ZN(n2334) );
  INV_X1 U2346 ( .A(n2333), .ZN(n2335) );
  INV_X1 U2347 ( .A(n863), .ZN(n2336) );
  INV_X1 U2348 ( .A(n863), .ZN(n2337) );
  INV_X1 U2349 ( .A(n864), .ZN(n2338) );
  INV_X1 U2350 ( .A(n2338), .ZN(n2339) );
  INV_X1 U2351 ( .A(n2338), .ZN(n23401) );
  INV_X1 U2352 ( .A(n4263), .ZN(n2341) );
  INV_X1 U2353 ( .A(n2341), .ZN(n2342) );
  INV_X1 U2354 ( .A(n4263), .ZN(n2343) );
  INV_X1 U2355 ( .A(n2342), .ZN(n2344) );
  INV_X1 U2356 ( .A(n4264), .ZN(n2345) );
  INV_X1 U2357 ( .A(n2345), .ZN(n2346) );
  INV_X1 U2358 ( .A(n2345), .ZN(n2347) );
  INV_X1 U2359 ( .A(n23601), .ZN(n2348) );
  INV_X1 U2360 ( .A(n2348), .ZN(n2349) );
  INV_X1 U2361 ( .A(n2348), .ZN(n23501) );
  INV_X1 U2362 ( .A(n23601), .ZN(n2351) );
  INV_X1 U2363 ( .A(n2351), .ZN(n2352) );
  INV_X1 U2364 ( .A(n2351), .ZN(n2353) );
  INV_X1 U2365 ( .A(n4264), .ZN(n2354) );
  INV_X1 U2366 ( .A(n2354), .ZN(n2355) );
  INV_X1 U2367 ( .A(n2354), .ZN(n2356) );
  INV_X1 U2368 ( .A(n866), .ZN(n2357) );
  INV_X1 U2369 ( .A(n2357), .ZN(n2358) );
  INV_X1 U2370 ( .A(n2357), .ZN(n2359) );
  INV_X1 U2371 ( .A(n4333), .ZN(n23601) );
  INV_X1 U2372 ( .A(n865), .ZN(n2361) );
  INV_X1 U2373 ( .A(n865), .ZN(n2362) );
  INV_X1 U2374 ( .A(n866), .ZN(n2363) );
  INV_X1 U2375 ( .A(n2363), .ZN(n2364) );
  INV_X1 U2376 ( .A(n2363), .ZN(n2365) );
  INV_X1 U2377 ( .A(n3964), .ZN(n2366) );
  INV_X1 U2378 ( .A(n2366), .ZN(n2367) );
  INV_X1 U2379 ( .A(n3964), .ZN(n2368) );
  INV_X1 U2380 ( .A(n2367), .ZN(n2369) );
  INV_X1 U2381 ( .A(n867), .ZN(n23701) );
  INV_X1 U2382 ( .A(n867), .ZN(n2371) );
  INV_X1 U2383 ( .A(n869), .ZN(n2372) );
  INV_X1 U2384 ( .A(n2372), .ZN(n2373) );
  INV_X1 U2385 ( .A(n2372), .ZN(n2374) );
  INV_X1 U2386 ( .A(n868), .ZN(n2375) );
  INV_X1 U2387 ( .A(n868), .ZN(n2376) );
  INV_X1 U2388 ( .A(n869), .ZN(n2377) );
  INV_X1 U2389 ( .A(n2377), .ZN(n2378) );
  INV_X1 U2390 ( .A(n2377), .ZN(n2379) );
  INV_X1 U2391 ( .A(n871), .ZN(n23801) );
  INV_X1 U2392 ( .A(n23801), .ZN(n2381) );
  INV_X1 U2393 ( .A(n23801), .ZN(n2382) );
  INV_X1 U2394 ( .A(n870), .ZN(n2383) );
  INV_X1 U2395 ( .A(n870), .ZN(n2384) );
  INV_X1 U2396 ( .A(n871), .ZN(n2385) );
  INV_X1 U2397 ( .A(n2385), .ZN(n2386) );
  INV_X1 U2398 ( .A(n2385), .ZN(n2387) );
  INV_X1 U2399 ( .A(n3866), .ZN(n2388) );
  INV_X1 U2400 ( .A(n2388), .ZN(n2389) );
  INV_X1 U2401 ( .A(n3866), .ZN(n23901) );
  INV_X1 U2402 ( .A(n2389), .ZN(n2391) );
  INV_X1 U2403 ( .A(n872), .ZN(n2392) );
  INV_X1 U2404 ( .A(n872), .ZN(n2393) );
  INV_X1 U2405 ( .A(n875), .ZN(n2394) );
  INV_X1 U2406 ( .A(n2394), .ZN(n2395) );
  INV_X1 U2407 ( .A(n2394), .ZN(n2396) );
  INV_X1 U2408 ( .A(n873), .ZN(n2397) );
  INV_X1 U2409 ( .A(n873), .ZN(n2398) );
  INV_X1 U2410 ( .A(n875), .ZN(n2399) );
  INV_X1 U2411 ( .A(n2399), .ZN(n24001) );
  INV_X1 U2412 ( .A(n2399), .ZN(n2401) );
  INV_X1 U2413 ( .A(n874), .ZN(n2402) );
  INV_X1 U2414 ( .A(n874), .ZN(n2403) );
  INV_X1 U2415 ( .A(n876), .ZN(n2404) );
  INV_X1 U2416 ( .A(n876), .ZN(n2405) );
  INV_X1 U2417 ( .A(n877), .ZN(n2406) );
  INV_X1 U2418 ( .A(n877), .ZN(n2407) );
  INV_X1 U2419 ( .A(n3697), .ZN(n2408) );
  INV_X1 U2420 ( .A(n3697), .ZN(n2409) );
  INV_X1 U2421 ( .A(n878), .ZN(n24101) );
  INV_X1 U2422 ( .A(n878), .ZN(n2411) );
  INV_X1 U2423 ( .A(n3723), .ZN(n2412) );
  INV_X1 U2424 ( .A(n2412), .ZN(n2413) );
  INV_X1 U2425 ( .A(n2412), .ZN(n2414) );
  INV_X1 U2426 ( .A(n2426), .ZN(n2415) );
  INV_X1 U2427 ( .A(n2415), .ZN(n2416) );
  INV_X1 U2428 ( .A(n2415), .ZN(n2417) );
  INV_X1 U2429 ( .A(n2426), .ZN(n2418) );
  INV_X1 U2430 ( .A(n2418), .ZN(n2419) );
  INV_X1 U2431 ( .A(n2418), .ZN(n24201) );
  INV_X1 U2432 ( .A(n3723), .ZN(n2421) );
  INV_X1 U2433 ( .A(n2421), .ZN(n2422) );
  INV_X1 U2434 ( .A(n2421), .ZN(n2423) );
  INV_X1 U2435 ( .A(n879), .ZN(n2424) );
  INV_X1 U2436 ( .A(n879), .ZN(n2425) );
  INV_X1 U2437 ( .A(n3757), .ZN(n2426) );
  INV_X1 U2438 ( .A(n880), .ZN(n2427) );
  INV_X1 U2439 ( .A(n880), .ZN(n2428) );
  INV_X1 U2440 ( .A(n881), .ZN(n2429) );
  INV_X1 U2441 ( .A(n881), .ZN(n24301) );
  INV_X1 U2442 ( .A(n3313), .ZN(n2431) );
  INV_X1 U2443 ( .A(n2431), .ZN(n2432) );
  INV_X1 U2444 ( .A(n2431), .ZN(n2433) );
  INV_X1 U2445 ( .A(n882), .ZN(n2434) );
  INV_X1 U2446 ( .A(n882), .ZN(n2435) );
  INV_X1 U2447 ( .A(n884), .ZN(n2436) );
  INV_X1 U2448 ( .A(n2436), .ZN(n2437) );
  INV_X1 U2449 ( .A(n2436), .ZN(n2438) );
  INV_X1 U2450 ( .A(n885), .ZN(n2439) );
  INV_X1 U2451 ( .A(n2439), .ZN(n24401) );
  INV_X1 U2452 ( .A(n2439), .ZN(n2441) );
  INV_X1 U2453 ( .A(n3698), .ZN(n2442) );
  INV_X1 U2454 ( .A(n2442), .ZN(n2443) );
  INV_X1 U2455 ( .A(n2442), .ZN(n2444) );
  INV_X1 U2456 ( .A(n885), .ZN(n2445) );
  INV_X1 U2457 ( .A(n2445), .ZN(n2446) );
  INV_X1 U2458 ( .A(n2445), .ZN(n2447) );
  INV_X1 U2459 ( .A(n883), .ZN(n2448) );
  INV_X1 U2460 ( .A(n883), .ZN(n2449) );
  INV_X1 U2461 ( .A(n886), .ZN(n24501) );
  INV_X1 U2462 ( .A(n886), .ZN(n2451) );
  INV_X1 U2463 ( .A(n887), .ZN(n2452) );
  INV_X1 U2464 ( .A(n887), .ZN(n2453) );
  INV_X1 U2465 ( .A(n888), .ZN(n2454) );
  INV_X1 U2466 ( .A(n888), .ZN(n2455) );
  INV_X1 U2467 ( .A(n889), .ZN(n2456) );
  INV_X1 U2468 ( .A(n889), .ZN(n2457) );
  INV_X1 U2469 ( .A(n892), .ZN(n2458) );
  INV_X1 U2470 ( .A(n2458), .ZN(n2459) );
  INV_X1 U2471 ( .A(n2458), .ZN(n24601) );
  INV_X1 U2472 ( .A(n891), .ZN(n2461) );
  INV_X1 U2473 ( .A(n2461), .ZN(n2462) );
  INV_X1 U2474 ( .A(n2461), .ZN(n2463) );
  INV_X1 U2475 ( .A(n892), .ZN(n2464) );
  INV_X1 U2476 ( .A(n2464), .ZN(n2465) );
  INV_X1 U2477 ( .A(n2464), .ZN(n2466) );
  INV_X1 U2478 ( .A(n1129), .ZN(n2467) );
  INV_X1 U2479 ( .A(n2467), .ZN(n2468) );
  INV_X1 U2480 ( .A(n2467), .ZN(n2469) );
  INV_X1 U2481 ( .A(n890), .ZN(n24701) );
  INV_X1 U2482 ( .A(n890), .ZN(n2471) );
  INV_X1 U2483 ( .A(n893), .ZN(n2472) );
  INV_X1 U2484 ( .A(n893), .ZN(n2473) );
  INV_X1 U2485 ( .A(n894), .ZN(n2474) );
  INV_X1 U2486 ( .A(n894), .ZN(n2475) );
  INV_X1 U2487 ( .A(n895), .ZN(n2476) );
  INV_X1 U2488 ( .A(n895), .ZN(n2477) );
  INV_X1 U2489 ( .A(n896), .ZN(n2478) );
  INV_X1 U2490 ( .A(n896), .ZN(n2479) );
  INV_X1 U2491 ( .A(n897), .ZN(n24801) );
  INV_X1 U2492 ( .A(n897), .ZN(n2481) );
  INV_X1 U2493 ( .A(n898), .ZN(n2482) );
  INV_X1 U2494 ( .A(n898), .ZN(n2483) );
  INV_X1 U2495 ( .A(n899), .ZN(n2484) );
  INV_X1 U2496 ( .A(n899), .ZN(n2485) );
  INV_X1 U2497 ( .A(n900), .ZN(n2486) );
  INV_X1 U2498 ( .A(n900), .ZN(n2487) );
  INV_X1 U2499 ( .A(n901), .ZN(n2488) );
  INV_X1 U2500 ( .A(n901), .ZN(n2489) );
  INV_X1 U2501 ( .A(n902), .ZN(n24901) );
  INV_X1 U2502 ( .A(n902), .ZN(n2491) );
  INV_X1 U2503 ( .A(n903), .ZN(n2492) );
  INV_X1 U2504 ( .A(n903), .ZN(n2493) );
  INV_X1 U2505 ( .A(n904), .ZN(n2494) );
  INV_X1 U2506 ( .A(n904), .ZN(n2495) );
  INV_X1 U2507 ( .A(n3312), .ZN(n2496) );
  INV_X1 U2508 ( .A(n2496), .ZN(n2497) );
  INV_X1 U2509 ( .A(n2496), .ZN(n2498) );
  INV_X1 U2510 ( .A(n905), .ZN(n2499) );
  INV_X1 U2511 ( .A(n905), .ZN(n25001) );
  INV_X1 U2512 ( .A(n906), .ZN(n2501) );
  INV_X1 U2513 ( .A(n906), .ZN(n2502) );
  INV_X1 U2514 ( .A(n907), .ZN(n2503) );
  INV_X1 U2515 ( .A(n907), .ZN(n2504) );
  INV_X1 U2516 ( .A(n909), .ZN(n2505) );
  INV_X1 U2517 ( .A(n2505), .ZN(n2506) );
  INV_X1 U2518 ( .A(n2505), .ZN(n2507) );
  INV_X1 U2519 ( .A(n908), .ZN(n2508) );
  INV_X1 U2520 ( .A(n908), .ZN(n2509) );
  INV_X1 U2521 ( .A(n3309), .ZN(n25101) );
  INV_X1 U2522 ( .A(n25101), .ZN(n2511) );
  INV_X1 U2523 ( .A(n25101), .ZN(n2512) );
  INV_X1 U2524 ( .A(n3311), .ZN(n2513) );
  INV_X1 U2525 ( .A(n2513), .ZN(n2514) );
  INV_X1 U2526 ( .A(n2513), .ZN(n2515) );
  INV_X1 U2527 ( .A(n3307), .ZN(n2516) );
  INV_X1 U2528 ( .A(n2516), .ZN(n2517) );
  INV_X1 U2529 ( .A(n2516), .ZN(n2518) );
  INV_X1 U2530 ( .A(n3308), .ZN(n2519) );
  INV_X1 U2531 ( .A(n2519), .ZN(n25201) );
  INV_X1 U2532 ( .A(n2519), .ZN(n2521) );
  INV_X1 U2533 ( .A(n3305), .ZN(n2522) );
  INV_X1 U2534 ( .A(n2522), .ZN(n2523) );
  INV_X1 U2535 ( .A(n2522), .ZN(n2524) );
  INV_X1 U2536 ( .A(n42001), .ZN(n2525) );
  INV_X1 U2537 ( .A(n42001), .ZN(n2526) );
  INV_X1 U2538 ( .A(n3758), .ZN(n2527) );
  INV_X1 U2539 ( .A(n3758), .ZN(n2528) );
  INV_X1 U2540 ( .A(n3303), .ZN(n2529) );
  INV_X1 U2541 ( .A(n2529), .ZN(n25301) );
  INV_X1 U2542 ( .A(n2529), .ZN(n2531) );
  INV_X1 U2543 ( .A(n910), .ZN(n2532) );
  INV_X1 U2544 ( .A(n910), .ZN(n2533) );
  INV_X1 U2545 ( .A(n3299), .ZN(n2534) );
  INV_X1 U2546 ( .A(n2534), .ZN(n2535) );
  INV_X1 U2547 ( .A(n2534), .ZN(n2536) );
  INV_X1 U2548 ( .A(n3715), .ZN(n2537) );
  INV_X1 U2549 ( .A(n2537), .ZN(n2538) );
  INV_X1 U2550 ( .A(n2537), .ZN(n2539) );
  INV_X1 U2551 ( .A(n3705), .ZN(n25401) );
  INV_X1 U2552 ( .A(n3705), .ZN(n2541) );
  INV_X1 U2553 ( .A(n913), .ZN(n2542) );
  INV_X1 U2554 ( .A(n913), .ZN(n2543) );
  INV_X1 U2555 ( .A(n1063), .ZN(n2544) );
  INV_X1 U2556 ( .A(n2544), .ZN(n2545) );
  INV_X1 U2557 ( .A(n3702), .ZN(n2546) );
  INV_X1 U2558 ( .A(n3702), .ZN(n2547) );
  INV_X1 U2559 ( .A(n914), .ZN(n2548) );
  INV_X1 U2560 ( .A(n914), .ZN(n2549) );
  INV_X1 U2561 ( .A(n916), .ZN(n25501) );
  INV_X1 U2562 ( .A(n916), .ZN(n2551) );
  INV_X1 U2563 ( .A(n917), .ZN(n2552) );
  INV_X1 U2564 ( .A(n917), .ZN(n2553) );
  INV_X1 U2565 ( .A(n3265), .ZN(n2554) );
  INV_X1 U2566 ( .A(n2554), .ZN(n2555) );
  INV_X1 U2567 ( .A(n2554), .ZN(n2556) );
  INV_X1 U2568 ( .A(n918), .ZN(n2557) );
  INV_X1 U2569 ( .A(n918), .ZN(n2558) );
  INV_X1 U2570 ( .A(n919), .ZN(n2559) );
  INV_X1 U2571 ( .A(n919), .ZN(n25601) );
  INV_X1 U2572 ( .A(n921), .ZN(n2561) );
  INV_X1 U2573 ( .A(n921), .ZN(n2562) );
  INV_X1 U2574 ( .A(n922), .ZN(n2563) );
  INV_X1 U2575 ( .A(n922), .ZN(n2564) );
  INV_X1 U2576 ( .A(n923), .ZN(n2565) );
  INV_X1 U2577 ( .A(n923), .ZN(n2566) );
  INV_X1 U2578 ( .A(n1618), .ZN(n2567) );
  INV_X1 U2579 ( .A(n2567), .ZN(n2568) );
  INV_X1 U2580 ( .A(n2567), .ZN(n2569) );
  INV_X1 U2581 ( .A(n1618), .ZN(n25701) );
  INV_X1 U2582 ( .A(n25701), .ZN(n2571) );
  INV_X1 U2583 ( .A(n25701), .ZN(n2572) );
  INV_X1 U2584 ( .A(n9240), .ZN(n2573) );
  INV_X1 U2585 ( .A(n9240), .ZN(n2574) );
  INV_X1 U2586 ( .A(n9250), .ZN(n2575) );
  INV_X1 U2587 ( .A(n1536), .ZN(n2576) );
  INV_X1 U2588 ( .A(n9260), .ZN(n2577) );
  INV_X1 U2589 ( .A(n9270), .ZN(n2578) );
  INV_X1 U2590 ( .A(n9270), .ZN(n2579) );
  INV_X1 U2591 ( .A(n3759), .ZN(n25801) );
  INV_X1 U2592 ( .A(n3759), .ZN(n2581) );
  INV_X1 U2593 ( .A(n9280), .ZN(n2582) );
  INV_X1 U2594 ( .A(n9280), .ZN(n2583) );
  INV_X1 U2595 ( .A(n9290), .ZN(n2584) );
  INV_X1 U2596 ( .A(n9290), .ZN(n2585) );
  INV_X1 U2597 ( .A(n3226), .ZN(n2586) );
  INV_X1 U2598 ( .A(n2586), .ZN(n2587) );
  INV_X1 U2599 ( .A(n2586), .ZN(n2588) );
  INV_X1 U2600 ( .A(n3421), .ZN(n2589) );
  INV_X1 U2601 ( .A(n3424), .ZN(n25901) );
  INV_X1 U2602 ( .A(n9300), .ZN(n2591) );
  INV_X1 U2603 ( .A(n9300), .ZN(n2592) );
  INV_X1 U2604 ( .A(n9310), .ZN(n2593) );
  INV_X1 U2605 ( .A(n9310), .ZN(n2594) );
  INV_X1 U2606 ( .A(n9320), .ZN(n2595) );
  INV_X1 U2607 ( .A(n9320), .ZN(n2596) );
  INV_X1 U2608 ( .A(n9330), .ZN(n2597) );
  INV_X1 U2609 ( .A(n9330), .ZN(n2598) );
  INV_X1 U2610 ( .A(n9340), .ZN(n2599) );
  INV_X1 U2611 ( .A(n9340), .ZN(n26001) );
  INV_X1 U2612 ( .A(n9350), .ZN(n2601) );
  INV_X1 U2613 ( .A(n9350), .ZN(n2602) );
  INV_X1 U2614 ( .A(n9360), .ZN(n2603) );
  INV_X1 U2615 ( .A(n9360), .ZN(n2604) );
  INV_X1 U2616 ( .A(n9370), .ZN(n2605) );
  INV_X1 U2617 ( .A(n9370), .ZN(n2606) );
  INV_X1 U2618 ( .A(n9380), .ZN(n2607) );
  INV_X1 U2619 ( .A(n9380), .ZN(n2608) );
  INV_X1 U2620 ( .A(n9390), .ZN(n2609) );
  INV_X1 U2621 ( .A(n9390), .ZN(n26101) );
  INV_X1 U2622 ( .A(n940), .ZN(n2611) );
  INV_X1 U2623 ( .A(n940), .ZN(n2612) );
  INV_X1 U2624 ( .A(n941), .ZN(n2613) );
  INV_X1 U2625 ( .A(n941), .ZN(n2614) );
  INV_X1 U2626 ( .A(n942), .ZN(n2615) );
  INV_X1 U2627 ( .A(n942), .ZN(n2616) );
  INV_X1 U2628 ( .A(n943), .ZN(n2617) );
  INV_X1 U2629 ( .A(n943), .ZN(n2618) );
  INV_X1 U2630 ( .A(n944), .ZN(n2619) );
  INV_X1 U2631 ( .A(n944), .ZN(n26201) );
  INV_X1 U2632 ( .A(n945), .ZN(n2621) );
  INV_X1 U2633 ( .A(n945), .ZN(n2622) );
  INV_X1 U2634 ( .A(n946), .ZN(n2623) );
  INV_X1 U2635 ( .A(n946), .ZN(n2624) );
  INV_X1 U2636 ( .A(n947), .ZN(n2625) );
  INV_X1 U2637 ( .A(n947), .ZN(n2626) );
  INV_X1 U2638 ( .A(n948), .ZN(n2627) );
  INV_X1 U2639 ( .A(n948), .ZN(n2628) );
  INV_X1 U2640 ( .A(n949), .ZN(n2629) );
  INV_X1 U2641 ( .A(n949), .ZN(n26301) );
  INV_X1 U2642 ( .A(n950), .ZN(n2631) );
  INV_X1 U2643 ( .A(n950), .ZN(n2632) );
  INV_X1 U2644 ( .A(n951), .ZN(n2633) );
  INV_X1 U2645 ( .A(n951), .ZN(n2634) );
  INV_X1 U2646 ( .A(n952), .ZN(n2635) );
  INV_X1 U2647 ( .A(n952), .ZN(n2636) );
  INV_X1 U2648 ( .A(n953), .ZN(n2637) );
  INV_X1 U2649 ( .A(n953), .ZN(n2638) );
  INV_X1 U2650 ( .A(n954), .ZN(n2639) );
  INV_X1 U2651 ( .A(n954), .ZN(n26401) );
  INV_X1 U2652 ( .A(n955), .ZN(n2641) );
  INV_X1 U2653 ( .A(n955), .ZN(n2642) );
  INV_X1 U2654 ( .A(n956), .ZN(n2643) );
  INV_X1 U2655 ( .A(n956), .ZN(n2644) );
  INV_X1 U2656 ( .A(n3969), .ZN(n2645) );
  INV_X1 U2657 ( .A(n3969), .ZN(n2646) );
  INV_X1 U2658 ( .A(n3972), .ZN(n2647) );
  INV_X1 U2659 ( .A(n3972), .ZN(n2648) );
  INV_X1 U2660 ( .A(n3974), .ZN(n2649) );
  INV_X1 U2661 ( .A(n3974), .ZN(n26501) );
  INV_X1 U2662 ( .A(n3976), .ZN(n2651) );
  INV_X1 U2663 ( .A(n3976), .ZN(n2652) );
  INV_X1 U2664 ( .A(n3978), .ZN(n2653) );
  INV_X1 U2665 ( .A(n3978), .ZN(n2654) );
  INV_X1 U2666 ( .A(n39801), .ZN(n2655) );
  INV_X1 U2667 ( .A(n39801), .ZN(n2656) );
  INV_X1 U2668 ( .A(n3982), .ZN(n2657) );
  INV_X1 U2669 ( .A(n3982), .ZN(n2658) );
  INV_X1 U2670 ( .A(n3984), .ZN(n2659) );
  INV_X1 U2671 ( .A(n3984), .ZN(n26601) );
  INV_X1 U2672 ( .A(n3986), .ZN(n2661) );
  INV_X1 U2673 ( .A(n3986), .ZN(n2662) );
  INV_X1 U2674 ( .A(n3988), .ZN(n2663) );
  INV_X1 U2675 ( .A(n3988), .ZN(n2664) );
  INV_X1 U2676 ( .A(n39901), .ZN(n2665) );
  INV_X1 U2677 ( .A(n39901), .ZN(n2666) );
  INV_X1 U2678 ( .A(n3992), .ZN(n2667) );
  INV_X1 U2679 ( .A(n3992), .ZN(n2668) );
  INV_X1 U2680 ( .A(n3994), .ZN(n2669) );
  INV_X1 U2681 ( .A(n3994), .ZN(n26701) );
  INV_X1 U2682 ( .A(n3996), .ZN(n2671) );
  INV_X1 U2683 ( .A(n3996), .ZN(n2672) );
  INV_X1 U2684 ( .A(n3998), .ZN(n2673) );
  INV_X1 U2685 ( .A(n3998), .ZN(n2674) );
  INV_X1 U2686 ( .A(n40001), .ZN(n2675) );
  INV_X1 U2687 ( .A(n40001), .ZN(n2676) );
  INV_X1 U2688 ( .A(n957), .ZN(n2677) );
  INV_X1 U2689 ( .A(n957), .ZN(n2678) );
  INV_X1 U2690 ( .A(n958), .ZN(n2679) );
  INV_X1 U2691 ( .A(n958), .ZN(n26801) );
  INV_X1 U2692 ( .A(n959), .ZN(n2681) );
  INV_X1 U2693 ( .A(n959), .ZN(n2682) );
  INV_X1 U2694 ( .A(n4272), .ZN(n2683) );
  INV_X1 U2695 ( .A(n2683), .ZN(n2684) );
  INV_X1 U2696 ( .A(n2683), .ZN(n2685) );
  INV_X1 U2697 ( .A(n960), .ZN(n2686) );
  INV_X1 U2698 ( .A(n960), .ZN(n2687) );
  INV_X1 U2699 ( .A(n4061), .ZN(n2688) );
  INV_X1 U2700 ( .A(n2688), .ZN(n2689) );
  INV_X1 U2701 ( .A(n962), .ZN(n26901) );
  INV_X1 U2702 ( .A(n962), .ZN(n2691) );
  INV_X1 U2703 ( .A(n963), .ZN(n2692) );
  INV_X1 U2704 ( .A(n963), .ZN(n2693) );
  INV_X1 U2705 ( .A(n964), .ZN(n2694) );
  INV_X1 U2706 ( .A(n2535), .ZN(n2695) );
  INV_X1 U2707 ( .A(n965), .ZN(n2696) );
  INV_X1 U2708 ( .A(n966), .ZN(n2697) );
  INV_X1 U2709 ( .A(n10301), .ZN(n2698) );
  INV_X1 U2710 ( .A(n2698), .ZN(n2699) );
  INV_X1 U2711 ( .A(n3468), .ZN(n27001) );
  INV_X1 U2712 ( .A(n27001), .ZN(n2701) );
  INV_X1 U2713 ( .A(n27001), .ZN(n2702) );
  INV_X1 U2714 ( .A(n3444), .ZN(n2703) );
  INV_X1 U2715 ( .A(n2703), .ZN(n2704) );
  INV_X1 U2716 ( .A(n3433), .ZN(n2705) );
  INV_X1 U2717 ( .A(n2705), .ZN(n2706) );
  INV_X1 U2718 ( .A(n3436), .ZN(n2707) );
  INV_X1 U2719 ( .A(n2707), .ZN(n2708) );
  INV_X1 U2720 ( .A(n2714), .ZN(n2709) );
  INV_X1 U2721 ( .A(n2709), .ZN(n27101) );
  INV_X1 U2722 ( .A(n968), .ZN(n2711) );
  INV_X1 U2723 ( .A(n2716), .ZN(n2712) );
  INV_X1 U2724 ( .A(n3415), .ZN(n2713) );
  INV_X1 U2725 ( .A(n2713), .ZN(n2714) );
  INV_X1 U2726 ( .A(n2713), .ZN(n2715) );
  INV_X1 U2727 ( .A(n969), .ZN(n2716) );
  INV_X1 U2728 ( .A(n2716), .ZN(n2717) );
  INV_X1 U2729 ( .A(n3308), .ZN(n2718) );
  INV_X1 U2730 ( .A(n2718), .ZN(n2719) );
  INV_X1 U2731 ( .A(n3408), .ZN(n27201) );
  INV_X1 U2732 ( .A(n27201), .ZN(n2721) );
  INV_X1 U2733 ( .A(n970), .ZN(n2722) );
  CLKBUF_X1 U2734 ( .A(n2724), .Z(n2723) );
  CLKBUF_X1 U2735 ( .A(n37001), .Z(n2724) );
  INV_X1 U2736 ( .A(n1113), .ZN(n2725) );
  INV_X1 U2737 ( .A(n2725), .ZN(n2726) );
  INV_X1 U2738 ( .A(n2725), .ZN(n2727) );
  CLKBUF_X1 U2739 ( .A(n1764), .Z(n3385) );
  INV_X1 U2740 ( .A(n3385), .ZN(n2728) );
  INV_X1 U2741 ( .A(n3385), .ZN(n2729) );
  INV_X1 U2742 ( .A(n2095), .ZN(n27301) );
  INV_X1 U2743 ( .A(n27301), .ZN(n2731) );
  INV_X1 U2744 ( .A(n27301), .ZN(n2732) );
  CLKBUF_X1 U2745 ( .A(n1762), .Z(n3383) );
  INV_X1 U2746 ( .A(n3383), .ZN(n2733) );
  INV_X1 U2747 ( .A(n3383), .ZN(n2734) );
  INV_X1 U2748 ( .A(n1111), .ZN(n2735) );
  INV_X1 U2749 ( .A(n2735), .ZN(n2736) );
  INV_X1 U2750 ( .A(n2735), .ZN(n2737) );
  CLKBUF_X1 U2751 ( .A(n17601), .Z(n3381) );
  INV_X1 U2752 ( .A(n3381), .ZN(n2738) );
  INV_X1 U2753 ( .A(n3381), .ZN(n2739) );
  INV_X1 U2754 ( .A(n11101), .ZN(n27401) );
  INV_X1 U2755 ( .A(n27401), .ZN(n2741) );
  INV_X1 U2756 ( .A(n27401), .ZN(n2742) );
  INV_X1 U2757 ( .A(n1109), .ZN(n2743) );
  INV_X1 U2758 ( .A(n2743), .ZN(n2744) );
  INV_X1 U2759 ( .A(n2738), .ZN(n2745) );
  INV_X1 U2760 ( .A(n2745), .ZN(n2746) );
  INV_X1 U2761 ( .A(n2749), .ZN(n2747) );
  INV_X1 U2762 ( .A(n2747), .ZN(n2748) );
  CLKBUF_X1 U2763 ( .A(n20801), .Z(n3376) );
  INV_X1 U2764 ( .A(n3376), .ZN(n2749) );
  INV_X1 U2765 ( .A(n3376), .ZN(n27501) );
  INV_X1 U2766 ( .A(n4118), .ZN(n2751) );
  INV_X1 U2767 ( .A(n2751), .ZN(n2752) );
  CLKBUF_X1 U2768 ( .A(n1759), .Z(n3373) );
  INV_X1 U2769 ( .A(n3373), .ZN(n2753) );
  INV_X1 U2770 ( .A(n2757), .ZN(n2754) );
  INV_X1 U2771 ( .A(n2754), .ZN(n2755) );
  CLKBUF_X1 U2772 ( .A(n2757), .Z(n2756) );
  CLKBUF_X1 U2773 ( .A(n41401), .Z(n2757) );
  CLKBUF_X1 U2774 ( .A(n2759), .Z(n2758) );
  CLKBUF_X1 U2775 ( .A(n4139), .Z(n2759) );
  INV_X1 U2776 ( .A(n3371), .ZN(n27601) );
  INV_X1 U2777 ( .A(n27601), .ZN(n2761) );
  INV_X1 U2778 ( .A(n3369), .ZN(n2762) );
  INV_X1 U2779 ( .A(n2762), .ZN(n2763) );
  INV_X1 U2780 ( .A(n1753), .ZN(n2764) );
  INV_X1 U2781 ( .A(n2764), .ZN(n2765) );
  INV_X1 U2782 ( .A(n1749), .ZN(n2766) );
  INV_X1 U2783 ( .A(n2766), .ZN(n2767) );
  INV_X1 U2784 ( .A(n2073), .ZN(n2768) );
  INV_X1 U2785 ( .A(n2768), .ZN(n2769) );
  INV_X1 U2786 ( .A(n3365), .ZN(n27701) );
  INV_X1 U2787 ( .A(n27701), .ZN(n2771) );
  INV_X1 U2788 ( .A(n1737), .ZN(n2772) );
  INV_X1 U2789 ( .A(n2772), .ZN(n2773) );
  INV_X1 U2790 ( .A(n17401), .ZN(n2774) );
  INV_X1 U2791 ( .A(n2774), .ZN(n2775) );
  INV_X1 U2792 ( .A(n1731), .ZN(n2776) );
  INV_X1 U2793 ( .A(n2776), .ZN(n2777) );
  INV_X1 U2794 ( .A(n1734), .ZN(n2778) );
  INV_X1 U2795 ( .A(n2778), .ZN(n2779) );
  INV_X1 U2796 ( .A(n1725), .ZN(n27801) );
  INV_X1 U2797 ( .A(n27801), .ZN(n2781) );
  INV_X1 U2798 ( .A(n1728), .ZN(n2782) );
  INV_X1 U2799 ( .A(n2782), .ZN(n2783) );
  INV_X1 U2800 ( .A(n1719), .ZN(n2784) );
  INV_X1 U2801 ( .A(n2784), .ZN(n2785) );
  INV_X1 U2802 ( .A(n2784), .ZN(n2786) );
  INV_X1 U2803 ( .A(n1722), .ZN(n2787) );
  INV_X1 U2804 ( .A(n2787), .ZN(n2788) );
  INV_X1 U2805 ( .A(n17101), .ZN(n2789) );
  INV_X1 U2806 ( .A(n2789), .ZN(n27901) );
  INV_X1 U2807 ( .A(n1715), .ZN(n2791) );
  INV_X1 U2808 ( .A(n2791), .ZN(n2792) );
  INV_X1 U2809 ( .A(n1704), .ZN(n2793) );
  INV_X1 U2810 ( .A(n2793), .ZN(n2794) );
  INV_X1 U2811 ( .A(n1707), .ZN(n2795) );
  INV_X1 U2812 ( .A(n2795), .ZN(n2796) );
  INV_X1 U2813 ( .A(n1698), .ZN(n2797) );
  INV_X1 U2814 ( .A(n2797), .ZN(n2798) );
  INV_X1 U2815 ( .A(n1701), .ZN(n2799) );
  INV_X1 U2816 ( .A(n2799), .ZN(n28001) );
  INV_X1 U2817 ( .A(n1692), .ZN(n2801) );
  INV_X1 U2818 ( .A(n2801), .ZN(n2802) );
  INV_X1 U2819 ( .A(n1695), .ZN(n2803) );
  INV_X1 U2820 ( .A(n2803), .ZN(n2804) );
  INV_X1 U2821 ( .A(n1686), .ZN(n2805) );
  INV_X1 U2822 ( .A(n2805), .ZN(n2806) );
  INV_X1 U2823 ( .A(n1689), .ZN(n2807) );
  INV_X1 U2824 ( .A(n2807), .ZN(n2808) );
  INV_X1 U2825 ( .A(n16801), .ZN(n2809) );
  INV_X1 U2826 ( .A(n2809), .ZN(n28101) );
  INV_X1 U2827 ( .A(n1683), .ZN(n2811) );
  INV_X1 U2828 ( .A(n2811), .ZN(n2812) );
  INV_X1 U2829 ( .A(n1677), .ZN(n2813) );
  INV_X1 U2830 ( .A(n2813), .ZN(n2814) );
  INV_X1 U2831 ( .A(n1298), .ZN(n2815) );
  INV_X1 U2832 ( .A(n1298), .ZN(n2816) );
  INV_X1 U2833 ( .A(n1299), .ZN(n2817) );
  INV_X1 U2834 ( .A(n1299), .ZN(n2818) );
  INV_X1 U2835 ( .A(n13001), .ZN(n2819) );
  INV_X1 U2836 ( .A(n13001), .ZN(n28201) );
  INV_X1 U2837 ( .A(n1301), .ZN(n2821) );
  INV_X1 U2838 ( .A(n1301), .ZN(n2822) );
  INV_X1 U2839 ( .A(n1302), .ZN(n2823) );
  INV_X1 U2840 ( .A(n1302), .ZN(n2824) );
  INV_X1 U2841 ( .A(n1303), .ZN(n2825) );
  INV_X1 U2842 ( .A(n1303), .ZN(n2826) );
  INV_X1 U2843 ( .A(n1304), .ZN(n2827) );
  INV_X1 U2844 ( .A(n1304), .ZN(n2828) );
  INV_X1 U2845 ( .A(n1305), .ZN(n2829) );
  INV_X1 U2846 ( .A(n1305), .ZN(n28301) );
  INV_X1 U2847 ( .A(n1306), .ZN(n2831) );
  INV_X1 U2848 ( .A(n1306), .ZN(n2832) );
  INV_X1 U2849 ( .A(n1307), .ZN(n2833) );
  INV_X1 U2850 ( .A(n1307), .ZN(n2834) );
  INV_X1 U2851 ( .A(n1308), .ZN(n2835) );
  INV_X1 U2852 ( .A(n1308), .ZN(n2836) );
  INV_X1 U2853 ( .A(n1309), .ZN(n2837) );
  INV_X1 U2854 ( .A(n1309), .ZN(n2838) );
  INV_X1 U2855 ( .A(n13101), .ZN(n2839) );
  INV_X1 U2856 ( .A(n13101), .ZN(n28401) );
  INV_X1 U2857 ( .A(n1311), .ZN(n2841) );
  INV_X1 U2858 ( .A(n1311), .ZN(n2842) );
  INV_X1 U2859 ( .A(n1312), .ZN(n2843) );
  INV_X1 U2860 ( .A(n1312), .ZN(n2844) );
  INV_X1 U2861 ( .A(n1313), .ZN(n2845) );
  INV_X1 U2862 ( .A(n1313), .ZN(n2846) );
  INV_X1 U2863 ( .A(n1314), .ZN(n2847) );
  INV_X1 U2864 ( .A(n1314), .ZN(n2848) );
  INV_X1 U2865 ( .A(n1315), .ZN(n2849) );
  INV_X1 U2866 ( .A(n1315), .ZN(n28501) );
  INV_X1 U2867 ( .A(n1316), .ZN(n2851) );
  INV_X1 U2868 ( .A(n1316), .ZN(n2852) );
  INV_X1 U2869 ( .A(n1317), .ZN(n2853) );
  INV_X1 U2870 ( .A(n1317), .ZN(n2854) );
  INV_X1 U2871 ( .A(n1318), .ZN(n2855) );
  INV_X1 U2872 ( .A(n1318), .ZN(n2856) );
  INV_X1 U2873 ( .A(n1319), .ZN(n2857) );
  INV_X1 U2874 ( .A(n1319), .ZN(n2858) );
  INV_X1 U2875 ( .A(n13201), .ZN(n2859) );
  INV_X1 U2876 ( .A(n13201), .ZN(n28601) );
  INV_X1 U2877 ( .A(n1321), .ZN(n2861) );
  INV_X1 U2878 ( .A(n1321), .ZN(n2862) );
  INV_X1 U2879 ( .A(n1322), .ZN(n2863) );
  INV_X1 U2880 ( .A(n1322), .ZN(n2864) );
  INV_X1 U2881 ( .A(n1323), .ZN(n2865) );
  INV_X1 U2882 ( .A(n1323), .ZN(n2866) );
  INV_X1 U2883 ( .A(n1324), .ZN(n2867) );
  INV_X1 U2884 ( .A(n1324), .ZN(n2868) );
  INV_X1 U2885 ( .A(n1325), .ZN(n2869) );
  INV_X1 U2886 ( .A(n1325), .ZN(n28701) );
  INV_X1 U2887 ( .A(n1326), .ZN(n2871) );
  INV_X1 U2888 ( .A(n1326), .ZN(n2872) );
  INV_X1 U2889 ( .A(n1327), .ZN(n2873) );
  INV_X1 U2890 ( .A(n1327), .ZN(n2874) );
  INV_X1 U2891 ( .A(n1328), .ZN(n2875) );
  INV_X1 U2892 ( .A(n1328), .ZN(n2876) );
  INV_X1 U2893 ( .A(n1329), .ZN(n2877) );
  INV_X1 U2894 ( .A(n1329), .ZN(n2878) );
  INV_X1 U2895 ( .A(n13301), .ZN(n2879) );
  INV_X1 U2896 ( .A(n13301), .ZN(n28801) );
  INV_X1 U2897 ( .A(n1331), .ZN(n2881) );
  INV_X1 U2898 ( .A(n1331), .ZN(n2882) );
  INV_X1 U2899 ( .A(n1332), .ZN(n2883) );
  INV_X1 U2900 ( .A(n1332), .ZN(n2884) );
  INV_X1 U2901 ( .A(n1333), .ZN(n2885) );
  INV_X1 U2902 ( .A(n1333), .ZN(n2886) );
  INV_X1 U2903 ( .A(n1334), .ZN(n2887) );
  INV_X1 U2904 ( .A(n1334), .ZN(n2888) );
  INV_X1 U2905 ( .A(n1335), .ZN(n2889) );
  INV_X1 U2906 ( .A(n1335), .ZN(n28901) );
  INV_X1 U2907 ( .A(n1336), .ZN(n2891) );
  INV_X1 U2908 ( .A(n1336), .ZN(n2892) );
  INV_X1 U2909 ( .A(n1337), .ZN(n2893) );
  INV_X1 U2910 ( .A(n1337), .ZN(n2894) );
  INV_X1 U2911 ( .A(n1338), .ZN(n2895) );
  INV_X1 U2912 ( .A(n1338), .ZN(n2896) );
  INV_X1 U2913 ( .A(n1339), .ZN(n2897) );
  INV_X1 U2914 ( .A(n1339), .ZN(n2898) );
  INV_X1 U2915 ( .A(n13401), .ZN(n2899) );
  INV_X1 U2916 ( .A(n13401), .ZN(n29001) );
  INV_X1 U2917 ( .A(n1341), .ZN(n2901) );
  INV_X1 U2918 ( .A(n1341), .ZN(n29020) );
  INV_X1 U2919 ( .A(n1342), .ZN(n2903) );
  INV_X1 U2920 ( .A(n1342), .ZN(n2904) );
  INV_X1 U2921 ( .A(n1343), .ZN(n2905) );
  INV_X1 U2922 ( .A(n1343), .ZN(n2906) );
  INV_X1 U2923 ( .A(n1344), .ZN(n2907) );
  INV_X1 U2924 ( .A(n1344), .ZN(n2908) );
  INV_X1 U2925 ( .A(n1345), .ZN(n2909) );
  INV_X1 U2926 ( .A(n1345), .ZN(n29101) );
  INV_X1 U2927 ( .A(n1346), .ZN(n2911) );
  INV_X1 U2928 ( .A(n1346), .ZN(n2912) );
  INV_X1 U2929 ( .A(n659), .ZN(n2913) );
  INV_X1 U2930 ( .A(n659), .ZN(n2914) );
  CLKBUF_X1 U2931 ( .A(n2109), .Z(n3399) );
  INV_X1 U2932 ( .A(n3399), .ZN(n2915) );
  INV_X1 U2933 ( .A(n3399), .ZN(n2916) );
  INV_X1 U2934 ( .A(n1021), .ZN(n2917) );
  INV_X1 U2935 ( .A(n1021), .ZN(n2918) );
  INV_X1 U2936 ( .A(n1348), .ZN(n2919) );
  INV_X1 U2937 ( .A(n1348), .ZN(n29201) );
  INV_X1 U2938 ( .A(n1349), .ZN(n2921) );
  INV_X1 U2939 ( .A(n1349), .ZN(n2922) );
  INV_X1 U2940 ( .A(n13501), .ZN(n2923) );
  INV_X1 U2941 ( .A(n13501), .ZN(n2924) );
  CLKBUF_X1 U2942 ( .A(n2104), .Z(n3395) );
  INV_X1 U2943 ( .A(n3395), .ZN(n2925) );
  INV_X1 U2944 ( .A(n3395), .ZN(n2926) );
  INV_X1 U2945 ( .A(n2724), .ZN(n2927) );
  INV_X1 U2946 ( .A(n1352), .ZN(n2928) );
  INV_X1 U2947 ( .A(n1352), .ZN(n2929) );
  INV_X1 U2948 ( .A(n1353), .ZN(n29301) );
  INV_X1 U2949 ( .A(n1353), .ZN(n2931) );
  INV_X1 U2950 ( .A(n1354), .ZN(n2932) );
  INV_X1 U2951 ( .A(n1354), .ZN(n2933) );
  INV_X1 U2952 ( .A(n1355), .ZN(n2934) );
  INV_X1 U2953 ( .A(n1355), .ZN(n2935) );
  INV_X1 U2954 ( .A(n2091), .ZN(n2936) );
  INV_X1 U2955 ( .A(n1357), .ZN(n2937) );
  INV_X1 U2956 ( .A(n1357), .ZN(n2938) );
  INV_X1 U2957 ( .A(n1358), .ZN(n2939) );
  INV_X1 U2958 ( .A(n1358), .ZN(n29401) );
  INV_X1 U2959 ( .A(n578), .ZN(n2941) );
  INV_X1 U2960 ( .A(n578), .ZN(n2942) );
  INV_X1 U2961 ( .A(n13601), .ZN(n2943) );
  INV_X1 U2962 ( .A(n1363), .ZN(n2944) );
  INV_X1 U2963 ( .A(n1363), .ZN(n2945) );
  INV_X1 U2964 ( .A(n1367), .ZN(n2946) );
  INV_X1 U2965 ( .A(n13701), .ZN(n2947) );
  INV_X1 U2966 ( .A(n13701), .ZN(n2948) );
  INV_X1 U2967 ( .A(n39001), .ZN(n2949) );
  INV_X1 U2968 ( .A(n1372), .ZN(n29501) );
  INV_X1 U2969 ( .A(n1375), .ZN(n2951) );
  INV_X1 U2970 ( .A(n1375), .ZN(n2952) );
  INV_X1 U2971 ( .A(n3898), .ZN(n2953) );
  INV_X1 U2972 ( .A(n1379), .ZN(n2954) );
  INV_X1 U2973 ( .A(n1382), .ZN(n2955) );
  INV_X1 U2974 ( .A(n1382), .ZN(n2956) );
  INV_X1 U2975 ( .A(n3896), .ZN(n2957) );
  INV_X1 U2976 ( .A(n1386), .ZN(n2958) );
  INV_X1 U2977 ( .A(n1389), .ZN(n2959) );
  INV_X1 U2978 ( .A(n1389), .ZN(n29601) );
  INV_X1 U2979 ( .A(n3894), .ZN(n2961) );
  INV_X1 U2980 ( .A(n1393), .ZN(n2962) );
  INV_X1 U2981 ( .A(n1396), .ZN(n2963) );
  INV_X1 U2982 ( .A(n1396), .ZN(n2964) );
  INV_X1 U2983 ( .A(n3892), .ZN(n2965) );
  INV_X1 U2984 ( .A(n1398), .ZN(n2966) );
  INV_X1 U2985 ( .A(n1401), .ZN(n2967) );
  INV_X1 U2986 ( .A(n1401), .ZN(n2968) );
  INV_X1 U2987 ( .A(n38901), .ZN(n2969) );
  INV_X1 U2988 ( .A(n1403), .ZN(n29701) );
  INV_X1 U2989 ( .A(n1406), .ZN(n2971) );
  INV_X1 U2990 ( .A(n1406), .ZN(n2972) );
  INV_X1 U2991 ( .A(n3888), .ZN(n2973) );
  INV_X1 U2992 ( .A(n1408), .ZN(n2974) );
  INV_X1 U2993 ( .A(n1411), .ZN(n2975) );
  INV_X1 U2994 ( .A(n1411), .ZN(n2976) );
  INV_X1 U2995 ( .A(n3886), .ZN(n2977) );
  INV_X1 U2996 ( .A(n1415), .ZN(n2978) );
  INV_X1 U2997 ( .A(n1418), .ZN(n2979) );
  INV_X1 U2998 ( .A(n1418), .ZN(n29801) );
  INV_X1 U2999 ( .A(n3884), .ZN(n2981) );
  INV_X1 U3000 ( .A(n14201), .ZN(n2982) );
  INV_X1 U3001 ( .A(n1423), .ZN(n2983) );
  INV_X1 U3002 ( .A(n1423), .ZN(n2984) );
  INV_X1 U3003 ( .A(n3882), .ZN(n2985) );
  INV_X1 U3004 ( .A(n1427), .ZN(n2986) );
  INV_X1 U3005 ( .A(n14301), .ZN(n2987) );
  INV_X1 U3006 ( .A(n14301), .ZN(n2988) );
  INV_X1 U3007 ( .A(n38801), .ZN(n2989) );
  INV_X1 U3008 ( .A(n1434), .ZN(n29901) );
  INV_X1 U3009 ( .A(n1437), .ZN(n2991) );
  INV_X1 U3010 ( .A(n1437), .ZN(n2992) );
  INV_X1 U3011 ( .A(n3878), .ZN(n2993) );
  INV_X1 U3012 ( .A(n1441), .ZN(n2994) );
  INV_X1 U3013 ( .A(n1444), .ZN(n2995) );
  INV_X1 U3014 ( .A(n1444), .ZN(n2996) );
  INV_X1 U3015 ( .A(n3876), .ZN(n2997) );
  INV_X1 U3016 ( .A(n1446), .ZN(n2998) );
  INV_X1 U3017 ( .A(n1449), .ZN(n2999) );
  INV_X1 U3018 ( .A(n1449), .ZN(n30001) );
  INV_X1 U3019 ( .A(n3874), .ZN(n3001) );
  INV_X1 U3020 ( .A(n1453), .ZN(n3002) );
  INV_X1 U3021 ( .A(n1456), .ZN(n3003) );
  INV_X1 U3022 ( .A(n1456), .ZN(n3004) );
  INV_X1 U3023 ( .A(n3872), .ZN(n3005) );
  INV_X1 U3024 ( .A(n14601), .ZN(n3006) );
  INV_X1 U3025 ( .A(n1464), .ZN(n3007) );
  INV_X1 U3026 ( .A(n1467), .ZN(n3008) );
  INV_X1 U3027 ( .A(n2941), .ZN(n3711) );
  INV_X1 U3028 ( .A(n3711), .ZN(n3009) );
  INV_X1 U3029 ( .A(n2939), .ZN(n3709) );
  INV_X1 U3030 ( .A(n3709), .ZN(n30101) );
  INV_X1 U3031 ( .A(n1477), .ZN(n3011) );
  INV_X1 U3032 ( .A(n14801), .ZN(n3012) );
  INV_X1 U3033 ( .A(n1483), .ZN(n3013) );
  INV_X1 U3034 ( .A(n1486), .ZN(n3014) );
  CLKBUF_X1 U3035 ( .A(n2711), .Z(n3425) );
  INV_X1 U3036 ( .A(n3425), .ZN(n3015) );
  CLKBUF_X1 U3037 ( .A(n1773), .Z(n34001) );
  INV_X1 U3038 ( .A(n34001), .ZN(n3016) );
  INV_X1 U3039 ( .A(n34001), .ZN(n3017) );
  INV_X1 U3040 ( .A(n3401), .ZN(n3018) );
  INV_X1 U3041 ( .A(n3018), .ZN(n3019) );
  INV_X1 U3042 ( .A(n3018), .ZN(n30201) );
  INV_X1 U3043 ( .A(n33801), .ZN(n3021) );
  INV_X1 U3044 ( .A(n3021), .ZN(n3022) );
  INV_X1 U3045 ( .A(n3021), .ZN(n3023) );
  INV_X1 U3046 ( .A(n1497), .ZN(n3024) );
  INV_X1 U3047 ( .A(n15001), .ZN(n3025) );
  INV_X1 U3048 ( .A(n1503), .ZN(n3026) );
  INV_X1 U3049 ( .A(n2673), .ZN(n3027) );
  INV_X1 U3050 ( .A(n2674), .ZN(n3028) );
  INV_X1 U3051 ( .A(n2673), .ZN(n3029) );
  INV_X1 U3052 ( .A(n2674), .ZN(n30301) );
  INV_X1 U3053 ( .A(n2675), .ZN(n3031) );
  INV_X1 U3054 ( .A(n2676), .ZN(n3032) );
  INV_X1 U3055 ( .A(n2675), .ZN(n3033) );
  INV_X1 U3056 ( .A(n2676), .ZN(n3034) );
  INV_X1 U3057 ( .A(n2669), .ZN(n3035) );
  INV_X1 U3058 ( .A(n26701), .ZN(n3036) );
  INV_X1 U3059 ( .A(n2669), .ZN(n3037) );
  INV_X1 U3060 ( .A(n26701), .ZN(n3038) );
  INV_X1 U3061 ( .A(n2671), .ZN(n3039) );
  INV_X1 U3062 ( .A(n2672), .ZN(n30401) );
  INV_X1 U3063 ( .A(n2671), .ZN(n3041) );
  INV_X1 U3064 ( .A(n2672), .ZN(n3042) );
  INV_X1 U3065 ( .A(n2665), .ZN(n3043) );
  INV_X1 U3066 ( .A(n2666), .ZN(n3044) );
  INV_X1 U3067 ( .A(n2665), .ZN(n3045) );
  INV_X1 U3068 ( .A(n2666), .ZN(n3046) );
  INV_X1 U3069 ( .A(n2667), .ZN(n3047) );
  INV_X1 U3070 ( .A(n2668), .ZN(n3048) );
  INV_X1 U3071 ( .A(n2667), .ZN(n3049) );
  INV_X1 U3072 ( .A(n2668), .ZN(n30501) );
  INV_X1 U3073 ( .A(n2661), .ZN(n3051) );
  INV_X1 U3074 ( .A(n2662), .ZN(n3052) );
  INV_X1 U3075 ( .A(n2661), .ZN(n3053) );
  INV_X1 U3076 ( .A(n2662), .ZN(n3054) );
  INV_X1 U3077 ( .A(n2663), .ZN(n3055) );
  INV_X1 U3078 ( .A(n2664), .ZN(n3056) );
  INV_X1 U3079 ( .A(n2663), .ZN(n3057) );
  INV_X1 U3080 ( .A(n2664), .ZN(n3058) );
  INV_X1 U3081 ( .A(n2657), .ZN(n3059) );
  INV_X1 U3082 ( .A(n2658), .ZN(n30601) );
  INV_X1 U3083 ( .A(n2657), .ZN(n3061) );
  INV_X1 U3084 ( .A(n2658), .ZN(n3062) );
  INV_X1 U3085 ( .A(n2659), .ZN(n3063) );
  INV_X1 U3086 ( .A(n26601), .ZN(n3064) );
  INV_X1 U3087 ( .A(n2659), .ZN(n3065) );
  INV_X1 U3088 ( .A(n26601), .ZN(n3066) );
  INV_X1 U3089 ( .A(n2653), .ZN(n3067) );
  INV_X1 U3090 ( .A(n2654), .ZN(n3068) );
  INV_X1 U3091 ( .A(n2653), .ZN(n3069) );
  INV_X1 U3092 ( .A(n2654), .ZN(n30701) );
  INV_X1 U3093 ( .A(n2655), .ZN(n3071) );
  INV_X1 U3094 ( .A(n2656), .ZN(n3072) );
  INV_X1 U3095 ( .A(n2655), .ZN(n3073) );
  INV_X1 U3096 ( .A(n2656), .ZN(n3074) );
  INV_X1 U3097 ( .A(n2649), .ZN(n3075) );
  INV_X1 U3098 ( .A(n26501), .ZN(n3076) );
  INV_X1 U3099 ( .A(n2649), .ZN(n3077) );
  INV_X1 U3100 ( .A(n26501), .ZN(n3078) );
  INV_X1 U3101 ( .A(n2651), .ZN(n3079) );
  INV_X1 U3102 ( .A(n2652), .ZN(n30801) );
  INV_X1 U3103 ( .A(n2651), .ZN(n3081) );
  INV_X1 U3104 ( .A(n2652), .ZN(n3082) );
  INV_X1 U3105 ( .A(n2645), .ZN(n3083) );
  INV_X1 U3106 ( .A(n2646), .ZN(n3084) );
  INV_X1 U3107 ( .A(n2645), .ZN(n3085) );
  INV_X1 U3108 ( .A(n2646), .ZN(n3086) );
  INV_X1 U3109 ( .A(n2647), .ZN(n3087) );
  INV_X1 U3110 ( .A(n2648), .ZN(n3088) );
  INV_X1 U3111 ( .A(n2647), .ZN(n3089) );
  INV_X1 U3112 ( .A(n2648), .ZN(n30901) );
  INV_X1 U3113 ( .A(n2641), .ZN(n3091) );
  INV_X1 U3114 ( .A(n2642), .ZN(n3092) );
  INV_X1 U3115 ( .A(n2642), .ZN(n3093) );
  INV_X1 U3116 ( .A(n2641), .ZN(n3094) );
  INV_X1 U3117 ( .A(n2643), .ZN(n3095) );
  INV_X1 U3118 ( .A(n2644), .ZN(n3096) );
  INV_X1 U3119 ( .A(n2644), .ZN(n3097) );
  INV_X1 U3120 ( .A(n2643), .ZN(n3098) );
  INV_X1 U3121 ( .A(n2638), .ZN(n3099) );
  INV_X1 U3122 ( .A(n2638), .ZN(n31001) );
  INV_X1 U3123 ( .A(n2637), .ZN(n3101) );
  INV_X1 U3124 ( .A(n2637), .ZN(n3102) );
  INV_X1 U3125 ( .A(n2639), .ZN(n3103) );
  INV_X1 U3126 ( .A(n26401), .ZN(n3104) );
  INV_X1 U3127 ( .A(n26401), .ZN(n3105) );
  INV_X1 U3128 ( .A(n2639), .ZN(n3106) );
  INV_X1 U3129 ( .A(n2633), .ZN(n3107) );
  INV_X1 U3130 ( .A(n2634), .ZN(n3108) );
  INV_X1 U3131 ( .A(n2634), .ZN(n3109) );
  INV_X1 U3132 ( .A(n2633), .ZN(n31101) );
  INV_X1 U3133 ( .A(n2635), .ZN(n3111) );
  INV_X1 U3134 ( .A(n2636), .ZN(n3112) );
  INV_X1 U3135 ( .A(n2636), .ZN(n3113) );
  INV_X1 U3136 ( .A(n2635), .ZN(n3114) );
  INV_X1 U3137 ( .A(n26301), .ZN(n3115) );
  INV_X1 U3138 ( .A(n26301), .ZN(n3116) );
  INV_X1 U3139 ( .A(n2629), .ZN(n3117) );
  INV_X1 U3140 ( .A(n2629), .ZN(n3118) );
  INV_X1 U3141 ( .A(n2631), .ZN(n3119) );
  INV_X1 U3142 ( .A(n2632), .ZN(n31201) );
  INV_X1 U3143 ( .A(n2632), .ZN(n3121) );
  INV_X1 U3144 ( .A(n2631), .ZN(n3122) );
  INV_X1 U3145 ( .A(n2625), .ZN(n3123) );
  INV_X1 U3146 ( .A(n2626), .ZN(n3124) );
  INV_X1 U3147 ( .A(n2626), .ZN(n3125) );
  INV_X1 U3148 ( .A(n2625), .ZN(n3126) );
  INV_X1 U3149 ( .A(n2627), .ZN(n3127) );
  INV_X1 U3150 ( .A(n2628), .ZN(n3128) );
  INV_X1 U3151 ( .A(n2628), .ZN(n3129) );
  INV_X1 U3152 ( .A(n2627), .ZN(n31301) );
  INV_X1 U3153 ( .A(n2622), .ZN(n3131) );
  INV_X1 U3154 ( .A(n2622), .ZN(n3132) );
  INV_X1 U3155 ( .A(n2621), .ZN(n3133) );
  INV_X1 U3156 ( .A(n2621), .ZN(n3134) );
  INV_X1 U3157 ( .A(n2623), .ZN(n3135) );
  INV_X1 U3158 ( .A(n2624), .ZN(n3136) );
  INV_X1 U3159 ( .A(n2624), .ZN(n3137) );
  INV_X1 U3160 ( .A(n2623), .ZN(n3138) );
  INV_X1 U3161 ( .A(n2617), .ZN(n3139) );
  INV_X1 U3162 ( .A(n2618), .ZN(n31401) );
  INV_X1 U3163 ( .A(n2618), .ZN(n3141) );
  INV_X1 U3164 ( .A(n2617), .ZN(n3142) );
  INV_X1 U3165 ( .A(n2619), .ZN(n3143) );
  INV_X1 U3166 ( .A(n26201), .ZN(n3144) );
  INV_X1 U3167 ( .A(n26201), .ZN(n3145) );
  INV_X1 U3168 ( .A(n2619), .ZN(n3146) );
  INV_X1 U3169 ( .A(n2613), .ZN(n3147) );
  INV_X1 U3170 ( .A(n2614), .ZN(n3148) );
  INV_X1 U3171 ( .A(n2613), .ZN(n3149) );
  INV_X1 U3172 ( .A(n2614), .ZN(n31501) );
  INV_X1 U3173 ( .A(n2615), .ZN(n3151) );
  INV_X1 U3174 ( .A(n2616), .ZN(n3152) );
  INV_X1 U3175 ( .A(n2616), .ZN(n3153) );
  INV_X1 U3176 ( .A(n2615), .ZN(n3154) );
  INV_X1 U3177 ( .A(n1126), .ZN(n3155) );
  INV_X1 U3178 ( .A(n11201), .ZN(n3156) );
  INV_X1 U3179 ( .A(n3156), .ZN(n3157) );
  INV_X1 U3180 ( .A(n3156), .ZN(n3158) );
  INV_X1 U3181 ( .A(n26101), .ZN(n3159) );
  INV_X1 U3182 ( .A(n2609), .ZN(n31601) );
  INV_X1 U3183 ( .A(n26101), .ZN(n3161) );
  INV_X1 U3184 ( .A(n2609), .ZN(n3162) );
  INV_X1 U3185 ( .A(n2612), .ZN(n3163) );
  INV_X1 U3186 ( .A(n2611), .ZN(n3164) );
  INV_X1 U3187 ( .A(n2612), .ZN(n3165) );
  INV_X1 U3188 ( .A(n2611), .ZN(n3166) );
  INV_X1 U3189 ( .A(n558), .ZN(n3167) );
  INV_X1 U3190 ( .A(n2606), .ZN(n3168) );
  INV_X1 U3191 ( .A(n2605), .ZN(n3169) );
  INV_X1 U3192 ( .A(n2606), .ZN(n31701) );
  INV_X1 U3193 ( .A(n2605), .ZN(n3171) );
  INV_X1 U3194 ( .A(n2608), .ZN(n3172) );
  INV_X1 U3195 ( .A(n2607), .ZN(n3173) );
  INV_X1 U3196 ( .A(n2608), .ZN(n3174) );
  INV_X1 U3197 ( .A(n2607), .ZN(n3175) );
  INV_X1 U3198 ( .A(n3704), .ZN(n3176) );
  INV_X1 U3199 ( .A(n1116), .ZN(n3177) );
  INV_X1 U3200 ( .A(n3177), .ZN(n3178) );
  INV_X1 U3201 ( .A(n3177), .ZN(n3179) );
  INV_X1 U3202 ( .A(n1128), .ZN(n4474) );
  INV_X1 U3203 ( .A(n2602), .ZN(n31801) );
  INV_X1 U3204 ( .A(n2601), .ZN(n3181) );
  INV_X1 U3205 ( .A(n2602), .ZN(n3182) );
  INV_X1 U3206 ( .A(n2601), .ZN(n3183) );
  INV_X1 U3207 ( .A(n2603), .ZN(n3184) );
  INV_X1 U3208 ( .A(n2604), .ZN(n3185) );
  INV_X1 U3209 ( .A(n2603), .ZN(n3186) );
  INV_X1 U3210 ( .A(n2604), .ZN(n3187) );
  INV_X1 U3211 ( .A(n2719), .ZN(n3188) );
  INV_X1 U3212 ( .A(n3188), .ZN(n3189) );
  INV_X1 U3213 ( .A(n3189), .ZN(n31901) );
  INV_X1 U3214 ( .A(n3189), .ZN(n3191) );
  INV_X1 U3215 ( .A(n2177), .ZN(n4338) );
  INV_X1 U3216 ( .A(n2598), .ZN(n3192) );
  INV_X1 U3217 ( .A(n2597), .ZN(n3193) );
  INV_X1 U3218 ( .A(n2598), .ZN(n3194) );
  INV_X1 U3219 ( .A(n2597), .ZN(n3195) );
  INV_X1 U3220 ( .A(n26001), .ZN(n3196) );
  INV_X1 U3221 ( .A(n2599), .ZN(n3197) );
  INV_X1 U3222 ( .A(n26001), .ZN(n3198) );
  INV_X1 U3223 ( .A(n2599), .ZN(n3199) );
  INV_X1 U3224 ( .A(n2722), .ZN(n32001) );
  INV_X1 U3225 ( .A(n32001), .ZN(n3201) );
  INV_X1 U3226 ( .A(n3201), .ZN(n3202) );
  INV_X1 U3227 ( .A(n3201), .ZN(n3203) );
  INV_X1 U3228 ( .A(n2678), .ZN(n4202) );
  INV_X1 U3229 ( .A(n2594), .ZN(n3204) );
  INV_X1 U3230 ( .A(n2593), .ZN(n3205) );
  INV_X1 U3231 ( .A(n2594), .ZN(n3206) );
  INV_X1 U3232 ( .A(n2593), .ZN(n3207) );
  INV_X1 U3233 ( .A(n2596), .ZN(n3208) );
  INV_X1 U3234 ( .A(n2595), .ZN(n3209) );
  INV_X1 U3235 ( .A(n2596), .ZN(n32101) );
  INV_X1 U3236 ( .A(n2595), .ZN(n3211) );
  INV_X1 U3237 ( .A(n2589), .ZN(n3212) );
  INV_X1 U3238 ( .A(n25901), .ZN(n3213) );
  INV_X1 U3239 ( .A(n2589), .ZN(n3214) );
  INV_X1 U3240 ( .A(n25901), .ZN(n3215) );
  INV_X1 U3241 ( .A(n2145), .ZN(n3421) );
  INV_X1 U3242 ( .A(n2591), .ZN(n3216) );
  INV_X1 U3243 ( .A(n2591), .ZN(n3217) );
  INV_X1 U3244 ( .A(n2592), .ZN(n3218) );
  INV_X1 U3245 ( .A(n2592), .ZN(n3219) );
  INV_X1 U3246 ( .A(n2584), .ZN(n32201) );
  INV_X1 U3247 ( .A(n2585), .ZN(n3221) );
  INV_X1 U3248 ( .A(n2584), .ZN(n3222) );
  INV_X1 U3249 ( .A(n2585), .ZN(n3223) );
  INV_X1 U3250 ( .A(n2912), .ZN(n3224) );
  INV_X1 U3251 ( .A(n1019), .ZN(n3225) );
  CLKBUF_X1 U3252 ( .A(n1769), .Z(n3226) );
  INV_X1 U3253 ( .A(n25801), .ZN(n3227) );
  INV_X1 U3254 ( .A(n2581), .ZN(n3228) );
  INV_X1 U3255 ( .A(n25801), .ZN(n3229) );
  INV_X1 U3256 ( .A(n2581), .ZN(n32301) );
  INV_X1 U3257 ( .A(n2583), .ZN(n3231) );
  INV_X1 U3258 ( .A(n2582), .ZN(n3232) );
  INV_X1 U3259 ( .A(n2583), .ZN(n3233) );
  INV_X1 U3260 ( .A(n2577), .ZN(n3234) );
  INV_X1 U3261 ( .A(n2577), .ZN(n3235) );
  INV_X1 U3262 ( .A(n2579), .ZN(n3236) );
  INV_X1 U3263 ( .A(n2579), .ZN(n3237) );
  INV_X1 U3264 ( .A(n2578), .ZN(n3238) );
  INV_X1 U3265 ( .A(n2575), .ZN(n3239) );
  INV_X1 U3266 ( .A(n2575), .ZN(n32401) );
  INV_X1 U3267 ( .A(n2576), .ZN(n3241) );
  INV_X1 U3268 ( .A(n576), .ZN(n3242) );
  INV_X1 U3269 ( .A(n1203), .ZN(n3243) );
  INV_X1 U3270 ( .A(n27101), .ZN(n3244) );
  INV_X1 U3271 ( .A(n3419), .ZN(n3245) );
  INV_X1 U3272 ( .A(n3245), .ZN(n3246) );
  INV_X1 U3273 ( .A(n3245), .ZN(n3247) );
  INV_X1 U3274 ( .A(n2574), .ZN(n3248) );
  INV_X1 U3275 ( .A(n2573), .ZN(n3249) );
  INV_X1 U3276 ( .A(n2566), .ZN(n32501) );
  INV_X1 U3277 ( .A(n2565), .ZN(n3251) );
  INV_X1 U3278 ( .A(n1208), .ZN(n3252) );
  INV_X1 U3279 ( .A(n2715), .ZN(n3253) );
  INV_X1 U3280 ( .A(n3417), .ZN(n3254) );
  INV_X1 U3281 ( .A(n3254), .ZN(n3255) );
  INV_X1 U3282 ( .A(n3254), .ZN(n3256) );
  INV_X1 U3283 ( .A(n2561), .ZN(n3257) );
  INV_X1 U3284 ( .A(n2562), .ZN(n3258) );
  INV_X1 U3285 ( .A(n2564), .ZN(n3259) );
  INV_X1 U3286 ( .A(n2563), .ZN(n32601) );
  INV_X1 U3287 ( .A(n2559), .ZN(n3261) );
  INV_X1 U3288 ( .A(n25601), .ZN(n3262) );
  INV_X1 U3289 ( .A(n1205), .ZN(n3263) );
  INV_X1 U3290 ( .A(n1206), .ZN(n3264) );
  CLKBUF_X1 U3291 ( .A(n3432), .Z(n3265) );
  INV_X1 U3292 ( .A(n2158), .ZN(n3432) );
  INV_X1 U3293 ( .A(n1212), .ZN(n3266) );
  INV_X1 U3294 ( .A(n2717), .ZN(n3267) );
  INV_X1 U3295 ( .A(n2557), .ZN(n3268) );
  INV_X1 U3296 ( .A(n2558), .ZN(n3269) );
  INV_X1 U3297 ( .A(n25501), .ZN(n32701) );
  INV_X1 U3298 ( .A(n25501), .ZN(n3271) );
  INV_X1 U3299 ( .A(n2551), .ZN(n3272) );
  INV_X1 U3300 ( .A(n2551), .ZN(n3273) );
  INV_X1 U3301 ( .A(n2552), .ZN(n3274) );
  INV_X1 U3302 ( .A(n2553), .ZN(n3275) );
  INV_X1 U3303 ( .A(n2549), .ZN(n3276) );
  INV_X1 U3304 ( .A(n2548), .ZN(n3277) );
  INV_X1 U3305 ( .A(n3706), .ZN(n3278) );
  INV_X1 U3306 ( .A(n3278), .ZN(n3279) );
  INV_X1 U3307 ( .A(n915), .ZN(n32801) );
  INV_X1 U3308 ( .A(n915), .ZN(n3281) );
  INV_X1 U3309 ( .A(n2545), .ZN(n3282) );
  INV_X1 U3310 ( .A(n2546), .ZN(n3283) );
  INV_X1 U3311 ( .A(n2546), .ZN(n3284) );
  INV_X1 U3312 ( .A(n2547), .ZN(n3285) );
  INV_X1 U3313 ( .A(n2547), .ZN(n3286) );
  INV_X1 U3314 ( .A(n25401), .ZN(n3287) );
  INV_X1 U3315 ( .A(n2541), .ZN(n3288) );
  INV_X1 U3316 ( .A(n25401), .ZN(n3289) );
  INV_X1 U3317 ( .A(n2541), .ZN(n32901) );
  INV_X1 U3318 ( .A(n2542), .ZN(n3291) );
  INV_X1 U3319 ( .A(n2542), .ZN(n3292) );
  INV_X1 U3320 ( .A(n911), .ZN(n3293) );
  INV_X1 U3321 ( .A(n912), .ZN(n3294) );
  INV_X1 U3322 ( .A(n911), .ZN(n3295) );
  INV_X1 U3323 ( .A(n2538), .ZN(n3296) );
  INV_X1 U3324 ( .A(n2538), .ZN(n3297) );
  INV_X1 U3325 ( .A(n2539), .ZN(n3298) );
  INV_X1 U3326 ( .A(n2533), .ZN(n3299) );
  INV_X1 U3327 ( .A(n2532), .ZN(n33001) );
  INV_X1 U3328 ( .A(n2532), .ZN(n3301) );
  INV_X1 U3329 ( .A(n2533), .ZN(n3302) );
  INV_X1 U3330 ( .A(n2528), .ZN(n3303) );
  INV_X1 U3331 ( .A(n2527), .ZN(n3304) );
  INV_X1 U3332 ( .A(n2527), .ZN(n3305) );
  INV_X1 U3333 ( .A(n2528), .ZN(n3306) );
  INV_X1 U3334 ( .A(n2525), .ZN(n3307) );
  INV_X1 U3335 ( .A(n2525), .ZN(n3308) );
  INV_X1 U3336 ( .A(n2526), .ZN(n3309) );
  INV_X1 U3337 ( .A(n2526), .ZN(n33101) );
  INV_X1 U3338 ( .A(n2685), .ZN(n3311) );
  INV_X1 U3339 ( .A(n1063), .ZN(n3312) );
  INV_X1 U3340 ( .A(n3703), .ZN(n3313) );
  INV_X1 U3341 ( .A(n3904), .ZN(n3314) );
  INV_X1 U3342 ( .A(n3868), .ZN(n3315) );
  INV_X1 U3343 ( .A(n4403), .ZN(n3316) );
  INV_X1 U3344 ( .A(n3761), .ZN(n3317) );
  INV_X1 U3345 ( .A(n2265), .ZN(n3318) );
  INV_X1 U3346 ( .A(n2266), .ZN(n3319) );
  INV_X1 U3347 ( .A(n2265), .ZN(n33201) );
  INV_X1 U3348 ( .A(n2266), .ZN(n3321) );
  INV_X1 U3349 ( .A(n1619), .ZN(n3322) );
  INV_X1 U3350 ( .A(n1622), .ZN(n3323) );
  INV_X1 U3351 ( .A(n16250), .ZN(n3324) );
  INV_X1 U3352 ( .A(n16280), .ZN(n3325) );
  INV_X1 U3353 ( .A(n16310), .ZN(n3326) );
  INV_X1 U3354 ( .A(n16340), .ZN(n3327) );
  INV_X1 U3355 ( .A(n16370), .ZN(n3328) );
  INV_X1 U3356 ( .A(n16401), .ZN(n3329) );
  INV_X1 U3357 ( .A(n1643), .ZN(n33301) );
  INV_X1 U3358 ( .A(n1646), .ZN(n3331) );
  INV_X1 U3359 ( .A(n1649), .ZN(n3332) );
  INV_X1 U3360 ( .A(n1652), .ZN(n3333) );
  INV_X1 U3361 ( .A(n1655), .ZN(n3334) );
  INV_X1 U3362 ( .A(n1658), .ZN(n3335) );
  INV_X1 U3363 ( .A(n1661), .ZN(n3336) );
  INV_X1 U3364 ( .A(n1664), .ZN(n3337) );
  INV_X1 U3365 ( .A(n1667), .ZN(n3338) );
  INV_X1 U3366 ( .A(n16701), .ZN(n3339) );
  INV_X1 U3367 ( .A(n1673), .ZN(n33401) );
  INV_X1 U3368 ( .A(n1676), .ZN(n3341) );
  INV_X1 U3369 ( .A(n1679), .ZN(n3342) );
  INV_X1 U3370 ( .A(n1682), .ZN(n3343) );
  INV_X1 U3371 ( .A(n1685), .ZN(n3344) );
  INV_X1 U3372 ( .A(n1688), .ZN(n3345) );
  INV_X1 U3373 ( .A(n1691), .ZN(n3346) );
  INV_X1 U3374 ( .A(n1694), .ZN(n3347) );
  INV_X1 U3375 ( .A(n1697), .ZN(n3348) );
  INV_X1 U3376 ( .A(n17001), .ZN(n3349) );
  INV_X1 U3377 ( .A(n1703), .ZN(n33501) );
  INV_X1 U3378 ( .A(n1706), .ZN(n3351) );
  INV_X1 U3379 ( .A(n1709), .ZN(n3352) );
  INV_X1 U3380 ( .A(n4267), .ZN(n3353) );
  INV_X1 U3381 ( .A(n1713), .ZN(n3354) );
  INV_X1 U3382 ( .A(n1714), .ZN(n3355) );
  INV_X1 U3383 ( .A(n3714), .ZN(n3356) );
  INV_X1 U3384 ( .A(n1718), .ZN(n3357) );
  INV_X1 U3385 ( .A(n1721), .ZN(n3358) );
  INV_X1 U3386 ( .A(n1724), .ZN(n3359) );
  INV_X1 U3387 ( .A(n1727), .ZN(n33601) );
  INV_X1 U3388 ( .A(n17301), .ZN(n3361) );
  INV_X1 U3389 ( .A(n1733), .ZN(n3362) );
  INV_X1 U3390 ( .A(n1736), .ZN(n3363) );
  INV_X1 U3391 ( .A(n1739), .ZN(n3364) );
  INV_X1 U3392 ( .A(n1743), .ZN(n3365) );
  INV_X1 U3393 ( .A(n1743), .ZN(n3366) );
  INV_X1 U3394 ( .A(n3718), .ZN(n3367) );
  INV_X1 U3395 ( .A(n1748), .ZN(n3368) );
  INV_X1 U3396 ( .A(n1751), .ZN(n3369) );
  INV_X1 U3397 ( .A(n1751), .ZN(n33701) );
  INV_X1 U3398 ( .A(n1755), .ZN(n3371) );
  INV_X1 U3399 ( .A(n1755), .ZN(n3372) );
  INV_X1 U3400 ( .A(n1759), .ZN(n3374) );
  INV_X1 U3401 ( .A(n20801), .ZN(n3375) );
  INV_X1 U3402 ( .A(n2081), .ZN(n3377) );
  INV_X1 U3403 ( .A(n2081), .ZN(n3378) );
  INV_X1 U3404 ( .A(n1204), .ZN(n3379) );
  CLKBUF_X1 U3405 ( .A(n43401), .Z(n33801) );
  INV_X1 U3406 ( .A(n1263), .ZN(n43401) );
  INV_X1 U3407 ( .A(n17601), .ZN(n3382) );
  INV_X1 U3408 ( .A(n1762), .ZN(n3384) );
  INV_X1 U3409 ( .A(n1764), .ZN(n3386) );
  INV_X1 U3410 ( .A(n2677), .ZN(n3387) );
  INV_X1 U3411 ( .A(n1766), .ZN(n3388) );
  INV_X1 U3412 ( .A(n2912), .ZN(n3389) );
  INV_X1 U3413 ( .A(n2103), .ZN(n33901) );
  INV_X1 U3414 ( .A(n2102), .ZN(n3391) );
  INV_X1 U3415 ( .A(n2103), .ZN(n3392) );
  INV_X1 U3416 ( .A(n2102), .ZN(n3393) );
  INV_X1 U3417 ( .A(n2105), .ZN(n3394) );
  INV_X1 U3418 ( .A(n2105), .ZN(n3396) );
  INV_X1 U3419 ( .A(n21101), .ZN(n3397) );
  INV_X1 U3420 ( .A(n21101), .ZN(n3398) );
  INV_X1 U3421 ( .A(n1773), .ZN(n3401) );
  INV_X1 U3422 ( .A(n1774), .ZN(n3402) );
  INV_X1 U3423 ( .A(n1774), .ZN(n3403) );
  INV_X1 U3424 ( .A(n1219), .ZN(n3404) );
  INV_X1 U3425 ( .A(n2722), .ZN(n3405) );
  INV_X1 U3426 ( .A(n1213), .ZN(n3406) );
  INV_X1 U3427 ( .A(n2719), .ZN(n3407) );
  INV_X1 U3428 ( .A(n1785), .ZN(n3408) );
  INV_X1 U3429 ( .A(n1785), .ZN(n3409) );
  INV_X1 U3430 ( .A(n12101), .ZN(n34101) );
  INV_X1 U3431 ( .A(n558), .ZN(n3411) );
  INV_X1 U3432 ( .A(n2717), .ZN(n3412) );
  INV_X1 U3433 ( .A(n2712), .ZN(n3413) );
  INV_X1 U3434 ( .A(n2712), .ZN(n3414) );
  INV_X1 U3435 ( .A(n3301), .ZN(n3415) );
  INV_X1 U3436 ( .A(n1208), .ZN(n3416) );
  INV_X1 U3437 ( .A(n2715), .ZN(n3417) );
  INV_X1 U3438 ( .A(n1203), .ZN(n3418) );
  INV_X1 U3439 ( .A(n27101), .ZN(n3419) );
  INV_X1 U3440 ( .A(matrix_index[0]), .ZN(n34201) );
  INV_X1 U3441 ( .A(n2146), .ZN(n3422) );
  INV_X1 U3442 ( .A(n2146), .ZN(n3423) );
  INV_X1 U3443 ( .A(n1204), .ZN(n3426) );
  INV_X1 U3444 ( .A(n2711), .ZN(n3427) );
  INV_X1 U3445 ( .A(n1769), .ZN(n3428) );
  INV_X1 U3446 ( .A(n1019), .ZN(n3429) );
  INV_X1 U3447 ( .A(matrix_index[2]), .ZN(n34301) );
  INV_X1 U3448 ( .A(n2159), .ZN(n3431) );
  INV_X1 U3449 ( .A(n1794), .ZN(n3433) );
  INV_X1 U3450 ( .A(n1794), .ZN(n3434) );
  BUF_X1 U3451 ( .A(n4128), .Z(n3435) );
  AND2_X1 U3452 ( .A1(n1603), .A2(n3438), .ZN(n4061) );
  BUF_X1 U3453 ( .A(n2941), .Z(n3436) );
  BUF_X1 U3454 ( .A(n2942), .Z(n3437) );
  BUF_X1 U3455 ( .A(n4059), .Z(n3438) );
  BUF_X1 U3456 ( .A(n4094), .Z(n3439) );
  NOR2_X1 U3457 ( .A1(n1247), .A2(n3457), .ZN(n4062) );
  INV_X1 U3458 ( .A(n4062), .ZN(n34401) );
  INV_X1 U3459 ( .A(n4062), .ZN(n3441) );
  OR3_X1 U3460 ( .A1(n2697), .A2(n3242), .A3(n2759), .ZN(n4197) );
  INV_X1 U3461 ( .A(n4197), .ZN(n3442) );
  INV_X1 U3462 ( .A(n4197), .ZN(n3443) );
  BUF_X1 U3463 ( .A(n2939), .Z(n3444) );
  BUF_X1 U3464 ( .A(n10301), .Z(n3445) );
  INV_X1 U3465 ( .A(n15400), .ZN(n3468) );
  NAND2_X1 U3466 ( .A1(n3227), .A2(n18001), .ZN(n3907) );
  NAND2_X1 U3467 ( .A1(n32301), .A2(n3903), .ZN(n3871) );
  NAND2_X1 U3468 ( .A1(n4675), .A2(n4001), .ZN(n4679) );
  NAND2_X1 U3469 ( .A1(n4125), .A2(n3439), .ZN(n4127) );
  NAND2_X1 U3470 ( .A1(n582), .A2(n4119), .ZN(n4098) );
  AND2_X1 U3471 ( .A1(n1296), .A2(n26801), .ZN(n4137) );
  AND2_X1 U3472 ( .A1(n582), .A2(n1801), .ZN(n41001) );
  NOR3_X1 U3473 ( .A1(n3447), .A2(n3448), .A3(n3449), .ZN(n3446) );
  NAND3_X1 U3474 ( .A1(n581), .A2(n1137), .A3(n1602), .ZN(n4123) );
  NOR2_X1 U3475 ( .A1(n2691), .A2(n1527), .ZN(n3715) );
  NAND2_X1 U3476 ( .A1(n3228), .A2(n3966), .ZN(n3942) );
  NAND2_X1 U3477 ( .A1(n32301), .A2(n2217), .ZN(n3967) );
  AND2_X1 U3478 ( .A1(n1297), .A2(n585), .ZN(n4134) );
  AND2_X1 U3479 ( .A1(n554), .A2(n1291), .ZN(n4135) );
  INV_X1 U3480 ( .A(n3795), .ZN(n3761) );
  INV_X1 U3481 ( .A(n4604), .ZN(n4538) );
  INV_X1 U3482 ( .A(n4469), .ZN(n4403) );
  INV_X1 U3483 ( .A(n4333), .ZN(n4264) );
  INV_X1 U3484 ( .A(n3902), .ZN(n3868) );
  INV_X1 U3485 ( .A(n3938), .ZN(n3904) );
  AND2_X1 U3486 ( .A1(n1296), .A2(n1294), .ZN(n4136) );
  INV_X1 U3487 ( .A(n3757), .ZN(n3723) );
  INV_X1 U3488 ( .A(n3537), .ZN(n3693) );
  INV_X1 U3489 ( .A(n3538), .ZN(n36901) );
  INV_X1 U3490 ( .A(n3539), .ZN(n3687) );
  INV_X1 U3491 ( .A(n35401), .ZN(n3684) );
  INV_X1 U3492 ( .A(n3541), .ZN(n3681) );
  INV_X1 U3493 ( .A(n3542), .ZN(n3678) );
  INV_X1 U3494 ( .A(n3543), .ZN(n3675) );
  INV_X1 U3495 ( .A(n3544), .ZN(n3672) );
  INV_X1 U3496 ( .A(n3545), .ZN(n3669) );
  INV_X1 U3497 ( .A(n3546), .ZN(n3666) );
  INV_X1 U3498 ( .A(n3547), .ZN(n3663) );
  INV_X1 U3499 ( .A(n3548), .ZN(n36601) );
  INV_X1 U3500 ( .A(n3549), .ZN(n3657) );
  INV_X1 U3501 ( .A(n35501), .ZN(n3654) );
  INV_X1 U3502 ( .A(n3551), .ZN(n3651) );
  INV_X1 U3503 ( .A(n3552), .ZN(n3696) );
  INV_X1 U3504 ( .A(n3584), .ZN(n3647) );
  INV_X1 U3505 ( .A(n3553), .ZN(n3624) );
  INV_X1 U3506 ( .A(n3555), .ZN(n3622) );
  INV_X1 U3507 ( .A(n3557), .ZN(n36201) );
  INV_X1 U3508 ( .A(n3559), .ZN(n3618) );
  INV_X1 U3509 ( .A(n3561), .ZN(n3646) );
  INV_X1 U3510 ( .A(n3563), .ZN(n3644) );
  INV_X1 U3511 ( .A(n3565), .ZN(n3642) );
  INV_X1 U3512 ( .A(n3567), .ZN(n36401) );
  INV_X1 U3513 ( .A(n3569), .ZN(n3638) );
  INV_X1 U3514 ( .A(n3571), .ZN(n3636) );
  INV_X1 U3515 ( .A(n3573), .ZN(n3634) );
  INV_X1 U3516 ( .A(n3575), .ZN(n3632) );
  INV_X1 U3517 ( .A(n3577), .ZN(n36301) );
  INV_X1 U3518 ( .A(n3579), .ZN(n3628) );
  INV_X1 U3519 ( .A(n3581), .ZN(n3626) );
  INV_X1 U3520 ( .A(n3583), .ZN(n3648) );
  INV_X1 U3521 ( .A(n1131), .ZN(n4142) );
  BUF_X1 U3522 ( .A(n4198), .Z(n3697) );
  BUF_X1 U3523 ( .A(n4198), .Z(n3698) );
  BUF_X1 U3524 ( .A(n29401), .Z(n37101) );
  BUF_X1 U3525 ( .A(n1128), .Z(n3703) );
  BUF_X1 U3526 ( .A(n1129), .Z(n3704) );
  XNOR2_X1 U3527 ( .A(n3455), .B(r317_carry_2_), .ZN(N1539) );
  XNOR2_X1 U3528 ( .A(n1795), .B(n3472), .ZN(n3447) );
  NAND2_X1 U3529 ( .A1(n1795), .A2(n3453), .ZN(n3472) );
  XOR2_X1 U3530 ( .A(n1796), .B(n3453), .Z(n3448) );
  XOR2_X1 U3531 ( .A(n3461), .B(n3456), .Z(n3449) );
  XNOR2_X1 U3532 ( .A(n34601), .B(n3451), .ZN(n3471) );
  XNOR2_X1 U3533 ( .A(n3459), .B(r317_carry_3_), .ZN(n34701) );
  AND2_X1 U3534 ( .A1(n1121), .A2(n3452), .ZN(n34501) );
  AND2_X1 U3535 ( .A1(n3459), .A2(r317_carry_3_), .ZN(n3451) );
  AND2_X1 U3536 ( .A1(n1186), .A2(n3712), .ZN(n3452) );
  AND2_X1 U3537 ( .A1(n3461), .A2(n3456), .ZN(n3453) );
  XOR2_X1 U3538 ( .A(n2214), .B(n3712), .Z(n3454) );
  XOR2_X1 U3539 ( .A(n1121), .B(n3452), .Z(n3455) );
  AND2_X1 U3540 ( .A1(n34601), .A2(n3451), .ZN(n3456) );
  OR2_X1 U3541 ( .A1(n3455), .A2(r317_carry_2_), .ZN(r317_carry_3_) );
  AND3_X1 U3542 ( .A1(n577), .A2(n1798), .A3(n4093), .ZN(n3457) );
  NAND2_X1 U3543 ( .A1(n4683), .A2(n4681), .ZN(N100) );
  NAND2_X1 U3544 ( .A1(n46801), .A2(n588), .ZN(N102) );
  INV_X1 U3545 ( .A(n3474), .ZN(n3691) );
  INV_X1 U3546 ( .A(n3476), .ZN(n3688) );
  INV_X1 U3547 ( .A(n3478), .ZN(n3685) );
  INV_X1 U3548 ( .A(n34801), .ZN(n3682) );
  INV_X1 U3549 ( .A(n3482), .ZN(n3679) );
  INV_X1 U3550 ( .A(n3484), .ZN(n3676) );
  INV_X1 U3551 ( .A(n3486), .ZN(n3673) );
  INV_X1 U3552 ( .A(n3488), .ZN(n36701) );
  INV_X1 U3553 ( .A(n34901), .ZN(n3667) );
  INV_X1 U3554 ( .A(n3492), .ZN(n3664) );
  INV_X1 U3555 ( .A(n3494), .ZN(n3661) );
  INV_X1 U3556 ( .A(n3496), .ZN(n3658) );
  INV_X1 U3557 ( .A(n3498), .ZN(n3655) );
  INV_X1 U3558 ( .A(n35001), .ZN(n3652) );
  INV_X1 U3559 ( .A(n3502), .ZN(n3649) );
  INV_X1 U3560 ( .A(n3504), .ZN(n3694) );
  INV_X1 U3561 ( .A(n3554), .ZN(n3623) );
  INV_X1 U3562 ( .A(n3556), .ZN(n3621) );
  INV_X1 U3563 ( .A(n3558), .ZN(n3619) );
  INV_X1 U3564 ( .A(n35601), .ZN(n3617) );
  INV_X1 U3565 ( .A(n3562), .ZN(n3645) );
  INV_X1 U3566 ( .A(n3564), .ZN(n3643) );
  INV_X1 U3567 ( .A(n3566), .ZN(n3641) );
  INV_X1 U3568 ( .A(n3568), .ZN(n3639) );
  INV_X1 U3569 ( .A(n35701), .ZN(n3637) );
  INV_X1 U3570 ( .A(n3572), .ZN(n3635) );
  INV_X1 U3571 ( .A(n3574), .ZN(n3633) );
  INV_X1 U3572 ( .A(n3576), .ZN(n3631) );
  INV_X1 U3573 ( .A(n3578), .ZN(n3629) );
  INV_X1 U3574 ( .A(n35801), .ZN(n3627) );
  INV_X1 U3575 ( .A(n3582), .ZN(n3625) );
  INV_X1 U3576 ( .A(n3586), .ZN(n3692) );
  INV_X1 U3577 ( .A(n3588), .ZN(n3689) );
  INV_X1 U3578 ( .A(n35901), .ZN(n3686) );
  INV_X1 U3579 ( .A(n3592), .ZN(n3683) );
  INV_X1 U3580 ( .A(n3594), .ZN(n36801) );
  INV_X1 U3581 ( .A(n3596), .ZN(n3677) );
  INV_X1 U3582 ( .A(n3598), .ZN(n3674) );
  INV_X1 U3583 ( .A(n36001), .ZN(n3671) );
  INV_X1 U3584 ( .A(n3602), .ZN(n3668) );
  INV_X1 U3585 ( .A(n3604), .ZN(n3665) );
  INV_X1 U3586 ( .A(n3606), .ZN(n3662) );
  INV_X1 U3587 ( .A(n3608), .ZN(n3659) );
  INV_X1 U3588 ( .A(n36101), .ZN(n3656) );
  INV_X1 U3589 ( .A(n3612), .ZN(n3653) );
  INV_X1 U3590 ( .A(n3614), .ZN(n36501) );
  INV_X1 U3591 ( .A(n3616), .ZN(n3695) );
  NAND2_X1 U3592 ( .A1(n1288), .A2(n4119), .ZN(n4267) );
  AND2_X1 U3593 ( .A1(n585), .A2(n10201), .ZN(n4611) );
  BUF_X1 U3594 ( .A(n2677), .Z(n37001) );
  BUF_X1 U3595 ( .A(n2678), .Z(n3701) );
  BUF_X1 U3596 ( .A(n4118), .Z(n3707) );
  BUF_X1 U3597 ( .A(n2178), .Z(n3699) );
  OR2_X1 U3598 ( .A1(n3454), .A2(n32201), .ZN(r317_carry_2_) );
  INV_X1 U3599 ( .A(n3422), .ZN(n3712) );
  AND2_X1 U3600 ( .A1(n580), .A2(n34501), .ZN(n3458) );
  XOR2_X1 U3601 ( .A(n2697), .B(n34501), .Z(n3459) );
  XOR2_X1 U3602 ( .A(n1463), .B(n3458), .Z(n34601) );
  XOR2_X1 U3603 ( .A(n3468), .B(n3462), .Z(n3461) );
  AND2_X1 U3604 ( .A1(n1465), .A2(n3458), .ZN(n3462) );
  AND2_X1 U3605 ( .A1(n1193), .A2(n3462), .ZN(n3463) );
  INV_X1 U3606 ( .A(r298_carry_5_), .ZN(n3469) );
  XOR2_X1 U3607 ( .A(n543), .B(n37), .Z(n3464) );
  XOR2_X1 U3608 ( .A(n15400), .B(n3467), .Z(n3465) );
  XNOR2_X1 U3609 ( .A(n541), .B(n37), .ZN(N1228) );
  XNOR2_X1 U3610 ( .A(n15510), .B(r298_carry_5_), .ZN(N1229) );
  OR2_X1 U3611 ( .A1(n542), .A2(n547), .ZN(r298_carry_5_) );
  AND2_X1 U3612 ( .A1(n1193), .A2(n3469), .ZN(n3466) );
  INV_X1 U3613 ( .A(n545), .ZN(r290_B_3_) );
  AND2_X1 U3614 ( .A1(n542), .A2(n35), .ZN(n3467) );
  MUX2_X1 U3615 ( .A(n21700), .B(n537), .S(n1543), .Z(n3473) );
  MUX2_X1 U3616 ( .A(n37800), .B(n45700), .S(n3263), .Z(n3474) );
  MUX2_X1 U3617 ( .A(n3693), .B(n3473), .S(n2119), .Z(N1623) );
  MUX2_X1 U3618 ( .A(n21300), .B(n532), .S(n15530), .Z(n3475) );
  MUX2_X1 U3619 ( .A(n37400), .B(n45200), .S(n3274), .Z(n3476) );
  MUX2_X1 U3620 ( .A(n36901), .B(n3475), .S(n850), .Z(N1624) );
  MUX2_X1 U3621 ( .A(n20900), .B(n527), .S(n21401), .Z(n3477) );
  MUX2_X1 U3622 ( .A(n37000), .B(n44700), .S(n3268), .Z(n3478) );
  MUX2_X1 U3623 ( .A(n3687), .B(n3477), .S(n3218), .Z(N1625) );
  MUX2_X1 U3624 ( .A(n20500), .B(n522), .S(n3256), .Z(n3479) );
  MUX2_X1 U3625 ( .A(n36600), .B(n44200), .S(n2556), .Z(n34801) );
  MUX2_X1 U3626 ( .A(n3684), .B(n3479), .S(n3215), .Z(N1626) );
  MUX2_X1 U3627 ( .A(n20100), .B(n517), .S(n3247), .Z(n3481) );
  MUX2_X1 U3628 ( .A(n36200), .B(n43700), .S(n3261), .Z(n3482) );
  MUX2_X1 U3629 ( .A(n3681), .B(n3481), .S(n30201), .Z(N1627) );
  MUX2_X1 U3630 ( .A(n19700), .B(n512), .S(n15490), .Z(n3483) );
  MUX2_X1 U3631 ( .A(n35800), .B(n43200), .S(n3267), .Z(n3484) );
  MUX2_X1 U3632 ( .A(n3678), .B(n3483), .S(n2257), .Z(N1628) );
  MUX2_X1 U3633 ( .A(n19300), .B(n507), .S(n1545), .Z(n3485) );
  MUX2_X1 U3634 ( .A(n35400), .B(n42700), .S(n1564), .Z(n3486) );
  MUX2_X1 U3635 ( .A(n3675), .B(n3485), .S(n2116), .Z(N1629) );
  MUX2_X1 U3636 ( .A(n18900), .B(n5020), .S(n15511), .Z(n3487) );
  MUX2_X1 U3637 ( .A(n35000), .B(n42200), .S(n1565), .Z(n3488) );
  MUX2_X1 U3638 ( .A(n3672), .B(n3487), .S(n3223), .Z(N1630) );
  MUX2_X1 U3639 ( .A(n18500), .B(n497), .S(n2143), .Z(n3489) );
  MUX2_X1 U3640 ( .A(n34600), .B(n41700), .S(n3272), .Z(n34901) );
  MUX2_X1 U3641 ( .A(n3669), .B(n3489), .S(n2254), .Z(N1631) );
  MUX2_X1 U3642 ( .A(n18100), .B(n4920), .S(n2137), .Z(n3491) );
  MUX2_X1 U3643 ( .A(n34200), .B(n41200), .S(n3264), .Z(n3492) );
  MUX2_X1 U3644 ( .A(n3666), .B(n3491), .S(n1498), .Z(N1632) );
  MUX2_X1 U3645 ( .A(n17700), .B(n4870), .S(n15390), .Z(n3493) );
  MUX2_X1 U3646 ( .A(n33800), .B(n40700), .S(n15701), .Z(n3494) );
  MUX2_X1 U3647 ( .A(n3663), .B(n3493), .S(n1217), .Z(N1633) );
  MUX2_X1 U3648 ( .A(n17300), .B(n4820), .S(n2569), .Z(n3495) );
  MUX2_X1 U3649 ( .A(n33400), .B(n40200), .S(n2122), .Z(n3496) );
  MUX2_X1 U3650 ( .A(n36601), .B(n3495), .S(n22601), .Z(N1634) );
  MUX2_X1 U3651 ( .A(n16900), .B(n4770), .S(n1541), .Z(n3497) );
  MUX2_X1 U3652 ( .A(n33000), .B(n39700), .S(n3414), .Z(n3498) );
  MUX2_X1 U3653 ( .A(n3657), .B(n3497), .S(n3219), .Z(N1635) );
  MUX2_X1 U3654 ( .A(n16500), .B(n4720), .S(n15470), .Z(n3499) );
  MUX2_X1 U3655 ( .A(n32600), .B(n39200), .S(n15580), .Z(n35001) );
  MUX2_X1 U3656 ( .A(n3654), .B(n3499), .S(n3403), .Z(N1636) );
  MUX2_X1 U3657 ( .A(n16100), .B(n46700), .S(n2572), .Z(n3501) );
  MUX2_X1 U3658 ( .A(n32200), .B(n38700), .S(n2128), .Z(n3502) );
  MUX2_X1 U3659 ( .A(n3651), .B(n3501), .S(n1218), .Z(N1637) );
  MUX2_X1 U3660 ( .A(n15700), .B(n46200), .S(n2134), .Z(n3503) );
  MUX2_X1 U3661 ( .A(n31800), .B(n38200), .S(n3266), .Z(n3504) );
  MUX2_X1 U3662 ( .A(n3696), .B(n3503), .S(n3017), .Z(N1638) );
  MUX2_X1 U3663 ( .A(n3623), .B(n3693), .S(n2257), .Z(N1581) );
  MUX2_X1 U3664 ( .A(n3621), .B(n36901), .S(n3214), .Z(N1582) );
  MUX2_X1 U3665 ( .A(n3619), .B(n3687), .S(n3019), .Z(N1583) );
  MUX2_X1 U3666 ( .A(n3617), .B(n3684), .S(n2259), .Z(N1584) );
  MUX2_X1 U3667 ( .A(n3645), .B(n3681), .S(n3222), .Z(N1585) );
  MUX2_X1 U3668 ( .A(n3643), .B(n3678), .S(n3024), .Z(N1586) );
  MUX2_X1 U3669 ( .A(n3641), .B(n3675), .S(n2253), .Z(N1587) );
  MUX2_X1 U3670 ( .A(n3639), .B(n3672), .S(n1522), .Z(N1588) );
  MUX2_X1 U3671 ( .A(n3637), .B(n3669), .S(n3217), .Z(N1589) );
  MUX2_X1 U3672 ( .A(n3635), .B(n3666), .S(n22601), .Z(N1590) );
  MUX2_X1 U3673 ( .A(n3633), .B(n3663), .S(n3401), .Z(N1591) );
  MUX2_X1 U3674 ( .A(n3631), .B(n36601), .S(n557), .Z(N1592) );
  MUX2_X1 U3675 ( .A(n3629), .B(n3657), .S(n1523), .Z(N1593) );
  MUX2_X1 U3676 ( .A(n3627), .B(n3654), .S(n2256), .Z(N1594) );
  MUX2_X1 U3677 ( .A(n3625), .B(n3651), .S(n2254), .Z(N1595) );
  MUX2_X1 U3678 ( .A(n3647), .B(n3696), .S(n2115), .Z(N1596) );
  MUX2_X1 U3679 ( .A(n3692), .B(n3623), .S(n2118), .Z(N1547) );
  MUX2_X1 U3680 ( .A(n3689), .B(n3621), .S(n30201), .Z(N1548) );
  MUX2_X1 U3681 ( .A(n3686), .B(n3619), .S(n1523), .Z(N1549) );
  MUX2_X1 U3682 ( .A(n3683), .B(n3617), .S(n1057), .Z(N1550) );
  MUX2_X1 U3683 ( .A(n36801), .B(n3645), .S(n3213), .Z(N1551) );
  MUX2_X1 U3684 ( .A(n3677), .B(n3643), .S(n3216), .Z(N1552) );
  MUX2_X1 U3685 ( .A(n3674), .B(n3641), .S(n3016), .Z(N1553) );
  MUX2_X1 U3686 ( .A(n3671), .B(n3639), .S(n3221), .Z(N1554) );
  MUX2_X1 U3687 ( .A(n3668), .B(n3637), .S(n2116), .Z(N1555) );
  MUX2_X1 U3688 ( .A(n3665), .B(n3635), .S(n1115), .Z(N1556) );
  MUX2_X1 U3689 ( .A(n3662), .B(n3633), .S(n1499), .Z(N1557) );
  MUX2_X1 U3690 ( .A(n3659), .B(n3631), .S(n3219), .Z(N1558) );
  MUX2_X1 U3691 ( .A(n3656), .B(n3629), .S(n1218), .Z(N1559) );
  MUX2_X1 U3692 ( .A(n3653), .B(n3627), .S(n1114), .Z(N1560) );
  MUX2_X1 U3693 ( .A(n36501), .B(n3625), .S(n3017), .Z(N1561) );
  MUX2_X1 U3694 ( .A(n3695), .B(n3647), .S(n3024), .Z(N1562) );
  MUX2_X1 U3695 ( .A(n3), .B(n21800), .S(n15550), .Z(n3505) );
  MUX2_X1 U3696 ( .A(n3505), .B(n3624), .S(n3246), .Z(n3506) );
  MUX2_X1 U3697 ( .A(n3506), .B(n3692), .S(n3212), .Z(N924) );
  MUX2_X1 U3698 ( .A(n4), .B(n21400), .S(n1567), .Z(n3507) );
  MUX2_X1 U3699 ( .A(n3507), .B(n3622), .S(n2133), .Z(n3508) );
  MUX2_X1 U3700 ( .A(n3508), .B(n3689), .S(n1498), .Z(N925) );
  MUX2_X1 U3701 ( .A(n5), .B(n21000), .S(n15590), .Z(n3509) );
  MUX2_X1 U3702 ( .A(n3509), .B(n36201), .S(n1119), .Z(n35101) );
  MUX2_X1 U3703 ( .A(n35101), .B(n3686), .S(n32201), .Z(N926) );
  MUX2_X1 U3704 ( .A(n6), .B(n20600), .S(n2556), .Z(n3511) );
  MUX2_X1 U3705 ( .A(n3511), .B(n3618), .S(n3253), .Z(n3512) );
  MUX2_X1 U3706 ( .A(n3512), .B(n3683), .S(n3218), .Z(N927) );
  MUX2_X1 U3707 ( .A(n7), .B(n20200), .S(n3263), .Z(n3513) );
  MUX2_X1 U3708 ( .A(n3513), .B(n3646), .S(n3251), .Z(n3514) );
  MUX2_X1 U3709 ( .A(n3514), .B(n36801), .S(n2119), .Z(N928) );
  MUX2_X1 U3710 ( .A(n8), .B(n19800), .S(n3267), .Z(n3515) );
  MUX2_X1 U3711 ( .A(n3515), .B(n3644), .S(n3259), .Z(n3516) );
  MUX2_X1 U3712 ( .A(n3516), .B(n3677), .S(n1522), .Z(N929) );
  MUX2_X1 U3713 ( .A(n9), .B(n19400), .S(n15610), .Z(n3517) );
  MUX2_X1 U3714 ( .A(n3517), .B(n3642), .S(n3249), .Z(n3518) );
  MUX2_X1 U3715 ( .A(n3518), .B(n3674), .S(n3402), .Z(N930) );
  MUX2_X1 U3716 ( .A(n10), .B(n19000), .S(n1565), .Z(n3519) );
  MUX2_X1 U3717 ( .A(n3519), .B(n36401), .S(n3257), .Z(n35201) );
  MUX2_X1 U3718 ( .A(n35201), .B(n3671), .S(n2115), .Z(N931) );
  MUX2_X1 U3719 ( .A(n11), .B(n18600), .S(n3262), .Z(n3521) );
  MUX2_X1 U3720 ( .A(n3521), .B(n3638), .S(n32501), .Z(n3522) );
  MUX2_X1 U3721 ( .A(n3522), .B(n3668), .S(n2256), .Z(N932) );
  MUX2_X1 U3722 ( .A(n12), .B(n18200), .S(n2122), .Z(n3523) );
  MUX2_X1 U3723 ( .A(n3523), .B(n3636), .S(n32601), .Z(n3524) );
  MUX2_X1 U3724 ( .A(n3524), .B(n3665), .S(n3215), .Z(N933) );
  MUX2_X1 U3725 ( .A(n13), .B(n17800), .S(n3414), .Z(n3525) );
  MUX2_X1 U3726 ( .A(n3525), .B(n3634), .S(n2139), .Z(n3526) );
  MUX2_X1 U3727 ( .A(n3526), .B(n3662), .S(n1057), .Z(N934) );
  MUX2_X1 U3728 ( .A(n14), .B(n17400), .S(n3271), .Z(n3527) );
  MUX2_X1 U3729 ( .A(n3527), .B(n3632), .S(n1118), .Z(n3528) );
  MUX2_X1 U3730 ( .A(n3528), .B(n3659), .S(n2253), .Z(N935) );
  MUX2_X1 U3731 ( .A(n15), .B(n17000), .S(n3269), .Z(n3529) );
  MUX2_X1 U3732 ( .A(n3529), .B(n36301), .S(n3244), .Z(n35301) );
  MUX2_X1 U3733 ( .A(n35301), .B(n3656), .S(n3217), .Z(N936) );
  MUX2_X1 U3734 ( .A(n16), .B(n16600), .S(n1791), .Z(n3531) );
  MUX2_X1 U3735 ( .A(n3531), .B(n3628), .S(n3258), .Z(n3532) );
  MUX2_X1 U3736 ( .A(n3532), .B(n3653), .S(n3223), .Z(N937) );
  MUX2_X1 U3737 ( .A(n17), .B(n16200), .S(n2128), .Z(n3533) );
  MUX2_X1 U3738 ( .A(n3533), .B(n3626), .S(n3248), .Z(n3534) );
  MUX2_X1 U3739 ( .A(n3534), .B(n36501), .S(n2259), .Z(N938) );
  MUX2_X1 U3740 ( .A(n26900), .B(n15800), .S(n3275), .Z(n3535) );
  MUX2_X1 U3741 ( .A(n3535), .B(n3648), .S(n3255), .Z(n3536) );
  MUX2_X1 U3742 ( .A(n3536), .B(n3695), .S(n3019), .Z(N939) );
  MUX2_X1 U3743 ( .A(n3691), .B(n825), .S(n15401), .Z(n3537) );
  MUX2_X1 U3744 ( .A(n3688), .B(n824), .S(n3417), .Z(n3538) );
  MUX2_X1 U3745 ( .A(n3685), .B(n823), .S(n2142), .Z(n3539) );
  MUX2_X1 U3746 ( .A(n3682), .B(n822), .S(n15520), .Z(n35401) );
  MUX2_X1 U3747 ( .A(n3679), .B(n821), .S(n1542), .Z(n3541) );
  MUX2_X1 U3748 ( .A(n3676), .B(n820), .S(n3416), .Z(n3542) );
  MUX2_X1 U3749 ( .A(n3673), .B(n819), .S(n3418), .Z(n3543) );
  MUX2_X1 U3750 ( .A(n36701), .B(n818), .S(n15540), .Z(n3544) );
  MUX2_X1 U3751 ( .A(n3667), .B(n817), .S(n3419), .Z(n3545) );
  MUX2_X1 U3752 ( .A(n3664), .B(n816), .S(n15480), .Z(n3546) );
  MUX2_X1 U3753 ( .A(n3661), .B(n815), .S(n1544), .Z(n3547) );
  MUX2_X1 U3754 ( .A(n3658), .B(n814), .S(n15500), .Z(n3548) );
  MUX2_X1 U3755 ( .A(n3655), .B(n813), .S(n2571), .Z(n3549) );
  MUX2_X1 U3756 ( .A(n3652), .B(n812), .S(n2568), .Z(n35501) );
  MUX2_X1 U3757 ( .A(n3649), .B(n811), .S(n1546), .Z(n3551) );
  MUX2_X1 U3758 ( .A(n3694), .B(n810), .S(n2136), .Z(n3552) );
  MUX2_X1 U3759 ( .A(n2817), .B(n1364), .S(n1566), .Z(n3553) );
  MUX2_X1 U3760 ( .A(n3553), .B(n39001), .S(n3249), .Z(n3554) );
  MUX2_X1 U3761 ( .A(n2815), .B(n3961), .S(n1117), .Z(n3555) );
  MUX2_X1 U3762 ( .A(n3555), .B(n3898), .S(n3259), .Z(n3556) );
  MUX2_X1 U3763 ( .A(n2821), .B(n1376), .S(n3269), .Z(n3557) );
  MUX2_X1 U3764 ( .A(n3557), .B(n3896), .S(n3247), .Z(n3558) );
  MUX2_X1 U3765 ( .A(n2819), .B(n1383), .S(n1566), .Z(n3559) );
  MUX2_X1 U3766 ( .A(n3559), .B(n3894), .S(n32601), .Z(n35601) );
  MUX2_X1 U3767 ( .A(n2825), .B(n13901), .S(n3262), .Z(n3561) );
  MUX2_X1 U3768 ( .A(n3561), .B(n3892), .S(n32501), .Z(n3562) );
  MUX2_X1 U3769 ( .A(n2823), .B(n3956), .S(n3275), .Z(n3563) );
  MUX2_X1 U3770 ( .A(n3563), .B(n38901), .S(n2134), .Z(n3564) );
  MUX2_X1 U3771 ( .A(n2829), .B(n3954), .S(n21301), .Z(n3565) );
  MUX2_X1 U3772 ( .A(n3565), .B(n3888), .S(n3243), .Z(n3566) );
  MUX2_X1 U3773 ( .A(n2827), .B(n3952), .S(n1568), .Z(n3567) );
  MUX2_X1 U3774 ( .A(n3567), .B(n3886), .S(n3258), .Z(n3568) );
  MUX2_X1 U3775 ( .A(n2833), .B(n1412), .S(n15620), .Z(n3569) );
  MUX2_X1 U3776 ( .A(n3569), .B(n3884), .S(n21401), .Z(n35701) );
  MUX2_X1 U3777 ( .A(n2831), .B(n3949), .S(n3412), .Z(n3571) );
  MUX2_X1 U3778 ( .A(n3571), .B(n3882), .S(n3244), .Z(n3572) );
  MUX2_X1 U3779 ( .A(n2837), .B(n1424), .S(n15560), .Z(n3573) );
  MUX2_X1 U3780 ( .A(n3573), .B(n38801), .S(n3251), .Z(n3574) );
  MUX2_X1 U3781 ( .A(n2835), .B(n1431), .S(n1792), .Z(n3575) );
  MUX2_X1 U3782 ( .A(n3575), .B(n3878), .S(n3248), .Z(n3576) );
  MUX2_X1 U3783 ( .A(n2841), .B(n1438), .S(n15600), .Z(n3577) );
  MUX2_X1 U3784 ( .A(n3577), .B(n3876), .S(n3257), .Z(n3578) );
  MUX2_X1 U3785 ( .A(n2839), .B(n3944), .S(n2124), .Z(n3579) );
  MUX2_X1 U3786 ( .A(n3579), .B(n3874), .S(n3253), .Z(n35801) );
  MUX2_X1 U3787 ( .A(n2845), .B(n14501), .S(n3413), .Z(n3581) );
  MUX2_X1 U3788 ( .A(n3581), .B(n3872), .S(n3256), .Z(n3582) );
  MUX2_X1 U3789 ( .A(n2843), .B(n1457), .S(n32701), .Z(n3583) );
  MUX2_X1 U3790 ( .A(n3583), .B(n3869), .S(n3252), .Z(n3584) );
  MUX2_X1 U3791 ( .A(n3793), .B(n825), .S(n2127), .Z(n3585) );
  MUX2_X1 U3792 ( .A(n3585), .B(n3691), .S(n2139), .Z(n3586) );
  MUX2_X1 U3793 ( .A(n3791), .B(n824), .S(n2555), .Z(n3587) );
  MUX2_X1 U3794 ( .A(n3587), .B(n3688), .S(n2133), .Z(n3588) );
  MUX2_X1 U3795 ( .A(n3789), .B(n823), .S(n15631), .Z(n3589) );
  MUX2_X1 U3796 ( .A(n3589), .B(n3685), .S(n2572), .Z(n35901) );
  MUX2_X1 U3797 ( .A(n3787), .B(n822), .S(n3273), .Z(n3591) );
  MUX2_X1 U3798 ( .A(n3591), .B(n3682), .S(n2137), .Z(n3592) );
  MUX2_X1 U3799 ( .A(n3785), .B(n821), .S(n15570), .Z(n3593) );
  MUX2_X1 U3800 ( .A(n3593), .B(n3679), .S(n1543), .Z(n3594) );
  MUX2_X1 U3801 ( .A(n3783), .B(n820), .S(n1569), .Z(n3595) );
  MUX2_X1 U3802 ( .A(n3595), .B(n3676), .S(n15511), .Z(n3596) );
  MUX2_X1 U3803 ( .A(n3781), .B(n819), .S(n3264), .Z(n3597) );
  MUX2_X1 U3804 ( .A(n3597), .B(n3673), .S(n15390), .Z(n3598) );
  MUX2_X1 U3805 ( .A(n3779), .B(n818), .S(n3274), .Z(n3599) );
  MUX2_X1 U3806 ( .A(n3599), .B(n36701), .S(n15470), .Z(n36001) );
  MUX2_X1 U3807 ( .A(n3777), .B(n817), .S(n3268), .Z(n3601) );
  MUX2_X1 U3808 ( .A(n3601), .B(n3667), .S(n1545), .Z(n3602) );
  MUX2_X1 U3809 ( .A(n3775), .B(n816), .S(n3266), .Z(n3603) );
  MUX2_X1 U3810 ( .A(n3603), .B(n3664), .S(n15530), .Z(n3604) );
  MUX2_X1 U3811 ( .A(n3773), .B(n815), .S(n3261), .Z(n3605) );
  MUX2_X1 U3812 ( .A(n3605), .B(n3661), .S(n3246), .Z(n3606) );
  MUX2_X1 U3813 ( .A(n3771), .B(n814), .S(n2125), .Z(n3607) );
  MUX2_X1 U3814 ( .A(n3607), .B(n3658), .S(n2569), .Z(n3608) );
  MUX2_X1 U3815 ( .A(n3769), .B(n813), .S(n920), .Z(n3609) );
  MUX2_X1 U3816 ( .A(n3609), .B(n3655), .S(n2143), .Z(n36101) );
  MUX2_X1 U3817 ( .A(n3767), .B(n812), .S(n2121), .Z(n3611) );
  MUX2_X1 U3818 ( .A(n3611), .B(n3652), .S(n15490), .Z(n3612) );
  MUX2_X1 U3819 ( .A(n3765), .B(n811), .S(n2131), .Z(n3613) );
  MUX2_X1 U3820 ( .A(n3613), .B(n3649), .S(n1541), .Z(n3614) );
  MUX2_X1 U3821 ( .A(n3762), .B(n810), .S(n3272), .Z(n3615) );
  MUX2_X1 U3822 ( .A(n3615), .B(n3694), .S(n3255), .Z(n3616) );
  NAND2_X1 U3823 ( .A1(n1292), .A2(n1031), .ZN(n3702) );
  AND2_X1 U3824 ( .A1(n1293), .A2(n2943), .ZN(n3705) );
  AND2_X1 U3825 ( .A1(n1294), .A2(n1362), .ZN(n3706) );
  NAND2_X1 U3826 ( .A1(n1289), .A2(n1801), .ZN(n3708) );
  INV_X1 U3827 ( .A(n3713), .ZN(n4685) );
  AOI22_X1 U3828 ( .A1(n2031), .A2(n2536), .B1(n1602), .B2(n3302), .ZN(n3713)
         );
  INV_X1 U3829 ( .A(n3716), .ZN(n4686) );
  AOI22_X1 U3830 ( .A1(n579), .A2(N1229), .B1(n1599), .B2(n3465), .ZN(n3716)
         );
  INV_X1 U3831 ( .A(n3717), .ZN(n4687) );
  AOI22_X1 U3832 ( .A1(n2035), .A2(N1228), .B1(n3292), .B2(n3464), .ZN(n3717)
         );
  OAI22_X1 U3833 ( .A1(n12401), .A2(n1798), .B1(n1614), .B2(n3719), .ZN(n4688)
         );
  INV_X1 U3834 ( .A(n2576), .ZN(n3719) );
  INV_X1 U3835 ( .A(n37201), .ZN(n4689) );
  AOI22_X1 U3836 ( .A1(n1719), .A2(n2914), .B1(n1603), .B2(n580), .ZN(n37201)
         );
  OAI22_X1 U3837 ( .A1(n1238), .A2(n577), .B1(n1611), .B2(n3722), .ZN(n46901)
         );
  INV_X1 U3838 ( .A(n3422), .ZN(n3722) );
  NOR2_X1 U3839 ( .A1(n3234), .A2(n2702), .ZN(N504) );
  NOR2_X1 U3840 ( .A1(n3235), .A2(n3007), .ZN(N503) );
  NOR2_X1 U3841 ( .A1(n1528), .A2(n1361), .ZN(N502) );
  NOR2_X1 U3842 ( .A1(n1528), .A2(n1537), .ZN(N501) );
  NOR2_X1 U3843 ( .A1(n3234), .A2(n2215), .ZN(N500) );
  NOR2_X1 U3844 ( .A1(n3235), .A2(n1136), .ZN(N499) );
  NOR2_X1 U3845 ( .A1(n3239), .A2(n1192), .ZN(N492) );
  NOR2_X1 U3846 ( .A1(n32401), .A2(n1465), .ZN(N491) );
  NOR2_X1 U3847 ( .A1(n1533), .A2(n1031), .ZN(N490) );
  NOR2_X1 U3848 ( .A1(n1533), .A2(n1535), .ZN(N489) );
  NOR2_X1 U3849 ( .A1(n3239), .A2(n2214), .ZN(N488) );
  NOR2_X1 U3850 ( .A1(n32401), .A2(n2694), .ZN(N487) );
  OAI22_X1 U3851 ( .A1(n2416), .A2(n2908), .B1(n3725), .B2(n1267), .ZN(N486)
         );
  OAI22_X1 U3852 ( .A1(n2413), .A2(n1018), .B1(n3728), .B2(n20201), .ZN(N485)
         );
  OAI22_X1 U3853 ( .A1(n2422), .A2(n2904), .B1(n37301), .B2(n1094), .ZN(N484)
         );
  OAI22_X1 U3854 ( .A1(n2419), .A2(n1016), .B1(n3732), .B2(n1094), .ZN(N483)
         );
  OAI22_X1 U3855 ( .A1(n2416), .A2(n29001), .B1(n3734), .B2(n2796), .ZN(N482)
         );
  OAI22_X1 U3856 ( .A1(n2414), .A2(n1014), .B1(n3736), .B2(n2021), .ZN(N481)
         );
  OAI22_X1 U3857 ( .A1(n2423), .A2(n1011), .B1(n3738), .B2(n3351), .ZN(N480)
         );
  OAI22_X1 U3858 ( .A1(n24201), .A2(n2898), .B1(n37401), .B2(n3351), .ZN(N479)
         );
  OAI22_X1 U3859 ( .A1(n2417), .A2(n1009), .B1(n3742), .B2(n1268), .ZN(N478)
         );
  OAI22_X1 U3860 ( .A1(n2413), .A2(n10101), .B1(n3744), .B2(n20201), .ZN(N477)
         );
  OAI22_X1 U3861 ( .A1(n2423), .A2(n1007), .B1(n3746), .B2(n1707), .ZN(N476)
         );
  OAI22_X1 U3862 ( .A1(n24201), .A2(n1008), .B1(n3748), .B2(n1708), .ZN(N475)
         );
  OAI22_X1 U3863 ( .A1(n2417), .A2(n2884), .B1(n37501), .B2(n2796), .ZN(N474)
         );
  OAI22_X1 U3864 ( .A1(n2414), .A2(n1006), .B1(n3752), .B2(n2021), .ZN(N473)
         );
  OAI22_X1 U3865 ( .A1(n2422), .A2(n1003), .B1(n3754), .B2(n2017), .ZN(N472)
         );
  OAI22_X1 U3866 ( .A1(n2419), .A2(n1004), .B1(n3756), .B2(n2017), .ZN(N471)
         );
  OAI21_X1 U3867 ( .B1(n1267), .B2(n3306), .A(n3298), .ZN(n3757) );
  NAND2_X1 U3868 ( .A1(n3229), .A2(n37601), .ZN(n3726) );
  OAI22_X1 U3869 ( .A1(n2279), .A2(n1001), .B1(n3763), .B2(n1261), .ZN(N470)
         );
  OAI22_X1 U3870 ( .A1(n2276), .A2(n1002), .B1(n3766), .B2(n2025), .ZN(N469)
         );
  OAI22_X1 U3871 ( .A1(n2285), .A2(n999), .B1(n3768), .B2(n1095), .ZN(N468) );
  OAI22_X1 U3872 ( .A1(n2282), .A2(n10001), .B1(n37701), .B2(n1095), .ZN(N467)
         );
  OAI22_X1 U3873 ( .A1(n2279), .A2(n997), .B1(n3772), .B2(n27901), .ZN(N466)
         );
  OAI22_X1 U3874 ( .A1(n2277), .A2(n998), .B1(n3774), .B2(n2026), .ZN(N465) );
  OAI22_X1 U3875 ( .A1(n2284), .A2(n995), .B1(n3776), .B2(n3352), .ZN(N464) );
  OAI22_X1 U3876 ( .A1(n2281), .A2(n996), .B1(n3778), .B2(n3352), .ZN(N463) );
  OAI22_X1 U3877 ( .A1(n22801), .A2(n993), .B1(n37801), .B2(n1262), .ZN(N462)
         );
  OAI22_X1 U3878 ( .A1(n2276), .A2(n994), .B1(n3782), .B2(n2025), .ZN(N461) );
  OAI22_X1 U3879 ( .A1(n2285), .A2(n991), .B1(n3784), .B2(n17101), .ZN(N460)
         );
  OAI22_X1 U3880 ( .A1(n2282), .A2(n992), .B1(n3786), .B2(n2022), .ZN(N459) );
  OAI22_X1 U3881 ( .A1(n22801), .A2(n989), .B1(n3788), .B2(n27901), .ZN(N458)
         );
  OAI22_X1 U3882 ( .A1(n2277), .A2(n990), .B1(n37901), .B2(n2026), .ZN(N457)
         );
  OAI22_X1 U3883 ( .A1(n2284), .A2(n987), .B1(n3792), .B2(n2022), .ZN(N456) );
  OAI22_X1 U3884 ( .A1(n2281), .A2(n988), .B1(n3794), .B2(n1711), .ZN(N455) );
  OAI22_X1 U3885 ( .A1(n2531), .A2(n1261), .B1(n2679), .B2(n1615), .ZN(n3795)
         );
  NAND2_X1 U3886 ( .A1(n3228), .A2(n583), .ZN(n3764) );
  OAI22_X1 U3887 ( .A1(n22401), .A2(n2844), .B1(n3798), .B2(n1271), .ZN(N454)
         );
  OAI22_X1 U3888 ( .A1(n2246), .A2(n2846), .B1(n3801), .B2(n20101), .ZN(N453)
         );
  OAI22_X1 U3889 ( .A1(n2244), .A2(n28401), .B1(n3803), .B2(n1092), .ZN(N452)
         );
  OAI22_X1 U3890 ( .A1(n2251), .A2(n2842), .B1(n3805), .B2(n1092), .ZN(N451)
         );
  OAI22_X1 U3891 ( .A1(n22401), .A2(n2836), .B1(n3807), .B2(n28001), .ZN(N450)
         );
  OAI22_X1 U3892 ( .A1(n2247), .A2(n2838), .B1(n3809), .B2(n2011), .ZN(N449)
         );
  OAI22_X1 U3893 ( .A1(n2243), .A2(n2832), .B1(n3811), .B2(n3349), .ZN(N448)
         );
  OAI22_X1 U3894 ( .A1(n22501), .A2(n2834), .B1(n3813), .B2(n3349), .ZN(N447)
         );
  OAI22_X1 U3895 ( .A1(n2241), .A2(n2828), .B1(n3815), .B2(n1272), .ZN(N446)
         );
  OAI22_X1 U3896 ( .A1(n2246), .A2(n28301), .B1(n3817), .B2(n20101), .ZN(N445)
         );
  OAI22_X1 U3897 ( .A1(n2243), .A2(n2824), .B1(n3819), .B2(n1701), .ZN(N444)
         );
  OAI22_X1 U3898 ( .A1(n22501), .A2(n2826), .B1(n3821), .B2(n2007), .ZN(N443)
         );
  OAI22_X1 U3899 ( .A1(n2241), .A2(n28201), .B1(n3823), .B2(n28001), .ZN(N442)
         );
  OAI22_X1 U3900 ( .A1(n2247), .A2(n2822), .B1(n3825), .B2(n2011), .ZN(N441)
         );
  OAI22_X1 U3901 ( .A1(n2244), .A2(n2816), .B1(n3827), .B2(n2007), .ZN(N440)
         );
  OAI22_X1 U3902 ( .A1(n2251), .A2(n2818), .B1(n3829), .B2(n1702), .ZN(N439)
         );
  OAI22_X1 U3903 ( .A1(n3303), .A2(n1271), .B1(n3831), .B2(n3296), .ZN(n38301)
         );
  NAND2_X1 U3904 ( .A1(n3227), .A2(n3832), .ZN(n3799) );
  OAI22_X1 U3905 ( .A1(n2381), .A2(n1181), .B1(n3834), .B2(n1265), .ZN(N438)
         );
  OAI22_X1 U3906 ( .A1(n2386), .A2(n1184), .B1(n3837), .B2(n2015), .ZN(N437)
         );
  OAI22_X1 U3907 ( .A1(n2384), .A2(n1175), .B1(n3839), .B2(n1093), .ZN(N436)
         );
  OAI22_X1 U3908 ( .A1(n2391), .A2(n1178), .B1(n3841), .B2(n1093), .ZN(N435)
         );
  OAI22_X1 U3909 ( .A1(n2381), .A2(n1169), .B1(n3843), .B2(n2794), .ZN(N434)
         );
  OAI22_X1 U3910 ( .A1(n2387), .A2(n1172), .B1(n3845), .B2(n2016), .ZN(N433)
         );
  OAI22_X1 U3911 ( .A1(n2383), .A2(n1163), .B1(n3847), .B2(n33501), .ZN(N432)
         );
  OAI22_X1 U3912 ( .A1(n23901), .A2(n1166), .B1(n3849), .B2(n33501), .ZN(N431)
         );
  OAI22_X1 U3913 ( .A1(n2382), .A2(n1157), .B1(n3851), .B2(n1266), .ZN(N430)
         );
  OAI22_X1 U3914 ( .A1(n2386), .A2(n11601), .B1(n3853), .B2(n2015), .ZN(N429)
         );
  OAI22_X1 U3915 ( .A1(n2383), .A2(n1151), .B1(n3855), .B2(n1704), .ZN(N428)
         );
  OAI22_X1 U3916 ( .A1(n23901), .A2(n1154), .B1(n3857), .B2(n1705), .ZN(N427)
         );
  OAI22_X1 U3917 ( .A1(n2382), .A2(n1145), .B1(n3859), .B2(n2794), .ZN(N426)
         );
  OAI22_X1 U3918 ( .A1(n2387), .A2(n1148), .B1(n3861), .B2(n2016), .ZN(N425)
         );
  OAI22_X1 U3919 ( .A1(n2384), .A2(n1139), .B1(n3863), .B2(n2012), .ZN(N424)
         );
  OAI22_X1 U3920 ( .A1(n2391), .A2(n1142), .B1(n3865), .B2(n2012), .ZN(N423)
         );
  OAI22_X1 U3921 ( .A1(n3867), .A2(n3297), .B1(n3304), .B2(n1265), .ZN(n3866)
         );
  NAND2_X1 U3922 ( .A1(n3229), .A2(n2681), .ZN(n3835) );
  OAI22_X1 U3923 ( .A1(n2373), .A2(n1468), .B1(n38701), .B2(n1259), .ZN(N422)
         );
  OAI22_X1 U3924 ( .A1(n23701), .A2(n1461), .B1(n3873), .B2(n2039), .ZN(N421)
         );
  OAI22_X1 U3925 ( .A1(n2379), .A2(n1454), .B1(n3875), .B2(n1097), .ZN(N420)
         );
  OAI22_X1 U3926 ( .A1(n2376), .A2(n1447), .B1(n3877), .B2(n1097), .ZN(N419)
         );
  OAI22_X1 U3927 ( .A1(n2373), .A2(n1442), .B1(n3879), .B2(n2788), .ZN(N418)
         );
  OAI22_X1 U3928 ( .A1(n2371), .A2(n1435), .B1(n3881), .B2(n20401), .ZN(N417)
         );
  OAI22_X1 U3929 ( .A1(n2378), .A2(n1428), .B1(n3883), .B2(n3358), .ZN(N416)
         );
  OAI22_X1 U3930 ( .A1(n2375), .A2(n1421), .B1(n3885), .B2(n3358), .ZN(N415)
         );
  OAI22_X1 U3931 ( .A1(n2374), .A2(n1416), .B1(n3887), .B2(n12601), .ZN(N414)
         );
  OAI22_X1 U3932 ( .A1(n23701), .A2(n1409), .B1(n3889), .B2(n2039), .ZN(N413)
         );
  OAI22_X1 U3933 ( .A1(n2379), .A2(n1404), .B1(n3891), .B2(n1722), .ZN(N412)
         );
  OAI22_X1 U3934 ( .A1(n2376), .A2(n1399), .B1(n3893), .B2(n2036), .ZN(N411)
         );
  OAI22_X1 U3935 ( .A1(n2374), .A2(n1394), .B1(n3895), .B2(n2788), .ZN(N410)
         );
  OAI22_X1 U3936 ( .A1(n2371), .A2(n1387), .B1(n3897), .B2(n20401), .ZN(N409)
         );
  OAI22_X1 U3937 ( .A1(n2378), .A2(n13801), .B1(n3899), .B2(n2036), .ZN(N408)
         );
  OAI22_X1 U3938 ( .A1(n2375), .A2(n1373), .B1(n3901), .B2(n1723), .ZN(N407)
         );
  OAI22_X1 U3939 ( .A1(n3305), .A2(n1259), .B1(n3242), .B2(n1614), .ZN(n3902)
         );
  OAI22_X1 U3940 ( .A1(n2395), .A2(n31501), .B1(n3906), .B2(n1257), .ZN(N406)
         );
  OAI22_X1 U3941 ( .A1(n2392), .A2(n3154), .B1(n3909), .B2(n2049), .ZN(N405)
         );
  OAI22_X1 U3942 ( .A1(n2401), .A2(n3142), .B1(n3911), .B2(n1099), .ZN(N404)
         );
  OAI22_X1 U3943 ( .A1(n2398), .A2(n3146), .B1(n3913), .B2(n1099), .ZN(N403)
         );
  OAI22_X1 U3944 ( .A1(n2395), .A2(n3134), .B1(n3915), .B2(n2783), .ZN(N402)
         );
  OAI22_X1 U3945 ( .A1(n2393), .A2(n3138), .B1(n3917), .B2(n20501), .ZN(N401)
         );
  OAI22_X1 U3946 ( .A1(n24001), .A2(n3126), .B1(n3919), .B2(n33601), .ZN(N400)
         );
  OAI22_X1 U3947 ( .A1(n2397), .A2(n31301), .B1(n3921), .B2(n33601), .ZN(N399)
         );
  OAI22_X1 U3948 ( .A1(n2396), .A2(n3118), .B1(n3923), .B2(n1258), .ZN(N398)
         );
  OAI22_X1 U3949 ( .A1(n2392), .A2(n3122), .B1(n3925), .B2(n2049), .ZN(N397)
         );
  OAI22_X1 U3950 ( .A1(n2401), .A2(n31101), .B1(n3927), .B2(n1728), .ZN(N396)
         );
  OAI22_X1 U3951 ( .A1(n2398), .A2(n3114), .B1(n3929), .B2(n2046), .ZN(N395)
         );
  OAI22_X1 U3952 ( .A1(n2396), .A2(n3102), .B1(n3931), .B2(n2783), .ZN(N394)
         );
  OAI22_X1 U3953 ( .A1(n2393), .A2(n3106), .B1(n3933), .B2(n20501), .ZN(N393)
         );
  OAI22_X1 U3954 ( .A1(n24001), .A2(n3094), .B1(n3935), .B2(n2046), .ZN(N392)
         );
  OAI22_X1 U3955 ( .A1(n2397), .A2(n3098), .B1(n3937), .B2(n1729), .ZN(N391)
         );
  OAI22_X1 U3956 ( .A1(n3939), .A2(n1615), .B1(n2523), .B2(n1257), .ZN(n3938)
         );
  OAI22_X1 U3957 ( .A1(n2358), .A2(n1457), .B1(n3941), .B2(n1255), .ZN(N390)
         );
  OAI22_X1 U3958 ( .A1(n2364), .A2(n14501), .B1(n3943), .B2(n2044), .ZN(N389)
         );
  OAI22_X1 U3959 ( .A1(n2362), .A2(n676), .B1(n3945), .B2(n1098), .ZN(N388) );
  OAI22_X1 U3960 ( .A1(n2369), .A2(n1438), .B1(n3946), .B2(n1098), .ZN(N387)
         );
  OAI22_X1 U3961 ( .A1(n2358), .A2(n1431), .B1(n3947), .B2(n2781), .ZN(N386)
         );
  OAI22_X1 U3962 ( .A1(n2365), .A2(n1424), .B1(n3948), .B2(n2045), .ZN(N385)
         );
  OAI22_X1 U3963 ( .A1(n2361), .A2(n2979), .B1(n39501), .B2(n3359), .ZN(N384)
         );
  OAI22_X1 U3964 ( .A1(n2368), .A2(n1412), .B1(n3951), .B2(n3359), .ZN(N383)
         );
  OAI22_X1 U3965 ( .A1(n2359), .A2(n2971), .B1(n3953), .B2(n1256), .ZN(N382)
         );
  OAI22_X1 U3966 ( .A1(n2364), .A2(n2967), .B1(n3955), .B2(n2044), .ZN(N381)
         );
  OAI22_X1 U3967 ( .A1(n2361), .A2(n2963), .B1(n3957), .B2(n1725), .ZN(N380)
         );
  OAI22_X1 U3968 ( .A1(n2368), .A2(n13901), .B1(n3958), .B2(n1726), .ZN(N379)
         );
  OAI22_X1 U3969 ( .A1(n2359), .A2(n1383), .B1(n3959), .B2(n2781), .ZN(N378)
         );
  OAI22_X1 U3970 ( .A1(n2365), .A2(n1376), .B1(n39601), .B2(n2045), .ZN(N377)
         );
  OAI22_X1 U3971 ( .A1(n2362), .A2(n663), .B1(n3962), .B2(n2041), .ZN(N376) );
  OAI22_X1 U3972 ( .A1(n2369), .A2(n1364), .B1(n3963), .B2(n2041), .ZN(N375)
         );
  OAI22_X1 U3973 ( .A1(n586), .A2(n1612), .B1(n25301), .B2(n1255), .ZN(n3964)
         );
  OAI22_X1 U3974 ( .A1(n1887), .A2(n3968), .B1(n3083), .B2(n1831), .ZN(N374)
         );
  OAI22_X1 U3975 ( .A1(n1884), .A2(n3971), .B1(n3087), .B2(n1828), .ZN(N373)
         );
  OAI22_X1 U3976 ( .A1(n33301), .A2(n3973), .B1(n3075), .B2(n3323), .ZN(N372)
         );
  OAI22_X1 U3977 ( .A1(n33301), .A2(n3975), .B1(n3079), .B2(n3323), .ZN(N371)
         );
  OAI22_X1 U3978 ( .A1(n1887), .A2(n3977), .B1(n3067), .B2(n1831), .ZN(N370)
         );
  OAI22_X1 U3979 ( .A1(n1885), .A2(n3979), .B1(n3071), .B2(n1829), .ZN(N369)
         );
  OAI22_X1 U3980 ( .A1(n1073), .A2(n3981), .B1(n3059), .B2(n1066), .ZN(N368)
         );
  OAI22_X1 U3981 ( .A1(n1073), .A2(n3983), .B1(n3063), .B2(n1066), .ZN(N367)
         );
  OAI22_X1 U3982 ( .A1(n1888), .A2(n3985), .B1(n3051), .B2(n1832), .ZN(N366)
         );
  OAI22_X1 U3983 ( .A1(n1884), .A2(n3987), .B1(n3055), .B2(n1828), .ZN(N365)
         );
  OAI22_X1 U3984 ( .A1(n1881), .A2(n3989), .B1(n3043), .B2(n16230), .ZN(N364)
         );
  OAI22_X1 U3985 ( .A1(n1881), .A2(n3991), .B1(n3047), .B2(n16240), .ZN(N363)
         );
  OAI22_X1 U3986 ( .A1(n1888), .A2(n3993), .B1(n3035), .B2(n1832), .ZN(N362)
         );
  OAI22_X1 U3987 ( .A1(n1885), .A2(n3995), .B1(n3039), .B2(n1829), .ZN(N361)
         );
  OAI22_X1 U3988 ( .A1(n1644), .A2(n3997), .B1(n3027), .B2(n1825), .ZN(N360)
         );
  OAI22_X1 U3989 ( .A1(n1645), .A2(n3999), .B1(n3031), .B2(n1825), .ZN(N359)
         );
  NAND2_X1 U3990 ( .A1(n3291), .A2(n4001), .ZN(n39701) );
  NOR2_X1 U3991 ( .A1(n1804), .A2(n9260), .ZN(n3759) );
  OAI22_X1 U3992 ( .A1(n3368), .A2(n1017), .B1(n1839), .B2(n4003), .ZN(N358)
         );
  INV_X1 U3993 ( .A(N1562), .ZN(n4003) );
  OAI22_X1 U3994 ( .A1(n1105), .A2(n29101), .B1(n1836), .B2(n4004), .ZN(N357)
         );
  INV_X1 U3995 ( .A(N1561), .ZN(n4004) );
  OAI22_X1 U3996 ( .A1(n12401), .A2(n1015), .B1(n3324), .B2(n4005), .ZN(N356)
         );
  INV_X1 U3997 ( .A(N1560), .ZN(n4005) );
  OAI22_X1 U3998 ( .A1(n2767), .A2(n2906), .B1(n16270), .B2(n4006), .ZN(N355)
         );
  INV_X1 U3999 ( .A(N1559), .ZN(n4006) );
  OAI22_X1 U4000 ( .A1(n2072), .A2(n1013), .B1(n1839), .B2(n4007), .ZN(N354)
         );
  INV_X1 U4001 ( .A(N1558), .ZN(n4007) );
  OAI22_X1 U4002 ( .A1(n2072), .A2(n29020), .B1(n1837), .B2(n4008), .ZN(N353)
         );
  INV_X1 U4003 ( .A(N1557), .ZN(n4008) );
  OAI22_X1 U4004 ( .A1(n2769), .A2(n2896), .B1(n1067), .B2(n4009), .ZN(N352)
         );
  INV_X1 U4005 ( .A(N1556), .ZN(n4009) );
  OAI22_X1 U4006 ( .A1(n1239), .A2(n1012), .B1(n1067), .B2(n40101), .ZN(N351)
         );
  INV_X1 U4007 ( .A(N1555), .ZN(n40101) );
  OAI22_X1 U4008 ( .A1(n1749), .A2(n2892), .B1(n18401), .B2(n4011), .ZN(N350)
         );
  INV_X1 U4009 ( .A(N1554), .ZN(n4011) );
  OAI22_X1 U4010 ( .A1(n17501), .A2(n2894), .B1(n1836), .B2(n4012), .ZN(N349)
         );
  INV_X1 U4011 ( .A(N1553), .ZN(n4012) );
  OAI22_X1 U4012 ( .A1(n2769), .A2(n2888), .B1(n1833), .B2(n4013), .ZN(N348)
         );
  INV_X1 U4013 ( .A(N1552), .ZN(n4013) );
  OAI22_X1 U4014 ( .A1(n2767), .A2(n28901), .B1(n3324), .B2(n4014), .ZN(N347)
         );
  INV_X1 U4015 ( .A(N1551), .ZN(n4014) );
  OAI22_X1 U4016 ( .A1(n1105), .A2(n1005), .B1(n18401), .B2(n4015), .ZN(N346)
         );
  INV_X1 U4017 ( .A(N1550), .ZN(n4015) );
  OAI22_X1 U4018 ( .A1(n3368), .A2(n2886), .B1(n1837), .B2(n4016), .ZN(N345)
         );
  INV_X1 U4019 ( .A(N1549), .ZN(n4016) );
  OAI22_X1 U4020 ( .A1(n1241), .A2(n28801), .B1(n16260), .B2(n4017), .ZN(N344)
         );
  INV_X1 U4021 ( .A(N1548), .ZN(n4017) );
  OAI22_X1 U4022 ( .A1(n1238), .A2(n2882), .B1(n1833), .B2(n4018), .ZN(N343)
         );
  INV_X1 U4023 ( .A(N1547), .ZN(n4018) );
  NAND2_X1 U4024 ( .A1(n3291), .A2(n4019), .ZN(n4002) );
  NAND3_X1 U4025 ( .A1(n1122), .A2(n2687), .A3(n40201), .ZN(n4019) );
  INV_X1 U4026 ( .A(n2786), .ZN(n3718) );
  OAI21_X1 U4027 ( .B1(n2876), .B2(n1815), .A(n4022), .ZN(N342) );
  NAND2_X1 U4028 ( .A1(N1596), .A2(n1251), .ZN(n4022) );
  OAI21_X1 U4029 ( .B1(n2878), .B2(n1812), .A(n4024), .ZN(N341) );
  NAND2_X1 U4030 ( .A1(N1595), .A2(n2054), .ZN(n4024) );
  OAI21_X1 U4031 ( .B1(n2872), .B2(n1809), .A(n4025), .ZN(N340) );
  NAND2_X1 U4032 ( .A1(N1594), .A2(n1731), .ZN(n4025) );
  OAI21_X1 U4033 ( .B1(n2874), .B2(n1806), .A(n4026), .ZN(N339) );
  NAND2_X1 U4034 ( .A1(N1593), .A2(n3361), .ZN(n4026) );
  OAI21_X1 U4035 ( .B1(n2868), .B2(n1816), .A(n4027), .ZN(N338) );
  NAND2_X1 U4036 ( .A1(N1592), .A2(n1252), .ZN(n4027) );
  OAI21_X1 U4037 ( .B1(n28701), .B2(n1813), .A(n4028), .ZN(N337) );
  NAND2_X1 U4038 ( .A1(N1591), .A2(n2055), .ZN(n4028) );
  OAI21_X1 U4039 ( .B1(n2864), .B2(n18101), .A(n4029), .ZN(N336) );
  NAND2_X1 U4040 ( .A1(N1590), .A2(n3361), .ZN(n4029) );
  OAI21_X1 U4041 ( .B1(n2866), .B2(n1807), .A(n40301), .ZN(N335) );
  NAND2_X1 U4042 ( .A1(N1589), .A2(n11001), .ZN(n40301) );
  OAI21_X1 U4043 ( .B1(n28601), .B2(n1815), .A(n4031), .ZN(N334) );
  NAND2_X1 U4044 ( .A1(N1588), .A2(n2777), .ZN(n4031) );
  OAI21_X1 U4045 ( .B1(n2862), .B2(n1812), .A(n4032), .ZN(N333) );
  NAND2_X1 U4046 ( .A1(N1587), .A2(n2054), .ZN(n4032) );
  OAI21_X1 U4047 ( .B1(n2856), .B2(n18101), .A(n4033), .ZN(N332) );
  NAND2_X1 U4048 ( .A1(N1586), .A2(n11001), .ZN(n4033) );
  OAI21_X1 U4049 ( .B1(n2858), .B2(n1807), .A(n4034), .ZN(N331) );
  NAND2_X1 U4050 ( .A1(N1585), .A2(n1732), .ZN(n4034) );
  OAI21_X1 U4051 ( .B1(n2852), .B2(n1816), .A(n4035), .ZN(N330) );
  NAND2_X1 U4052 ( .A1(N1584), .A2(n2777), .ZN(n4035) );
  OAI21_X1 U4053 ( .B1(n2854), .B2(n1813), .A(n4036), .ZN(N329) );
  NAND2_X1 U4054 ( .A1(N1583), .A2(n2055), .ZN(n4036) );
  OAI21_X1 U4055 ( .B1(n2848), .B2(n1809), .A(n4037), .ZN(N328) );
  NAND2_X1 U4056 ( .A1(N1582), .A2(n2051), .ZN(n4037) );
  OAI21_X1 U4057 ( .B1(n28501), .B2(n1806), .A(n4038), .ZN(N327) );
  NAND2_X1 U4058 ( .A1(N1581), .A2(n2051), .ZN(n4038) );
  NAND2_X1 U4059 ( .A1(n3357), .A2(n4039), .ZN(n4021) );
  NAND3_X1 U4060 ( .A1(n3722), .A2(n1799), .A3(n40401), .ZN(n4039) );
  OAI22_X1 U4061 ( .A1(n1951), .A2(n4042), .B1(n2843), .B2(n1247), .ZN(N326)
         );
  INV_X1 U4062 ( .A(N1638), .ZN(n4042) );
  OAI22_X1 U4063 ( .A1(n1948), .A2(n4044), .B1(n2845), .B2(n2064), .ZN(N325)
         );
  INV_X1 U4064 ( .A(N1637), .ZN(n4044) );
  OAI22_X1 U4065 ( .A1(n1668), .A2(n4045), .B1(n2839), .B2(n1102), .ZN(N324)
         );
  INV_X1 U4066 ( .A(N1636), .ZN(n4045) );
  OAI22_X1 U4067 ( .A1(n1945), .A2(n4046), .B1(n2841), .B2(n1102), .ZN(N323)
         );
  INV_X1 U4068 ( .A(N1635), .ZN(n4046) );
  OAI22_X1 U4069 ( .A1(n1951), .A2(n4047), .B1(n2835), .B2(n2773), .ZN(N322)
         );
  INV_X1 U4070 ( .A(N1634), .ZN(n4047) );
  OAI22_X1 U4071 ( .A1(n1949), .A2(n4048), .B1(n2837), .B2(n2065), .ZN(N321)
         );
  INV_X1 U4072 ( .A(N1633), .ZN(n4048) );
  OAI22_X1 U4073 ( .A1(n1945), .A2(n4049), .B1(n2831), .B2(n3363), .ZN(N320)
         );
  INV_X1 U4074 ( .A(N1632), .ZN(n4049) );
  OAI22_X1 U4075 ( .A1(n3338), .A2(n40501), .B1(n2833), .B2(n3363), .ZN(N319)
         );
  INV_X1 U4076 ( .A(N1631), .ZN(n40501) );
  OAI22_X1 U4077 ( .A1(n1952), .A2(n4051), .B1(n2827), .B2(n1248), .ZN(N318)
         );
  INV_X1 U4078 ( .A(N1630), .ZN(n4051) );
  OAI22_X1 U4079 ( .A1(n1948), .A2(n4052), .B1(n2829), .B2(n2064), .ZN(N317)
         );
  INV_X1 U4080 ( .A(N1629), .ZN(n4052) );
  OAI22_X1 U4081 ( .A1(n3338), .A2(n4053), .B1(n2823), .B2(n1737), .ZN(N316)
         );
  INV_X1 U4082 ( .A(N1628), .ZN(n4053) );
  OAI22_X1 U4083 ( .A1(n1669), .A2(n4054), .B1(n2825), .B2(n2061), .ZN(N315)
         );
  INV_X1 U4084 ( .A(N1627), .ZN(n4054) );
  OAI22_X1 U4085 ( .A1(n1952), .A2(n4055), .B1(n2819), .B2(n2773), .ZN(N314)
         );
  INV_X1 U4086 ( .A(N1626), .ZN(n4055) );
  OAI22_X1 U4087 ( .A1(n1949), .A2(n4056), .B1(n2821), .B2(n2065), .ZN(N313)
         );
  INV_X1 U4088 ( .A(N1625), .ZN(n4056) );
  OAI22_X1 U4089 ( .A1(n1081), .A2(n4057), .B1(n2815), .B2(n2061), .ZN(N312)
         );
  INV_X1 U4090 ( .A(N1624), .ZN(n4057) );
  OAI22_X1 U4091 ( .A1(n1081), .A2(n4058), .B1(n2817), .B2(n1738), .ZN(N311)
         );
  INV_X1 U4092 ( .A(N1623), .ZN(n4058) );
  INV_X1 U4093 ( .A(n4059), .ZN(n40201) );
  OAI22_X1 U4094 ( .A1(n40601), .A2(n2163), .B1(n1182), .B2(n2183), .ZN(N310)
         );
  INV_X1 U4095 ( .A(n4063), .ZN(n40601) );
  OAI22_X1 U4096 ( .A1(n4064), .A2(n2166), .B1(n1185), .B2(n2186), .ZN(N309)
         );
  INV_X1 U4097 ( .A(n4065), .ZN(n4064) );
  OAI22_X1 U4098 ( .A1(n4066), .A2(n2168), .B1(n1176), .B2(n2189), .ZN(N308)
         );
  INV_X1 U4099 ( .A(n4067), .ZN(n4066) );
  OAI22_X1 U4100 ( .A1(n4068), .A2(n2163), .B1(n1179), .B2(n2183), .ZN(N307)
         );
  INV_X1 U4101 ( .A(n4069), .ZN(n4068) );
  OAI22_X1 U4102 ( .A1(n40701), .A2(n2166), .B1(n11701), .B2(n2186), .ZN(N306)
         );
  INV_X1 U4103 ( .A(n4071), .ZN(n40701) );
  OAI22_X1 U4104 ( .A1(n4072), .A2(n2168), .B1(n1173), .B2(n2189), .ZN(N305)
         );
  INV_X1 U4105 ( .A(n4073), .ZN(n4072) );
  OAI22_X1 U4106 ( .A1(n4074), .A2(n2164), .B1(n1164), .B2(n2184), .ZN(N304)
         );
  INV_X1 U4107 ( .A(n4075), .ZN(n4074) );
  OAI22_X1 U4108 ( .A1(n4076), .A2(n2167), .B1(n1167), .B2(n2187), .ZN(N303)
         );
  INV_X1 U4109 ( .A(n4077), .ZN(n4076) );
  OAI22_X1 U4110 ( .A1(n4078), .A2(n2169), .B1(n1158), .B2(n21901), .ZN(N302)
         );
  INV_X1 U4111 ( .A(n4079), .ZN(n4078) );
  OAI22_X1 U4112 ( .A1(n40801), .A2(n2164), .B1(n1161), .B2(n2184), .ZN(N301)
         );
  INV_X1 U4113 ( .A(n4081), .ZN(n40801) );
  OAI22_X1 U4114 ( .A1(n4082), .A2(n2167), .B1(n1152), .B2(n2187), .ZN(N300)
         );
  INV_X1 U4115 ( .A(n4083), .ZN(n4082) );
  OAI22_X1 U4116 ( .A1(n4084), .A2(n2169), .B1(n1155), .B2(n21901), .ZN(N299)
         );
  INV_X1 U4117 ( .A(n4085), .ZN(n4084) );
  OAI22_X1 U4118 ( .A1(n4086), .A2(n2161), .B1(n1146), .B2(n21801), .ZN(N298)
         );
  INV_X1 U4119 ( .A(n4087), .ZN(n4086) );
  OAI22_X1 U4120 ( .A1(n4088), .A2(n2161), .B1(n1149), .B2(n21801), .ZN(N297)
         );
  INV_X1 U4121 ( .A(n4089), .ZN(n4088) );
  OAI22_X1 U4122 ( .A1(n40901), .A2(n2162), .B1(n11401), .B2(n2181), .ZN(N296)
         );
  INV_X1 U4123 ( .A(n4091), .ZN(n40901) );
  OAI22_X1 U4124 ( .A1(n4092), .A2(n2162), .B1(n1143), .B2(n2181), .ZN(N295)
         );
  INV_X1 U4125 ( .A(n557), .ZN(n3721) );
  NAND2_X1 U4126 ( .A1(n2692), .A2(n4095), .ZN(n4059) );
  INV_X1 U4127 ( .A(n4096), .ZN(n4092) );
  OAI221_X1 U4128 ( .B1(n1052), .B2(n1249), .C1(n3084), .C2(n1895), .A(n4099), 
        .ZN(N294) );
  AOI22_X1 U4129 ( .A1(n1072), .A2(n46400), .B1(n1065), .B2(n56), .ZN(n4099)
         );
  OAI221_X1 U4130 ( .B1(n1051), .B2(n2069), .C1(n3088), .C2(n1892), .A(n4102), 
        .ZN(N293) );
  AOI22_X1 U4131 ( .A1(n18801), .A2(n46900), .B1(n1824), .B2(n58), .ZN(n4102)
         );
  OAI221_X1 U4132 ( .B1(n10501), .B2(n1103), .C1(n3076), .C2(n1074), .A(n4103), 
        .ZN(N292) );
  AOI22_X1 U4133 ( .A1(n1876), .A2(n4740), .B1(n18201), .B2(n60), .ZN(n4103)
         );
  OAI221_X1 U4134 ( .B1(n1049), .B2(n1103), .C1(n30801), .C2(n1648), .A(n4104), 
        .ZN(N291) );
  AOI22_X1 U4135 ( .A1(n1072), .A2(n4790), .B1(n3322), .B2(n62), .ZN(n4104) );
  OAI221_X1 U4136 ( .B1(n1048), .B2(n2775), .C1(n3068), .C2(n1895), .A(n4105), 
        .ZN(N290) );
  AOI22_X1 U4137 ( .A1(n3329), .A2(n4840), .B1(n3322), .B2(n64), .ZN(n4105) );
  OAI221_X1 U4138 ( .B1(n1047), .B2(n20701), .C1(n3072), .C2(n1893), .A(n4106), 
        .ZN(N289) );
  AOI22_X1 U4139 ( .A1(n1879), .A2(n4890), .B1(n1823), .B2(n66), .ZN(n4106) );
  OAI221_X1 U4140 ( .B1(n1046), .B2(n3364), .C1(n30601), .C2(n3331), .A(n4107), 
        .ZN(N288) );
  AOI22_X1 U4141 ( .A1(n1877), .A2(n494), .B1(n1821), .B2(n68), .ZN(n4107) );
  OAI221_X1 U4142 ( .B1(n1045), .B2(n3364), .C1(n3064), .C2(n1074), .A(n4108), 
        .ZN(N287) );
  AOI22_X1 U4143 ( .A1(n3329), .A2(n4990), .B1(n1817), .B2(n70), .ZN(n4108) );
  OAI221_X1 U4144 ( .B1(n1043), .B2(n12501), .C1(n3052), .C2(n1896), .A(n4109), 
        .ZN(N286) );
  AOI22_X1 U4145 ( .A1(n1873), .A2(n5040), .B1(n1817), .B2(n72), .ZN(n4109) );
  OAI221_X1 U4146 ( .B1(n1042), .B2(n2069), .C1(n3056), .C2(n1892), .A(n41101), 
        .ZN(N285) );
  AOI22_X1 U4147 ( .A1(n18801), .A2(n509), .B1(n1824), .B2(n74), .ZN(n41101)
         );
  OAI221_X1 U4148 ( .B1(n10401), .B2(n17401), .C1(n3044), .C2(n1889), .A(n4111), .ZN(N284) );
  AOI22_X1 U4149 ( .A1(n1876), .A2(n514), .B1(n18201), .B2(n76), .ZN(n4111) );
  OAI221_X1 U4150 ( .B1(n1038), .B2(n2066), .C1(n3048), .C2(n1889), .A(n4112), 
        .ZN(N283) );
  AOI22_X1 U4151 ( .A1(n1873), .A2(n519), .B1(n16201), .B2(n78), .ZN(n4112) );
  OAI221_X1 U4152 ( .B1(n1036), .B2(n2775), .C1(n3036), .C2(n1896), .A(n4113), 
        .ZN(N282) );
  AOI22_X1 U4153 ( .A1(n1641), .A2(n524), .B1(n1621), .B2(n80), .ZN(n4113) );
  OAI221_X1 U4154 ( .B1(n1035), .B2(n20701), .C1(n30401), .C2(n1893), .A(n4114), .ZN(N281) );
  AOI22_X1 U4155 ( .A1(n1879), .A2(n529), .B1(n1823), .B2(n82), .ZN(n4114) );
  OAI221_X1 U4156 ( .B1(n1034), .B2(n2066), .C1(n3028), .C2(n1647), .A(n4115), 
        .ZN(N280) );
  AOI22_X1 U4157 ( .A1(n1877), .A2(n534), .B1(n1821), .B2(n84), .ZN(n4115) );
  OAI221_X1 U4158 ( .B1(n1033), .B2(n1741), .C1(n3032), .C2(n3331), .A(n4116), 
        .ZN(N279) );
  AOI22_X1 U4159 ( .A1(n1642), .A2(n539), .B1(n1065), .B2(n86), .ZN(n4116) );
  AND2_X1 U4160 ( .A1(n4117), .A2(n2078), .ZN(n4101) );
  NOR2_X1 U4161 ( .A1(n1611), .A2(n41201), .ZN(n4117) );
  AOI21_X1 U4162 ( .B1(N1539), .B2(n1797), .A(n4121), .ZN(n41201) );
  OAI222_X1 U4163 ( .A1(n3148), .A2(n1959), .B1(n1458), .B2(n1935), .C1(n3085), 
        .C2(n1927), .ZN(N278) );
  OAI222_X1 U4164 ( .A1(n3152), .A2(n1956), .B1(n1451), .B2(n1932), .C1(n3089), 
        .C2(n1924), .ZN(N277) );
  OAI222_X1 U4165 ( .A1(n31401), .A2(n3339), .B1(n676), .B2(n3336), .C1(n3077), 
        .C2(n1078), .ZN(N276) );
  OAI222_X1 U4166 ( .A1(n3144), .A2(n3339), .B1(n1439), .B2(n3336), .C1(n3081), 
        .C2(n1078), .ZN(N275) );
  OAI222_X1 U4167 ( .A1(n3132), .A2(n1959), .B1(n1432), .B2(n1935), .C1(n3069), 
        .C2(n1928), .ZN(N274) );
  OAI222_X1 U4168 ( .A1(n3136), .A2(n1957), .B1(n1425), .B2(n1933), .C1(n3073), 
        .C2(n1925), .ZN(N273) );
  OAI222_X1 U4169 ( .A1(n3124), .A2(n1082), .B1(n2979), .B2(n1079), .C1(n3061), 
        .C2(n3335), .ZN(N272) );
  OAI222_X1 U4170 ( .A1(n3128), .A2(n1082), .B1(n1413), .B2(n1079), .C1(n3065), 
        .C2(n3335), .ZN(N271) );
  OAI222_X1 U4171 ( .A1(n3116), .A2(n19601), .B1(n2971), .B2(n1936), .C1(n3053), .C2(n1927), .ZN(N270) );
  OAI222_X1 U4172 ( .A1(n31201), .A2(n1956), .B1(n2967), .B2(n1932), .C1(n3057), .C2(n1924), .ZN(N269) );
  OAI222_X1 U4173 ( .A1(n3108), .A2(n1671), .B1(n2963), .B2(n1662), .C1(n3045), 
        .C2(n1659), .ZN(N268) );
  OAI222_X1 U4174 ( .A1(n3112), .A2(n1672), .B1(n1391), .B2(n1663), .C1(n3049), 
        .C2(n16601), .ZN(N267) );
  OAI222_X1 U4175 ( .A1(n31001), .A2(n19601), .B1(n1384), .B2(n1936), .C1(
        n3037), .C2(n1928), .ZN(N266) );
  OAI222_X1 U4176 ( .A1(n3104), .A2(n1957), .B1(n1377), .B2(n1933), .C1(n3041), 
        .C2(n1925), .ZN(N265) );
  OAI222_X1 U4177 ( .A1(n3092), .A2(n1953), .B1(n663), .B2(n1929), .C1(n3029), 
        .C2(n1921), .ZN(N264) );
  OAI222_X1 U4178 ( .A1(n3096), .A2(n1953), .B1(n1365), .B2(n1929), .C1(n3033), 
        .C2(n1921), .ZN(N263) );
  NAND3_X1 U4179 ( .A1(n1599), .A2(n581), .A3(n3319), .ZN(n4124) );
  OAI21_X1 U4180 ( .B1(n2686), .B2(n809), .A(n2693), .ZN(n4121) );
  OAI22_X1 U4181 ( .A1(n3086), .A2(n1943), .B1(n3003), .B2(n1919), .ZN(N262)
         );
  OAI22_X1 U4182 ( .A1(n30901), .A2(n19401), .B1(n2999), .B2(n1916), .ZN(N261)
         );
  OAI22_X1 U4183 ( .A1(n3078), .A2(n3337), .B1(n2995), .B2(n3334), .ZN(N260)
         );
  OAI22_X1 U4184 ( .A1(n3082), .A2(n3337), .B1(n2991), .B2(n3334), .ZN(N259)
         );
  OAI22_X1 U4185 ( .A1(n30701), .A2(n1943), .B1(n2987), .B2(n1919), .ZN(N258)
         );
  OAI22_X1 U4186 ( .A1(n3074), .A2(n1941), .B1(n2983), .B2(n1917), .ZN(N257)
         );
  OAI22_X1 U4187 ( .A1(n3062), .A2(n10801), .B1(n29801), .B2(n1077), .ZN(N256)
         );
  OAI22_X1 U4188 ( .A1(n3066), .A2(n10801), .B1(n2975), .B2(n1077), .ZN(N255)
         );
  OAI22_X1 U4189 ( .A1(n3054), .A2(n1944), .B1(n2972), .B2(n19201), .ZN(N254)
         );
  OAI22_X1 U4190 ( .A1(n3058), .A2(n19401), .B1(n2968), .B2(n1916), .ZN(N253)
         );
  OAI22_X1 U4191 ( .A1(n3046), .A2(n1937), .B1(n2964), .B2(n1656), .ZN(N252)
         );
  OAI22_X1 U4192 ( .A1(n30501), .A2(n1937), .B1(n2959), .B2(n1657), .ZN(N251)
         );
  OAI22_X1 U4193 ( .A1(n3038), .A2(n1944), .B1(n2955), .B2(n19201), .ZN(N250)
         );
  OAI22_X1 U4194 ( .A1(n3042), .A2(n1941), .B1(n2951), .B2(n1917), .ZN(N249)
         );
  OAI22_X1 U4195 ( .A1(n30301), .A2(n1665), .B1(n2947), .B2(n1913), .ZN(N248)
         );
  OAI22_X1 U4196 ( .A1(n3034), .A2(n1666), .B1(n2944), .B2(n1913), .ZN(N247)
         );
  INV_X1 U4197 ( .A(n40401), .ZN(n4094) );
  NOR2_X1 U4198 ( .A1(n4128), .A2(n33001), .ZN(n40401) );
  INV_X1 U4199 ( .A(n1249), .ZN(n4125) );
  INV_X1 U4200 ( .A(n2693), .ZN(n41301) );
  NOR3_X1 U4201 ( .A1(n1122), .A2(n2686), .A3(n809), .ZN(n4129) );
  INV_X1 U4202 ( .A(N1539), .ZN(n4095) );
  OAI211_X1 U4203 ( .C1(n3085), .C2(n1083), .A(n4132), .B(n4133), .ZN(N246) );
  AOI222_X1 U4204 ( .A1(n16360), .A2(n54), .B1(n1865), .B2(n31700), .C1(n16300), .C2(n22200), .ZN(n4133) );
  AOI22_X1 U4205 ( .A1(n1075), .A2(n27000), .B1(n2234), .B2(n4063), .ZN(n4132)
         );
  OAI221_X1 U4206 ( .B1(n1106), .B2(n3004), .C1(n1107), .C2(n3147), .A(n4141), 
        .ZN(n4063) );
  AOI22_X1 U4207 ( .A1(n1245), .A2(n38300), .B1(n15970), .B2(n12280), .ZN(
        n4141) );
  OAI211_X1 U4208 ( .C1(n3089), .C2(n1965), .A(n4143), .B(n4144), .ZN(N245) );
  AOI222_X1 U4209 ( .A1(n1863), .A2(n53), .B1(n1871), .B2(n32100), .C1(n1847), 
        .C2(n22500), .ZN(n4144) );
  AOI22_X1 U4210 ( .A1(n1903), .A2(n27300), .B1(n2232), .B2(n4065), .ZN(n4143)
         );
  OAI221_X1 U4211 ( .B1(n2765), .B2(n30001), .C1(n2755), .C2(n3151), .A(n4145), 
        .ZN(n4065) );
  AOI22_X1 U4212 ( .A1(n38800), .A2(n2771), .B1(n16390), .B2(n12260), .ZN(
        n4145) );
  OAI211_X1 U4213 ( .C1(n3077), .C2(n1964), .A(n4146), .B(n4147), .ZN(N244) );
  AOI222_X1 U4214 ( .A1(n18601), .A2(n52), .B1(n1868), .B2(n32500), .C1(n1844), 
        .C2(n22800), .ZN(n4147) );
  AOI22_X1 U4215 ( .A1(n19001), .A2(n27600), .B1(n2229), .B2(n4067), .ZN(n4146) );
  OAI221_X1 U4216 ( .B1(n2763), .B2(n2996), .C1(n2761), .C2(n3139), .A(n4148), 
        .ZN(n4067) );
  AOI22_X1 U4217 ( .A1(n39300), .A2(n2071), .B1(n16700), .B2(n2079), .ZN(n4148) );
  OAI211_X1 U4218 ( .C1(n3081), .C2(n33401), .A(n4149), .B(n41501), .ZN(N243)
         );
  AOI222_X1 U4219 ( .A1(n3327), .A2(n51), .B1(n1071), .B2(n32900), .C1(n1068), 
        .C2(n23100), .ZN(n41501) );
  AOI22_X1 U4220 ( .A1(n1897), .A2(n27900), .B1(n2238), .B2(n4069), .ZN(n4149)
         );
  OAI221_X1 U4221 ( .B1(n33701), .B2(n2992), .C1(n3372), .C2(n3143), .A(n4151), 
        .ZN(n4069) );
  AOI22_X1 U4222 ( .A1(n39800), .A2(n2071), .B1(n17100), .B2(n12280), .ZN(
        n4151) );
  OAI211_X1 U4223 ( .C1(n3069), .C2(n1961), .A(n4152), .B(n4153), .ZN(N242) );
  AOI222_X1 U4224 ( .A1(n3327), .A2(n50), .B1(n1071), .B2(n33300), .C1(n1068), 
        .C2(n23400), .ZN(n4153) );
  AOI22_X1 U4225 ( .A1(n1897), .A2(n28200), .B1(n2234), .B2(n4071), .ZN(n4152)
         );
  OAI221_X1 U4226 ( .B1(n3369), .B2(n2988), .C1(n3371), .C2(n3131), .A(n4154), 
        .ZN(n4071) );
  AOI22_X1 U4227 ( .A1(n40300), .A2(n556), .B1(n17500), .B2(n2753), .ZN(n4154)
         );
  OAI211_X1 U4228 ( .C1(n3073), .C2(n1966), .A(n4155), .B(n4156), .ZN(N241) );
  AOI222_X1 U4229 ( .A1(n1863), .A2(n49), .B1(n1872), .B2(n33700), .C1(n1848), 
        .C2(n23700), .ZN(n4156) );
  AOI22_X1 U4230 ( .A1(n1903), .A2(n28500), .B1(n2232), .B2(n4073), .ZN(n4155)
         );
  OAI221_X1 U4231 ( .B1(n1237), .B2(n2984), .C1(n1231), .C2(n3135), .A(n4157), 
        .ZN(n4073) );
  AOI22_X1 U4232 ( .A1(n40800), .A2(n1243), .B1(n17900), .B2(n2752), .ZN(n4157) );
  OAI211_X1 U4233 ( .C1(n3061), .C2(n1963), .A(n4158), .B(n4159), .ZN(N240) );
  AOI222_X1 U4234 ( .A1(n1861), .A2(n48), .B1(n1869), .B2(n34100), .C1(n1845), 
        .C2(n24000), .ZN(n4159) );
  AOI22_X1 U4235 ( .A1(n1901), .A2(n28800), .B1(n22301), .B2(n4075), .ZN(n4158) );
  OAI221_X1 U4236 ( .B1(n1235), .B2(n1044), .C1(n1233), .C2(n3123), .A(n41601), 
        .ZN(n4075) );
  AOI22_X1 U4237 ( .A1(n41300), .A2(n1104), .B1(n18300), .B2(n1108), .ZN(
        n41601) );
  OAI211_X1 U4238 ( .C1(n3065), .C2(n1083), .A(n4161), .B(n4162), .ZN(N239) );
  AOI222_X1 U4239 ( .A1(n10701), .A2(n47), .B1(n3328), .B2(n34500), .C1(n3325), 
        .C2(n24300), .ZN(n4162) );
  AOI22_X1 U4240 ( .A1(n3332), .A2(n29100), .B1(n2237), .B2(n4077), .ZN(n4161)
         );
  OAI221_X1 U4241 ( .B1(n33701), .B2(n2976), .C1(n3372), .C2(n3127), .A(n4163), 
        .ZN(n4077) );
  AOI22_X1 U4242 ( .A1(n41800), .A2(n3366), .B1(n18700), .B2(n2076), .ZN(n4163) );
  OAI211_X1 U4243 ( .C1(n3053), .C2(n33401), .A(n4164), .B(n4165), .ZN(N238)
         );
  AOI222_X1 U4244 ( .A1(n10701), .A2(n46), .B1(n3328), .B2(n34900), .C1(n3325), 
        .C2(n24600), .ZN(n4165) );
  AOI22_X1 U4245 ( .A1(n3332), .A2(n29400), .B1(n2235), .B2(n4079), .ZN(n4164)
         );
  OAI221_X1 U4246 ( .B1(n1753), .B2(n1041), .C1(n2756), .C2(n3115), .A(n4166), 
        .ZN(n4079) );
  AOI22_X1 U4247 ( .A1(n42300), .A2(n1246), .B1(n19100), .B2(n2076), .ZN(n4166) );
  OAI211_X1 U4248 ( .C1(n3057), .C2(n1965), .A(n4167), .B(n4168), .ZN(N237) );
  AOI222_X1 U4249 ( .A1(n1864), .A2(n45), .B1(n1871), .B2(n35300), .C1(n1847), 
        .C2(n24900), .ZN(n4168) );
  AOI22_X1 U4250 ( .A1(n1904), .A2(n29700), .B1(n2233), .B2(n4081), .ZN(n4167)
         );
  OAI221_X1 U4251 ( .B1(n2765), .B2(n1039), .C1(n2755), .C2(n3119), .A(n4169), 
        .ZN(n4081) );
  AOI22_X1 U4252 ( .A1(n42800), .A2(n2771), .B1(n19500), .B2(n1227), .ZN(n4169) );
  OAI211_X1 U4253 ( .C1(n3045), .C2(n1963), .A(n41701), .B(n4171), .ZN(N236)
         );
  AOI222_X1 U4254 ( .A1(n18601), .A2(n44), .B1(n1868), .B2(n35700), .C1(n1844), 
        .C2(n25200), .ZN(n4171) );
  AOI22_X1 U4255 ( .A1(n19001), .A2(n30000), .B1(n2229), .B2(n4083), .ZN(
        n41701) );
  OAI221_X1 U4256 ( .B1(n2763), .B2(n1037), .C1(n2761), .C2(n3107), .A(n4172), 
        .ZN(n4083) );
  AOI22_X1 U4257 ( .A1(n43300), .A2(n3365), .B1(n19900), .B2(n12290), .ZN(
        n4172) );
  OAI211_X1 U4258 ( .C1(n3049), .C2(n1961), .A(n4173), .B(n4174), .ZN(N235) );
  AOI222_X1 U4259 ( .A1(n16350), .A2(n43), .B1(n1865), .B2(n36100), .C1(n16290), .C2(n25500), .ZN(n4174) );
  AOI22_X1 U4260 ( .A1(n1075), .A2(n30300), .B1(n2238), .B2(n4085), .ZN(n4173)
         );
  OAI221_X1 U4261 ( .B1(n1754), .B2(n29601), .C1(n2756), .C2(n3111), .A(n4175), 
        .ZN(n4085) );
  AOI22_X1 U4262 ( .A1(n43800), .A2(n3366), .B1(n20300), .B2(n2078), .ZN(n4175) );
  OAI211_X1 U4263 ( .C1(n3037), .C2(n1675), .A(n4176), .B(n4177), .ZN(N234) );
  AOI222_X1 U4264 ( .A1(n1857), .A2(n42), .B1(n16391), .B2(n36500), .C1(n1841), 
        .C2(n25800), .ZN(n4177) );
  AOI22_X1 U4265 ( .A1(n1651), .A2(n30600), .B1(n2235), .B2(n4087), .ZN(n4176)
         );
  OAI221_X1 U4266 ( .B1(n2758), .B2(n2956), .C1(n1757), .C2(n3099), .A(n4178), 
        .ZN(n4087) );
  AOI22_X1 U4267 ( .A1(n44300), .A2(n556), .B1(n20700), .B2(n2079), .ZN(n4178)
         );
  OAI211_X1 U4268 ( .C1(n3041), .C2(n1966), .A(n4179), .B(n41801), .ZN(N233)
         );
  AOI222_X1 U4269 ( .A1(n1864), .A2(n41), .B1(n1872), .B2(n36900), .C1(n1848), 
        .C2(n26100), .ZN(n41801) );
  AOI22_X1 U4270 ( .A1(n1904), .A2(n30900), .B1(n2233), .B2(n4089), .ZN(n4179)
         );
  OAI221_X1 U4271 ( .B1(n1236), .B2(n2952), .C1(n12301), .C2(n3103), .A(n4181), 
        .ZN(n4089) );
  AOI22_X1 U4272 ( .A1(n44800), .A2(n1242), .B1(n21100), .B2(n2752), .ZN(n4181) );
  OAI211_X1 U4273 ( .C1(n3029), .C2(n1964), .A(n4182), .B(n4183), .ZN(N232) );
  AOI222_X1 U4274 ( .A1(n1861), .A2(n40), .B1(n1869), .B2(n37300), .C1(n1845), 
        .C2(n26400), .ZN(n4183) );
  AOI22_X1 U4275 ( .A1(n1901), .A2(n31200), .B1(n22301), .B2(n4091), .ZN(n4182) );
  OAI221_X1 U4276 ( .B1(n1234), .B2(n2948), .C1(n1232), .C2(n3091), .A(n4184), 
        .ZN(n4091) );
  AOI22_X1 U4277 ( .A1(n45300), .A2(n1745), .B1(n21500), .B2(n2075), .ZN(n4184) );
  OAI211_X1 U4278 ( .C1(n3033), .C2(n1674), .A(n4185), .B(n4186), .ZN(N231) );
  AOI222_X1 U4279 ( .A1(n1857), .A2(n39), .B1(n16380), .B2(n37700), .C1(n1841), 
        .C2(n26700), .ZN(n4186) );
  AOI22_X1 U4280 ( .A1(n16501), .A2(n31500), .B1(n2237), .B2(n4096), .ZN(n4185) );
  OAI221_X1 U4281 ( .B1(n2758), .B2(n2945), .C1(n1758), .C2(n3095), .A(n41901), 
        .ZN(n4096) );
  AOI22_X1 U4282 ( .A1(n45800), .A2(n1746), .B1(n21900), .B2(n3374), .ZN(
        n41901) );
  AND2_X1 U4283 ( .A1(n554), .A2(n2125), .ZN(n4138) );
  NOR2_X1 U4284 ( .A1(n2543), .A2(n2692), .ZN(n4187) );
  INV_X1 U4285 ( .A(n4093), .ZN(n4128) );
  NOR4_X1 U4286 ( .A1(N1228), .A2(n1347), .A3(n3466), .A4(N1229), .ZN(n4093)
         );
  AND3_X1 U4287 ( .A1(n3222), .A2(n3301), .A3(n15570), .ZN(n4191) );
  OAI22_X1 U4288 ( .A1(n2334), .A2(n2907), .B1(n3725), .B2(n1275), .ZN(N230)
         );
  INV_X1 U4289 ( .A(n4193), .ZN(n3725) );
  OAI211_X1 U4290 ( .C1(n1285), .C2(n1001), .A(n4195), .B(n4196), .ZN(n4193)
         );
  AOI221_X1 U4291 ( .B1(n38300), .B2(n2196), .C1(n46200), .C2(n2444), .A(n4199), .ZN(n4196) );
  OAI22_X1 U4292 ( .A1(n33101), .A2(n1468), .B1(n2779), .B2(n3147), .ZN(n4199)
         );
  AOI22_X1 U4293 ( .A1(n31900), .A2(n3411), .B1(n22100), .B2(n1776), .ZN(n4195) );
  OAI22_X1 U4294 ( .A1(n2339), .A2(n2909), .B1(n3728), .B2(n20001), .ZN(N229)
         );
  INV_X1 U4295 ( .A(n4203), .ZN(n3728) );
  OAI211_X1 U4296 ( .C1(n19701), .C2(n1002), .A(n4204), .B(n4205), .ZN(n4203)
         );
  AOI221_X1 U4297 ( .B1(n38900), .B2(n2198), .C1(n46800), .C2(n2447), .A(n4206), .ZN(n4205) );
  OAI22_X1 U4298 ( .A1(n2511), .A2(n1461), .B1(n20601), .B2(n3152), .ZN(n4206)
         );
  AOI22_X1 U4299 ( .A1(n32200), .A2(n549), .B1(n33), .B2(n1779), .ZN(n4204) );
  OAI22_X1 U4300 ( .A1(n2337), .A2(n2903), .B1(n37301), .B2(n10901), .ZN(N228)
         );
  INV_X1 U4301 ( .A(n4207), .ZN(n37301) );
  OAI211_X1 U4302 ( .C1(n1084), .C2(n999), .A(n4208), .B(n4209), .ZN(n4207) );
  AOI221_X1 U4303 ( .B1(n39400), .B2(n2201), .C1(n4730), .C2(n2411), .A(n42101), .ZN(n4209) );
  OAI22_X1 U4304 ( .A1(n2457), .A2(n1454), .B1(n1254), .B2(n31401), .ZN(n42101) );
  AOI22_X1 U4305 ( .A1(n32600), .A2(n3172), .B1(n32), .B2(n3208), .ZN(n4208)
         );
  OAI22_X1 U4306 ( .A1(n2344), .A2(n2905), .B1(n3732), .B2(n10901), .ZN(N227)
         );
  INV_X1 U4307 ( .A(n4211), .ZN(n3732) );
  OAI211_X1 U4308 ( .C1(n1084), .C2(n10001), .A(n4212), .B(n4213), .ZN(n4211)
         );
  AOI221_X1 U4309 ( .B1(n39900), .B2(n2195), .C1(n4780), .C2(n2405), .A(n4214), 
        .ZN(n4213) );
  OAI22_X1 U4310 ( .A1(n2451), .A2(n1447), .B1(n2059), .B2(n3144), .ZN(n4214)
         );
  AOI22_X1 U4311 ( .A1(n33000), .A2(n3168), .B1(n31), .B2(n3204), .ZN(n4212)
         );
  OAI22_X1 U4312 ( .A1(n2334), .A2(n2899), .B1(n3734), .B2(n2804), .ZN(N226)
         );
  INV_X1 U4313 ( .A(n4215), .ZN(n3734) );
  OAI211_X1 U4314 ( .C1(n2814), .C2(n997), .A(n4216), .B(n4217), .ZN(n4215) );
  AOI221_X1 U4315 ( .B1(n40100), .B2(n2199), .C1(n4840), .C2(n2438), .A(n4218), 
        .ZN(n4217) );
  OAI22_X1 U4316 ( .A1(n2521), .A2(n1442), .B1(n2056), .B2(n3132), .ZN(n4218)
         );
  AOI22_X1 U4317 ( .A1(n33400), .A2(n34101), .B1(n30), .B2(n3202), .ZN(n4216)
         );
  OAI22_X1 U4318 ( .A1(n23401), .A2(n2901), .B1(n3736), .B2(n2001), .ZN(N225)
         );
  INV_X1 U4319 ( .A(n4219), .ZN(n3736) );
  OAI211_X1 U4320 ( .C1(n1971), .C2(n998), .A(n42201), .B(n4221), .ZN(n4219)
         );
  AOI221_X1 U4321 ( .B1(n40900), .B2(n2201), .C1(n4880), .C2(n2441), .A(n4222), 
        .ZN(n4221) );
  OAI22_X1 U4322 ( .A1(n2518), .A2(n1435), .B1(n3362), .B2(n3136), .ZN(n4222)
         );
  AOI22_X1 U4323 ( .A1(n33800), .A2(n1786), .B1(n29), .B2(n15201), .ZN(n42201)
         );
  OAI22_X1 U4324 ( .A1(n2336), .A2(n2895), .B1(n3738), .B2(n3347), .ZN(N224)
         );
  INV_X1 U4325 ( .A(n4223), .ZN(n3738) );
  OAI211_X1 U4326 ( .C1(n3341), .C2(n995), .A(n4224), .B(n4225), .ZN(n4223) );
  AOI221_X1 U4327 ( .B1(n41400), .B2(n2195), .C1(n493), .C2(n2407), .A(n4226), 
        .ZN(n4225) );
  OAI22_X1 U4328 ( .A1(n2453), .A2(n1428), .B1(n3362), .B2(n3124), .ZN(n4226)
         );
  AOI22_X1 U4329 ( .A1(n34200), .A2(n3173), .B1(n28), .B2(n3209), .ZN(n4224)
         );
  OAI22_X1 U4330 ( .A1(n2343), .A2(n2897), .B1(n37401), .B2(n3347), .ZN(N223)
         );
  INV_X1 U4331 ( .A(n4227), .ZN(n37401) );
  OAI211_X1 U4332 ( .C1(n3341), .C2(n996), .A(n4228), .B(n4229), .ZN(n4227) );
  AOI221_X1 U4333 ( .B1(n41900), .B2(n2199), .C1(n498), .C2(n2402), .A(n42301), 
        .ZN(n4229) );
  OAI22_X1 U4334 ( .A1(n2448), .A2(n1421), .B1(n2056), .B2(n3128), .ZN(n42301)
         );
  AOI22_X1 U4335 ( .A1(n34600), .A2(n3169), .B1(n27), .B2(n3205), .ZN(n4228)
         );
  OAI22_X1 U4336 ( .A1(n2335), .A2(n2891), .B1(n3742), .B2(n1276), .ZN(N222)
         );
  INV_X1 U4337 ( .A(n4231), .ZN(n3742) );
  OAI211_X1 U4338 ( .C1(n1286), .C2(n993), .A(n4232), .B(n4233), .ZN(n4231) );
  AOI221_X1 U4339 ( .B1(n42100), .B2(n2202), .C1(n5040), .C2(n2443), .A(n4234), 
        .ZN(n4233) );
  OAI22_X1 U4340 ( .A1(n3309), .A2(n1416), .B1(n1253), .B2(n3116), .ZN(n4234)
         );
  AOI22_X1 U4341 ( .A1(n35000), .A2(n10601), .B1(n26), .B2(n3404), .ZN(n4232)
         );
  OAI22_X1 U4342 ( .A1(n2339), .A2(n2893), .B1(n3744), .B2(n20001), .ZN(N221)
         );
  INV_X1 U4343 ( .A(n4235), .ZN(n3744) );
  OAI211_X1 U4344 ( .C1(n19701), .C2(n994), .A(n4236), .B(n4237), .ZN(n4235)
         );
  AOI221_X1 U4345 ( .B1(n42900), .B2(n2196), .C1(n508), .C2(n2446), .A(n4238), 
        .ZN(n4237) );
  OAI22_X1 U4346 ( .A1(n2512), .A2(n1409), .B1(n20601), .B2(n31201), .ZN(n4238) );
  AOI22_X1 U4347 ( .A1(n35400), .A2(n3167), .B1(n25), .B2(n3405), .ZN(n4236)
         );
  OAI22_X1 U4348 ( .A1(n2336), .A2(n2887), .B1(n3746), .B2(n1695), .ZN(N220)
         );
  INV_X1 U4349 ( .A(n4239), .ZN(n3746) );
  OAI211_X1 U4350 ( .C1(n1677), .C2(n991), .A(n42401), .B(n4241), .ZN(n4239)
         );
  AOI221_X1 U4351 ( .B1(n43400), .B2(n2198), .C1(n513), .C2(n24101), .A(n4242), 
        .ZN(n4241) );
  OAI22_X1 U4352 ( .A1(n2456), .A2(n1404), .B1(n2779), .B2(n3108), .ZN(n4242)
         );
  AOI22_X1 U4353 ( .A1(n35800), .A2(n3174), .B1(n24), .B2(n32101), .ZN(n42401)
         );
  OAI22_X1 U4354 ( .A1(n2343), .A2(n2889), .B1(n3748), .B2(n1997), .ZN(N219)
         );
  INV_X1 U4355 ( .A(n4243), .ZN(n3748) );
  OAI211_X1 U4356 ( .C1(n1678), .C2(n992), .A(n4244), .B(n4245), .ZN(n4243) );
  AOI221_X1 U4357 ( .B1(n43900), .B2(n2202), .C1(n518), .C2(n2404), .A(n4246), 
        .ZN(n4245) );
  OAI22_X1 U4358 ( .A1(n24501), .A2(n1399), .B1(n2059), .B2(n3112), .ZN(n4246)
         );
  AOI22_X1 U4359 ( .A1(n36200), .A2(n31701), .B1(n23), .B2(n3206), .ZN(n4244)
         );
  OAI22_X1 U4360 ( .A1(n2335), .A2(n2883), .B1(n37501), .B2(n2804), .ZN(N218)
         );
  INV_X1 U4361 ( .A(n4247), .ZN(n37501) );
  OAI211_X1 U4362 ( .C1(n2814), .C2(n989), .A(n4248), .B(n4249), .ZN(n4247) );
  AOI221_X1 U4363 ( .B1(n44100), .B2(n2193), .C1(n524), .C2(n2437), .A(n42501), 
        .ZN(n4249) );
  OAI22_X1 U4364 ( .A1(n25201), .A2(n1394), .B1(n1734), .B2(n31001), .ZN(
        n42501) );
  AOI22_X1 U4365 ( .A1(n36600), .A2(n1789), .B1(n22), .B2(n3203), .ZN(n4248)
         );
  OAI22_X1 U4366 ( .A1(n23401), .A2(n2885), .B1(n3752), .B2(n2001), .ZN(N217)
         );
  INV_X1 U4367 ( .A(n4251), .ZN(n3752) );
  OAI211_X1 U4368 ( .C1(n1971), .C2(n990), .A(n4252), .B(n4253), .ZN(n4251) );
  AOI221_X1 U4369 ( .B1(n44900), .B2(n2192), .C1(n528), .C2(n24401), .A(n4254), 
        .ZN(n4253) );
  OAI22_X1 U4370 ( .A1(n2517), .A2(n1387), .B1(n1101), .B2(n3104), .ZN(n4254)
         );
  AOI22_X1 U4371 ( .A1(n37000), .A2(n15101), .B1(n21), .B2(n1062), .ZN(n4252)
         );
  OAI22_X1 U4372 ( .A1(n2337), .A2(n2879), .B1(n3754), .B2(n1997), .ZN(N216)
         );
  INV_X1 U4373 ( .A(n4255), .ZN(n3754) );
  OAI211_X1 U4374 ( .C1(n1967), .C2(n987), .A(n4256), .B(n4257), .ZN(n4255) );
  AOI221_X1 U4375 ( .B1(n45400), .B2(n2192), .C1(n533), .C2(n2406), .A(n4258), 
        .ZN(n4257) );
  OAI22_X1 U4376 ( .A1(n2452), .A2(n13801), .B1(n1101), .B2(n3092), .ZN(n4258)
         );
  AOI22_X1 U4377 ( .A1(n37400), .A2(n3175), .B1(n20), .B2(n3211), .ZN(n4256)
         );
  OAI22_X1 U4378 ( .A1(n2344), .A2(n2881), .B1(n3756), .B2(n1696), .ZN(N215)
         );
  INV_X1 U4379 ( .A(n4259), .ZN(n3756) );
  OAI211_X1 U4380 ( .C1(n1967), .C2(n988), .A(n42601), .B(n4261), .ZN(n4259)
         );
  AOI221_X1 U4381 ( .B1(n45900), .B2(n2193), .C1(n538), .C2(n2403), .A(n4262), 
        .ZN(n4261) );
  OAI22_X1 U4382 ( .A1(n2449), .A2(n1373), .B1(n1735), .B2(n3096), .ZN(n4262)
         );
  AOI22_X1 U4383 ( .A1(n37800), .A2(n3171), .B1(n19), .B2(n3207), .ZN(n42601)
         );
  OAI21_X1 U4384 ( .B1(n2524), .B2(n1275), .A(n1368), .ZN(n4263) );
  NAND2_X1 U4385 ( .A1(n2035), .A2(n37601), .ZN(n4192) );
  OR2_X1 U4386 ( .A1(n3796), .A2(n2212), .ZN(n37601) );
  OAI22_X1 U4387 ( .A1(n2349), .A2(n2875), .B1(n3763), .B2(n1269), .ZN(N214)
         );
  INV_X1 U4388 ( .A(n4266), .ZN(n3763) );
  OAI211_X1 U4389 ( .C1(n1017), .C2(n1263), .A(n4268), .B(n4269), .ZN(n4266)
         );
  AOI221_X1 U4390 ( .B1(n2441), .B2(n38100), .C1(n1199), .C2(n46400), .A(n4271), .ZN(n4269) );
  OAI22_X1 U4391 ( .A1(n1052), .A2(n2506), .B1(n3149), .B2(n2177), .ZN(n4271)
         );
  AOI22_X1 U4392 ( .A1(n1775), .A2(n31700), .B1(n3396), .B2(n34), .ZN(n4268)
         );
  OAI22_X1 U4393 ( .A1(n2346), .A2(n2877), .B1(n3766), .B2(n2005), .ZN(N213)
         );
  INV_X1 U4394 ( .A(n4273), .ZN(n3766) );
  OAI211_X1 U4395 ( .C1(n29101), .C2(n20301), .A(n4274), .B(n4275), .ZN(n4273)
         );
  AOI221_X1 U4396 ( .B1(n38700), .B2(n2443), .C1(n46600), .C2(n2706), .A(n4276), .ZN(n4275) );
  OAI22_X1 U4397 ( .A1(n2473), .A2(n1051), .B1(n2178), .B2(n3153), .ZN(n4276)
         );
  AOI22_X1 U4398 ( .A1(n32300), .A2(n1519), .B1(n22400), .B2(n3391), .ZN(n4274) );
  OAI22_X1 U4399 ( .A1(n2356), .A2(n2871), .B1(n3768), .B2(n1091), .ZN(N212)
         );
  INV_X1 U4400 ( .A(n4277), .ZN(n3768) );
  OAI211_X1 U4401 ( .C1(n1015), .C2(n3355), .A(n4278), .B(n4279), .ZN(n4277)
         );
  AOI221_X1 U4402 ( .B1(n39200), .B2(n2411), .C1(n4710), .C2(n3166), .A(n42801), .ZN(n4279) );
  OAI22_X1 U4403 ( .A1(n2503), .A2(n10501), .B1(n2456), .B2(n3141), .ZN(n42801) );
  AOI22_X1 U4404 ( .A1(n32700), .A2(n3405), .B1(n22700), .B2(n3236), .ZN(n4278) );
  OAI22_X1 U4405 ( .A1(n2353), .A2(n2873), .B1(n37701), .B2(n1091), .ZN(N211)
         );
  INV_X1 U4406 ( .A(n4281), .ZN(n37701) );
  OAI211_X1 U4407 ( .C1(n2906), .C2(n3355), .A(n4282), .B(n4283), .ZN(n4281)
         );
  AOI221_X1 U4408 ( .B1(n39700), .B2(n2405), .C1(n4760), .C2(n3162), .A(n4284), 
        .ZN(n4283) );
  OAI22_X1 U4409 ( .A1(n2507), .A2(n1049), .B1(n24501), .B2(n3145), .ZN(n4284)
         );
  AOI22_X1 U4410 ( .A1(n33100), .A2(n3208), .B1(n23000), .B2(n2919), .ZN(n4282) );
  OAI22_X1 U4411 ( .A1(n2349), .A2(n2867), .B1(n3772), .B2(n2798), .ZN(N210)
         );
  INV_X1 U4412 ( .A(n4285), .ZN(n3772) );
  OAI211_X1 U4413 ( .C1(n1013), .C2(n2792), .A(n4286), .B(n4287), .ZN(n4285)
         );
  AOI221_X1 U4414 ( .B1(n40200), .B2(n2446), .C1(n4810), .C2(n3155), .A(n4288), 
        .ZN(n4287) );
  OAI22_X1 U4415 ( .A1(n2487), .A2(n1048), .B1(n2512), .B2(n3133), .ZN(n4288)
         );
  AOI22_X1 U4416 ( .A1(n33500), .A2(n3202), .B1(n23300), .B2(n29301), .ZN(
        n4286) );
  OAI22_X1 U4417 ( .A1(n2347), .A2(n2869), .B1(n3774), .B2(n2006), .ZN(N209)
         );
  INV_X1 U4418 ( .A(n4289), .ZN(n3774) );
  OAI211_X1 U4419 ( .C1(n29020), .C2(n829), .A(n42901), .B(n4291), .ZN(n4289)
         );
  AOI221_X1 U4420 ( .B1(n40700), .B2(n2438), .C1(n4860), .C2(n3155), .A(n4292), 
        .ZN(n4291) );
  OAI22_X1 U4421 ( .A1(n2475), .A2(n1047), .B1(n2521), .B2(n3137), .ZN(n4292)
         );
  AOI22_X1 U4422 ( .A1(n33900), .A2(n3204), .B1(n23600), .B2(n21501), .ZN(
        n42901) );
  OAI22_X1 U4423 ( .A1(n2355), .A2(n2863), .B1(n3776), .B2(n3348), .ZN(N208)
         );
  INV_X1 U4424 ( .A(n4293), .ZN(n3776) );
  OAI211_X1 U4425 ( .C1(n2896), .C2(n3354), .A(n4294), .B(n4295), .ZN(n4293)
         );
  AOI221_X1 U4426 ( .B1(n41200), .B2(n2406), .C1(n4910), .C2(n3165), .A(n4296), 
        .ZN(n4295) );
  OAI22_X1 U4427 ( .A1(n2483), .A2(n1046), .B1(n2457), .B2(n3125), .ZN(n4296)
         );
  AOI22_X1 U4428 ( .A1(n34300), .A2(n1062), .B1(n23900), .B2(n3231), .ZN(n4294) );
  OAI22_X1 U4429 ( .A1(n2352), .A2(n2865), .B1(n3778), .B2(n3348), .ZN(N207)
         );
  INV_X1 U4430 ( .A(n4297), .ZN(n3778) );
  OAI211_X1 U4431 ( .C1(n1012), .C2(n3354), .A(n4298), .B(n4299), .ZN(n4297)
         );
  AOI221_X1 U4432 ( .B1(n41700), .B2(n2403), .C1(n496), .C2(n3161), .A(n43001), 
        .ZN(n4299) );
  OAI22_X1 U4433 ( .A1(n2509), .A2(n1045), .B1(n2453), .B2(n3129), .ZN(n43001)
         );
  AOI22_X1 U4434 ( .A1(n34700), .A2(n32001), .B1(n24200), .B2(n2921), .ZN(
        n4298) );
  OAI22_X1 U4435 ( .A1(n23501), .A2(n2859), .B1(n37801), .B2(n12701), .ZN(N206) );
  INV_X1 U4436 ( .A(n4301), .ZN(n37801) );
  OAI211_X1 U4437 ( .C1(n2892), .C2(n1264), .A(n4302), .B(n4303), .ZN(n4301)
         );
  AOI221_X1 U4438 ( .B1(n42200), .B2(n24401), .C1(n5010), .C2(n3158), .A(n4304), .ZN(n4303) );
  OAI22_X1 U4439 ( .A1(n2481), .A2(n1043), .B1(n2518), .B2(n3117), .ZN(n4304)
         );
  AOI22_X1 U4440 ( .A1(n35100), .A2(n3209), .B1(n24500), .B2(n2923), .ZN(n4302) );
  OAI22_X1 U4441 ( .A1(n2346), .A2(n2861), .B1(n3782), .B2(n2005), .ZN(N205)
         );
  INV_X1 U4442 ( .A(n4305), .ZN(n3782) );
  OAI211_X1 U4443 ( .C1(n2894), .C2(n20301), .A(n4306), .B(n4307), .ZN(n4305)
         );
  AOI221_X1 U4444 ( .B1(n42700), .B2(n2444), .C1(n506), .C2(n3157), .A(n4308), 
        .ZN(n4307) );
  OAI22_X1 U4445 ( .A1(n24701), .A2(n1042), .B1(n33101), .B2(n3121), .ZN(n4308) );
  AOI22_X1 U4446 ( .A1(n35500), .A2(n32101), .B1(n24800), .B2(n3389), .ZN(
        n4306) );
  OAI22_X1 U4447 ( .A1(n2356), .A2(n2855), .B1(n3784), .B2(n1698), .ZN(N204)
         );
  INV_X1 U4448 ( .A(n4309), .ZN(n3784) );
  OAI211_X1 U4449 ( .C1(n2888), .C2(n1715), .A(n43101), .B(n4311), .ZN(n4309)
         );
  AOI221_X1 U4450 ( .B1(n43200), .B2(n24101), .C1(n511), .C2(n3164), .A(n4312), 
        .ZN(n4311) );
  OAI22_X1 U4451 ( .A1(n2471), .A2(n10401), .B1(n2451), .B2(n3109), .ZN(n4312)
         );
  AOI22_X1 U4452 ( .A1(n35900), .A2(n3205), .B1(n25100), .B2(n33901), .ZN(
        n43101) );
  OAI22_X1 U4453 ( .A1(n2353), .A2(n2857), .B1(n3786), .B2(n1699), .ZN(N203)
         );
  INV_X1 U4454 ( .A(n4313), .ZN(n3786) );
  OAI211_X1 U4455 ( .C1(n28901), .C2(n2027), .A(n4314), .B(n4315), .ZN(n4313)
         );
  AOI221_X1 U4456 ( .B1(n43700), .B2(n2404), .C1(n516), .C2(n31601), .A(n4316), 
        .ZN(n4315) );
  OAI22_X1 U4457 ( .A1(n2502), .A2(n1038), .B1(n2448), .B2(n3113), .ZN(n4316)
         );
  AOI22_X1 U4458 ( .A1(n36300), .A2(n3404), .B1(n25400), .B2(n2917), .ZN(n4314) );
  OAI22_X1 U4459 ( .A1(n23501), .A2(n2851), .B1(n3788), .B2(n2798), .ZN(N202)
         );
  INV_X1 U4460 ( .A(n4317), .ZN(n3788) );
  OAI211_X1 U4461 ( .C1(n1005), .C2(n2792), .A(n4318), .B(n4319), .ZN(n4317)
         );
  AOI221_X1 U4462 ( .B1(n44200), .B2(n2447), .C1(n521), .C2(n11201), .A(n43201), .ZN(n4319) );
  OAI22_X1 U4463 ( .A1(n2504), .A2(n1036), .B1(n25201), .B2(n3101), .ZN(n43201) );
  AOI22_X1 U4464 ( .A1(n36700), .A2(n3206), .B1(n25700), .B2(n1771), .ZN(n4318) );
  OAI22_X1 U4465 ( .A1(n2347), .A2(n2853), .B1(n37901), .B2(n2006), .ZN(N201)
         );
  INV_X1 U4466 ( .A(n4321), .ZN(n37901) );
  OAI211_X1 U4467 ( .C1(n2886), .C2(n829), .A(n4322), .B(n4323), .ZN(n4321) );
  AOI221_X1 U4468 ( .B1(n44700), .B2(n2437), .C1(n526), .C2(n3434), .A(n4324), 
        .ZN(n4323) );
  OAI22_X1 U4469 ( .A1(n2482), .A2(n1035), .B1(n2511), .B2(n3105), .ZN(n4324)
         );
  AOI22_X1 U4470 ( .A1(n37100), .A2(n1778), .B1(n26000), .B2(n21001), .ZN(
        n4322) );
  OAI22_X1 U4471 ( .A1(n2355), .A2(n2847), .B1(n3792), .B2(n2002), .ZN(N200)
         );
  INV_X1 U4472 ( .A(n4325), .ZN(n3792) );
  OAI211_X1 U4473 ( .C1(n28801), .C2(n2027), .A(n4326), .B(n4327), .ZN(n4325)
         );
  AOI221_X1 U4474 ( .B1(n45200), .B2(n2407), .C1(n531), .C2(n3163), .A(n4328), 
        .ZN(n4327) );
  OAI22_X1 U4475 ( .A1(n2479), .A2(n1034), .B1(n2452), .B2(n3093), .ZN(n4328)
         );
  AOI22_X1 U4476 ( .A1(n37500), .A2(n3211), .B1(n26300), .B2(n2155), .ZN(n4326) );
  OAI22_X1 U4477 ( .A1(n2352), .A2(n2849), .B1(n3794), .B2(n2002), .ZN(N199)
         );
  INV_X1 U4478 ( .A(n4329), .ZN(n3794) );
  OAI211_X1 U4479 ( .C1(n2882), .C2(n1716), .A(n43301), .B(n4331), .ZN(n4329)
         );
  AOI221_X1 U4480 ( .B1(n45700), .B2(n2402), .C1(n536), .C2(n3159), .A(n4332), 
        .ZN(n4331) );
  OAI22_X1 U4481 ( .A1(n2485), .A2(n1033), .B1(n2449), .B2(n3097), .ZN(n4332)
         );
  NOR3_X1 U4482 ( .A1(n2943), .A2(n3241), .A3(n12301), .ZN(n4198) );
  AOI22_X1 U4483 ( .A1(n37900), .A2(n3207), .B1(n26600), .B2(n3397), .ZN(
        n43301) );
  OAI22_X1 U4484 ( .A1(n2524), .A2(n1269), .B1(n26801), .B2(n1032), .ZN(n4333)
         );
  NAND2_X1 U4485 ( .A1(n17201), .A2(n583), .ZN(n4265) );
  OR2_X1 U4486 ( .A1(n2681), .A2(n1187), .ZN(n3796) );
  OAI22_X1 U4487 ( .A1(n2311), .A2(n985), .B1(n3798), .B2(n1279), .ZN(N198) );
  INV_X1 U4488 ( .A(n4335), .ZN(n3798) );
  OAI211_X1 U4489 ( .C1(n2908), .C2(n1196), .A(n4336), .B(n4337), .ZN(n4335)
         );
  AOI221_X1 U4490 ( .B1(n12001), .B2(n38200), .C1(n3407), .C2(n46100), .A(
        n4339), .ZN(n4337) );
  OAI22_X1 U4491 ( .A1(n3008), .A2(n2934), .B1(n3148), .B2(n2484), .ZN(n4339)
         );
  AOI22_X1 U4492 ( .A1(n1529), .A2(n31800), .B1(n2749), .B2(n12200), .ZN(n4336) );
  OAI22_X1 U4493 ( .A1(n2317), .A2(n986), .B1(n3801), .B2(n19901), .ZN(N197)
         );
  INV_X1 U4494 ( .A(n4341), .ZN(n3801) );
  OAI211_X1 U4495 ( .C1(n1018), .C2(n1055), .A(n4342), .B(n4343), .ZN(n4341)
         );
  AOI221_X1 U4496 ( .B1(n38800), .B2(n2706), .C1(n46700), .C2(n1783), .A(n4344), .ZN(n4343) );
  OAI22_X1 U4497 ( .A1(n2934), .A2(n3006), .B1(n2487), .B2(n3151), .ZN(n4344)
         );
  AOI22_X1 U4498 ( .A1(n32100), .A2(n1022), .B1(n1489), .B2(n12400), .ZN(n4342) );
  OAI22_X1 U4499 ( .A1(n2315), .A2(n983), .B1(n3803), .B2(n1088), .ZN(N196) );
  INV_X1 U4500 ( .A(n4345), .ZN(n3803) );
  OAI211_X1 U4501 ( .C1(n2904), .C2(n2699), .A(n4346), .B(n4347), .ZN(n4345)
         );
  AOI221_X1 U4502 ( .B1(n39300), .B2(n3166), .C1(n4720), .C2(n3196), .A(n4348), 
        .ZN(n4347) );
  OAI22_X1 U4503 ( .A1(n2098), .A2(n3002), .B1(n2471), .B2(n3139), .ZN(n4348)
         );
  AOI22_X1 U4504 ( .A1(n32500), .A2(n2107), .B1(n20901), .B2(n12600), .ZN(
        n4346) );
  OAI22_X1 U4505 ( .A1(n2322), .A2(n984), .B1(n3805), .B2(n1088), .ZN(N195) );
  INV_X1 U4506 ( .A(n4349), .ZN(n3805) );
  OAI211_X1 U4507 ( .C1(n1016), .C2(n3011), .A(n43501), .B(n4351), .ZN(n4349)
         );
  AOI221_X1 U4508 ( .B1(n39800), .B2(n3162), .C1(n4770), .C2(n3192), .A(n4352), 
        .ZN(n4351) );
  OAI22_X1 U4509 ( .A1(n2094), .A2(n2998), .B1(n2501), .B2(n3143), .ZN(n4352)
         );
  AOI22_X1 U4510 ( .A1(n32900), .A2(n33901), .B1(n2086), .B2(n12800), .ZN(
        n43501) );
  OAI22_X1 U4511 ( .A1(n2311), .A2(n981), .B1(n3807), .B2(n2808), .ZN(N194) );
  INV_X1 U4512 ( .A(n4353), .ZN(n3807) );
  OAI211_X1 U4513 ( .C1(n29001), .C2(n1201), .A(n4354), .B(n4355), .ZN(n4353)
         );
  AOI221_X1 U4514 ( .B1(n40300), .B2(n1507), .C1(n4820), .C2(n17801), .A(n4356), .ZN(n4355) );
  OAI22_X1 U4515 ( .A1(n2937), .A2(n2994), .B1(n2504), .B2(n3131), .ZN(n4356)
         );
  AOI22_X1 U4516 ( .A1(n33300), .A2(n2156), .B1(n3023), .B2(n13000), .ZN(n4354) );
  OAI22_X1 U4517 ( .A1(n2318), .A2(n982), .B1(n3809), .B2(n1991), .ZN(N193) );
  INV_X1 U4518 ( .A(n4357), .ZN(n3809) );
  OAI211_X1 U4519 ( .C1(n1014), .C2(n11901), .A(n4358), .B(n4359), .ZN(n4357)
         );
  AOI221_X1 U4520 ( .B1(n40800), .B2(n1508), .C1(n4870), .C2(n31901), .A(
        n43601), .ZN(n4359) );
  OAI22_X1 U4521 ( .A1(n2928), .A2(n29901), .B1(n2481), .B2(n3135), .ZN(n43601) );
  AOI22_X1 U4522 ( .A1(n33700), .A2(n1023), .B1(n2741), .B2(n13200), .ZN(n4358) );
  OAI22_X1 U4523 ( .A1(n2314), .A2(n979), .B1(n3811), .B2(n3345), .ZN(N192) );
  INV_X1 U4524 ( .A(n4361), .ZN(n3811) );
  OAI211_X1 U4525 ( .C1(n1011), .C2(n1475), .A(n4362), .B(n4363), .ZN(n4361)
         );
  AOI221_X1 U4526 ( .B1(n41300), .B2(n3165), .C1(n4920), .C2(n3197), .A(n4364), 
        .ZN(n4363) );
  OAI22_X1 U4527 ( .A1(n1027), .A2(n2986), .B1(n2483), .B2(n3123), .ZN(n4364)
         );
  AOI22_X1 U4528 ( .A1(n34100), .A2(n1026), .B1(n1058), .B2(n13400), .ZN(n4362) );
  OAI22_X1 U4529 ( .A1(n2321), .A2(n980), .B1(n3813), .B2(n3345), .ZN(N191) );
  INV_X1 U4530 ( .A(n4365), .ZN(n3813) );
  OAI211_X1 U4531 ( .C1(n2898), .C2(n1198), .A(n4366), .B(n4367), .ZN(n4365)
         );
  AOI221_X1 U4532 ( .B1(n41800), .B2(n3161), .C1(n497), .C2(n3193), .A(n4368), 
        .ZN(n4367) );
  OAI22_X1 U4533 ( .A1(n2097), .A2(n2982), .B1(n2478), .B2(n3127), .ZN(n4368)
         );
  AOI22_X1 U4534 ( .A1(n34500), .A2(n2151), .B1(n550), .B2(n13600), .ZN(n4366)
         );
  OAI22_X1 U4535 ( .A1(n2312), .A2(n977), .B1(n3815), .B2(n12801), .ZN(N190)
         );
  INV_X1 U4536 ( .A(n4369), .ZN(n3815) );
  OAI211_X1 U4537 ( .C1(n1009), .C2(n3013), .A(n43701), .B(n4371), .ZN(n4369)
         );
  AOI221_X1 U4538 ( .B1(n42300), .B2(n3158), .C1(n5020), .C2(n3406), .A(n4372), 
        .ZN(n4371) );
  OAI22_X1 U4539 ( .A1(n2737), .A2(n2978), .B1(n2507), .B2(n3115), .ZN(n4372)
         );
  AOI22_X1 U4540 ( .A1(n34900), .A2(n2588), .B1(n2087), .B2(n13800), .ZN(
        n43701) );
  OAI22_X1 U4541 ( .A1(n2317), .A2(n978), .B1(n3817), .B2(n19901), .ZN(N189)
         );
  INV_X1 U4542 ( .A(n4373), .ZN(n3817) );
  OAI211_X1 U4543 ( .C1(n10101), .C2(n1485), .A(n4374), .B(n4375), .ZN(n4373)
         );
  AOI221_X1 U4544 ( .B1(n42800), .B2(n3157), .C1(n507), .C2(n1061), .A(n4376), 
        .ZN(n4375) );
  OAI22_X1 U4545 ( .A1(n1767), .A2(n2974), .B1(n2472), .B2(n3119), .ZN(n4376)
         );
  AOI22_X1 U4546 ( .A1(n35300), .A2(n2112), .B1(n1222), .B2(n14000), .ZN(n4374) );
  OAI22_X1 U4547 ( .A1(n2314), .A2(n975), .B1(n3819), .B2(n1689), .ZN(N188) );
  INV_X1 U4548 ( .A(n4377), .ZN(n3819) );
  OAI211_X1 U4549 ( .C1(n1007), .C2(n1053), .A(n4378), .B(n4379), .ZN(n4377)
         );
  AOI221_X1 U4550 ( .B1(n43300), .B2(n3164), .C1(n512), .C2(n3198), .A(n43801), 
        .ZN(n4379) );
  OAI22_X1 U4551 ( .A1(n2726), .A2(n29701), .B1(n2484), .B2(n3107), .ZN(n43801) );
  AOI22_X1 U4552 ( .A1(n35700), .A2(n1024), .B1(n2084), .B2(n14200), .ZN(n4378) );
  OAI22_X1 U4553 ( .A1(n2321), .A2(n976), .B1(n3821), .B2(n16901), .ZN(N187)
         );
  INV_X1 U4554 ( .A(n4381), .ZN(n3821) );
  OAI211_X1 U4555 ( .C1(n1008), .C2(n1479), .A(n4382), .B(n4383), .ZN(n4381)
         );
  AOI221_X1 U4556 ( .B1(n43800), .B2(n31601), .C1(n517), .C2(n3194), .A(n4384), 
        .ZN(n4383) );
  OAI22_X1 U4557 ( .A1(n2732), .A2(n2966), .B1(n2474), .B2(n3111), .ZN(n4384)
         );
  AOI22_X1 U4558 ( .A1(n36100), .A2(n3391), .B1(n1714), .B2(n14400), .ZN(n4382) );
  OAI22_X1 U4559 ( .A1(n2312), .A2(n973), .B1(n3823), .B2(n2808), .ZN(N186) );
  INV_X1 U4560 ( .A(n4385), .ZN(n3823) );
  OAI211_X1 U4561 ( .C1(n2884), .C2(n3014), .A(n4386), .B(n4387), .ZN(n4385)
         );
  AOI221_X1 U4562 ( .B1(n44300), .B2(n3434), .C1(n522), .C2(n3188), .A(n4388), 
        .ZN(n4387) );
  OAI22_X1 U4563 ( .A1(n2734), .A2(n2962), .B1(n2508), .B2(n3099), .ZN(n4388)
         );
  AOI22_X1 U4564 ( .A1(n36500), .A2(n3237), .B1(n1224), .B2(n14600), .ZN(n4386) );
  OAI22_X1 U4565 ( .A1(n2318), .A2(n974), .B1(n3825), .B2(n1991), .ZN(N185) );
  INV_X1 U4566 ( .A(n4389), .ZN(n3825) );
  OAI211_X1 U4567 ( .C1(n1006), .C2(n1488), .A(n43901), .B(n4391), .ZN(n4389)
         );
  AOI221_X1 U4568 ( .B1(n44800), .B2(n3433), .C1(n527), .C2(n1516), .A(n4392), 
        .ZN(n4391) );
  OAI22_X1 U4569 ( .A1(n2736), .A2(n2958), .B1(n2502), .B2(n3103), .ZN(n4392)
         );
  AOI22_X1 U4570 ( .A1(n36900), .A2(n2916), .B1(n3379), .B2(n14800), .ZN(
        n43901) );
  OAI22_X1 U4571 ( .A1(n2315), .A2(n971), .B1(n3827), .B2(n1987), .ZN(N184) );
  INV_X1 U4572 ( .A(n4393), .ZN(n3827) );
  OAI211_X1 U4573 ( .C1(n1003), .C2(n1054), .A(n4394), .B(n4395), .ZN(n4393)
         );
  AOI221_X1 U4574 ( .B1(n45300), .B2(n3163), .C1(n532), .C2(n3199), .A(n4396), 
        .ZN(n4395) );
  OAI22_X1 U4575 ( .A1(n2935), .A2(n2954), .B1(n2486), .B2(n3091), .ZN(n4396)
         );
  AOI22_X1 U4576 ( .A1(n37300), .A2(n2925), .B1(n12201), .B2(n15000), .ZN(
        n4394) );
  OAI22_X1 U4577 ( .A1(n2322), .A2(n972), .B1(n3829), .B2(n1987), .ZN(N183) );
  INV_X1 U4578 ( .A(n4397), .ZN(n3829) );
  OAI211_X1 U4579 ( .C1(n1004), .C2(n1482), .A(n4398), .B(n4399), .ZN(n4397)
         );
  AOI221_X1 U4580 ( .B1(n45800), .B2(n3159), .C1(n537), .C2(n3195), .A(n44001), 
        .ZN(n4399) );
  OAI22_X1 U4581 ( .A1(n2731), .A2(n29501), .B1(n24801), .B2(n3095), .ZN(
        n44001) );
  INV_X1 U4582 ( .A(n1253), .ZN(n42701) );
  NAND3_X1 U4583 ( .A1(n35), .A2(n1567), .A3(n2753), .ZN(n4201) );
  AOI22_X1 U4584 ( .A1(n37700), .A2(n2155), .B1(n3025), .B2(n15200), .ZN(n4398) );
  OAI22_X1 U4585 ( .A1(n2531), .A2(n1279), .B1(n3831), .B2(n2946), .ZN(n4401)
         );
  NOR2_X1 U4586 ( .A1(n1617), .A2(n1569), .ZN(n3831) );
  NAND2_X1 U4587 ( .A1(n2031), .A2(n3832), .ZN(n4334) );
  INV_X1 U4588 ( .A(n4402), .ZN(n3832) );
  AOI21_X1 U4589 ( .B1(n2211), .B2(n1186), .A(n2682), .ZN(n4402) );
  OAI22_X1 U4590 ( .A1(n2326), .A2(n563), .B1(n3834), .B2(n1273), .ZN(N182) );
  INV_X1 U4591 ( .A(n4405), .ZN(n3834) );
  OAI211_X1 U4592 ( .C1(n2876), .C2(n3009), .A(n4406), .B(n4407), .ZN(n4405)
         );
  AOI221_X1 U4593 ( .B1(n1781), .B2(n38400), .C1(n1787), .C2(n46300), .A(n4408), .ZN(n4407) );
  OAI22_X1 U4594 ( .A1(n2907), .A2(n2462), .B1(n31501), .B2(n2937), .ZN(n4408)
         );
  INV_X1 U4595 ( .A(n18), .ZN(n3724) );
  AOI22_X1 U4596 ( .A1(n2926), .A2(n15970), .B1(n3378), .B2(n22200), .ZN(n4406) );
  OAI22_X1 U4597 ( .A1(n2323), .A2(n560), .B1(n3837), .B2(n1995), .ZN(N181) );
  INV_X1 U4598 ( .A(n4409), .ZN(n3837) );
  OAI211_X1 U4599 ( .C1(n2878), .C2(n1056), .A(n44101), .B(n4411), .ZN(n4409)
         );
  AOI221_X1 U4600 ( .B1(n38600), .B2(n31901), .C1(n46900), .C2(n549), .A(n4412), .ZN(n4411) );
  OAI22_X1 U4601 ( .A1(n2909), .A2(n2434), .B1(n2932), .B2(n3154), .ZN(n4412)
         );
  INV_X1 U4602 ( .A(n27200), .ZN(n3727) );
  AOI22_X1 U4603 ( .A1(n16390), .A2(n29201), .B1(n3026), .B2(n22500), .ZN(
        n44101) );
  OAI22_X1 U4604 ( .A1(n2332), .A2(n561), .B1(n3839), .B2(n1089), .ZN(N180) );
  INV_X1 U4605 ( .A(n4413), .ZN(n3839) );
  OAI211_X1 U4606 ( .C1(n2872), .C2(n30101), .A(n4414), .B(n4415), .ZN(n4413)
         );
  AOI221_X1 U4607 ( .B1(n39100), .B2(n1784), .C1(n4740), .C2(n17901), .A(n4416), .ZN(n4415) );
  OAI22_X1 U4608 ( .A1(n2903), .A2(n2465), .B1(n2935), .B2(n3142), .ZN(n4416)
         );
  INV_X1 U4609 ( .A(n27500), .ZN(n3729) );
  AOI22_X1 U4610 ( .A1(n16700), .A2(n2918), .B1(n3025), .B2(n22800), .ZN(n4414) );
  OAI22_X1 U4611 ( .A1(n2329), .A2(n562), .B1(n3841), .B2(n1089), .ZN(N179) );
  INV_X1 U4612 ( .A(n4417), .ZN(n3841) );
  OAI211_X1 U4613 ( .C1(n2874), .C2(n3012), .A(n4418), .B(n4419), .ZN(n4417)
         );
  AOI221_X1 U4614 ( .B1(n39600), .B2(n3407), .C1(n4790), .C2(n34101), .A(
        n44201), .ZN(n4419) );
  OAI22_X1 U4615 ( .A1(n2905), .A2(n2428), .B1(n2097), .B2(n3146), .ZN(n44201)
         );
  INV_X1 U4616 ( .A(n27800), .ZN(n3731) );
  AOI22_X1 U4617 ( .A1(n17100), .A2(n2931), .B1(n2748), .B2(n23100), .ZN(n4418) );
  OAI22_X1 U4618 ( .A1(n2326), .A2(n567), .B1(n3843), .B2(n2802), .ZN(N178) );
  INV_X1 U4619 ( .A(n4421), .ZN(n3843) );
  OAI211_X1 U4620 ( .C1(n2868), .C2(n1195), .A(n4422), .B(n4423), .ZN(n4421)
         );
  AOI221_X1 U4621 ( .B1(n40400), .B2(n3198), .C1(n4830), .C2(n3174), .A(n4424), 
        .ZN(n4423) );
  OAI22_X1 U4622 ( .A1(n2899), .A2(n2469), .B1(n2928), .B2(n3134), .ZN(n4424)
         );
  INV_X1 U4623 ( .A(n28100), .ZN(n3733) );
  AOI22_X1 U4624 ( .A1(n17500), .A2(n2923), .B1(n12250), .B2(n23400), .ZN(
        n4422) );
  OAI22_X1 U4625 ( .A1(n2324), .A2(n564), .B1(n3845), .B2(n1996), .ZN(N177) );
  INV_X1 U4626 ( .A(n4425), .ZN(n3845) );
  OAI211_X1 U4627 ( .C1(n28701), .C2(n2708), .A(n4426), .B(n4427), .ZN(n4425)
         );
  AOI221_X1 U4628 ( .B1(n40600), .B2(n3194), .C1(n4890), .C2(n31701), .A(n4428), .ZN(n4427) );
  OAI22_X1 U4629 ( .A1(n2901), .A2(n2435), .B1(n2093), .B2(n3138), .ZN(n4428)
         );
  INV_X1 U4630 ( .A(n28400), .ZN(n3735) );
  AOI22_X1 U4631 ( .A1(n17900), .A2(n3238), .B1(n1492), .B2(n23700), .ZN(n4426) );
  OAI22_X1 U4632 ( .A1(n2331), .A2(n565), .B1(n3847), .B2(n3346), .ZN(N176) );
  INV_X1 U4633 ( .A(n4429), .ZN(n3847) );
  OAI211_X1 U4634 ( .C1(n2864), .C2(n2704), .A(n44301), .B(n4431), .ZN(n4429)
         );
  AOI221_X1 U4635 ( .B1(n41100), .B2(n3406), .C1(n494), .C2(n3411), .A(n4432), 
        .ZN(n4431) );
  OAI22_X1 U4636 ( .A1(n2895), .A2(n2459), .B1(n2726), .B2(n3126), .ZN(n4432)
         );
  INV_X1 U4637 ( .A(n28700), .ZN(n3737) );
  AOI22_X1 U4638 ( .A1(n18300), .A2(n2587), .B1(n3382), .B2(n24000), .ZN(
        n44301) );
  OAI22_X1 U4639 ( .A1(n2328), .A2(n566), .B1(n3849), .B2(n3346), .ZN(N175) );
  INV_X1 U4640 ( .A(n4433), .ZN(n3849) );
  OAI211_X1 U4641 ( .C1(n2866), .C2(n1189), .A(n4434), .B(n4435), .ZN(n4433)
         );
  AOI221_X1 U4642 ( .B1(n41600), .B2(n3191), .C1(n4990), .C2(n1511), .A(n4436), 
        .ZN(n4435) );
  OAI22_X1 U4643 ( .A1(n2897), .A2(n2427), .B1(n1029), .B2(n31301), .ZN(n4436)
         );
  INV_X1 U4644 ( .A(n29000), .ZN(n3739) );
  AOI22_X1 U4645 ( .A1(n18700), .A2(n3397), .B1(n2083), .B2(n24300), .ZN(n4434) );
  OAI22_X1 U4646 ( .A1(n2327), .A2(n571), .B1(n3851), .B2(n1274), .ZN(N174) );
  INV_X1 U4647 ( .A(n4437), .ZN(n3851) );
  OAI211_X1 U4648 ( .C1(n28601), .C2(n3009), .A(n4438), .B(n4439), .ZN(n4437)
         );
  AOI221_X1 U4649 ( .B1(n42400), .B2(n3196), .C1(n5030), .C2(n3172), .A(n44401), .ZN(n4439) );
  OAI22_X1 U4650 ( .A1(n2891), .A2(n2468), .B1(n2731), .B2(n3118), .ZN(n44401)
         );
  INV_X1 U4651 ( .A(n29300), .ZN(n3741) );
  AOI22_X1 U4652 ( .A1(n19100), .A2(n3231), .B1(n1223), .B2(n24600), .ZN(n4438) );
  OAI22_X1 U4653 ( .A1(n2323), .A2(n568), .B1(n3853), .B2(n1995), .ZN(N173) );
  INV_X1 U4654 ( .A(n4441), .ZN(n3853) );
  OAI211_X1 U4655 ( .C1(n2862), .C2(n683), .A(n4442), .B(n4443), .ZN(n4441) );
  AOI221_X1 U4656 ( .B1(n42600), .B2(n3199), .C1(n509), .C2(n3175), .A(n4444), 
        .ZN(n4443) );
  OAI22_X1 U4657 ( .A1(n2893), .A2(n2429), .B1(n2091), .B2(n3122), .ZN(n4444)
         );
  INV_X1 U4658 ( .A(n29600), .ZN(n3743) );
  AOI22_X1 U4659 ( .A1(n19500), .A2(n1771), .B1(n1059), .B2(n24900), .ZN(n4442) );
  OAI22_X1 U4660 ( .A1(n2332), .A2(n569), .B1(n3855), .B2(n1692), .ZN(N172) );
  INV_X1 U4661 ( .A(n4445), .ZN(n3855) );
  OAI211_X1 U4662 ( .C1(n2856), .C2(n30101), .A(n4446), .B(n4447), .ZN(n4445)
         );
  AOI221_X1 U4663 ( .B1(n43100), .B2(n3192), .C1(n514), .C2(n3168), .A(n4448), 
        .ZN(n4447) );
  OAI22_X1 U4664 ( .A1(n2887), .A2(n24601), .B1(n3386), .B2(n31101), .ZN(n4448) );
  INV_X1 U4665 ( .A(n29900), .ZN(n3745) );
  AOI22_X1 U4666 ( .A1(n19900), .A2(n21501), .B1(n1504), .B2(n25200), .ZN(
        n4446) );
  OAI22_X1 U4667 ( .A1(n2329), .A2(n570), .B1(n3857), .B2(n1992), .ZN(N171) );
  INV_X1 U4668 ( .A(n4449), .ZN(n3857) );
  OAI211_X1 U4669 ( .C1(n2858), .C2(n1476), .A(n44501), .B(n4451), .ZN(n4449)
         );
  AOI221_X1 U4670 ( .B1(n43600), .B2(n3195), .C1(n519), .C2(n3171), .A(n4452), 
        .ZN(n4451) );
  OAI22_X1 U4671 ( .A1(n2889), .A2(n2424), .B1(n2723), .B2(n3114), .ZN(n4452)
         );
  INV_X1 U4672 ( .A(n30200), .ZN(n3747) );
  AOI22_X1 U4673 ( .A1(n20300), .A2(n3233), .B1(n3015), .B2(n25500), .ZN(
        n44501) );
  OAI22_X1 U4674 ( .A1(n2327), .A2(n575), .B1(n3859), .B2(n2802), .ZN(N170) );
  INV_X1 U4675 ( .A(n4453), .ZN(n3859) );
  OAI211_X1 U4676 ( .C1(n2852), .C2(n559), .A(n4454), .B(n4455), .ZN(n4453) );
  AOI221_X1 U4677 ( .B1(n44400), .B2(n1061), .C1(n523), .C2(n10601), .A(n4456), 
        .ZN(n4455) );
  OAI22_X1 U4678 ( .A1(n2883), .A2(n2463), .B1(n1027), .B2(n3102), .ZN(n4456)
         );
  INV_X1 U4679 ( .A(n30500), .ZN(n3749) );
  AOI22_X1 U4680 ( .A1(n20700), .A2(n2922), .B1(n2087), .B2(n25800), .ZN(n4454) );
  OAI22_X1 U4681 ( .A1(n2324), .A2(n572), .B1(n3861), .B2(n1996), .ZN(N169) );
  INV_X1 U4682 ( .A(n4457), .ZN(n3861) );
  OAI211_X1 U4683 ( .C1(n2854), .C2(n1202), .A(n4458), .B(n4459), .ZN(n4457)
         );
  AOI221_X1 U4684 ( .B1(n44600), .B2(n1517), .C1(n529), .C2(n1511), .A(n44601), 
        .ZN(n4459) );
  OAI22_X1 U4685 ( .A1(n2885), .A2(n24301), .B1(n1768), .B2(n3106), .ZN(n44601) );
  INV_X1 U4686 ( .A(n30800), .ZN(n3751) );
  AOI22_X1 U4687 ( .A1(n21100), .A2(n2924), .B1(n2149), .B2(n26100), .ZN(n4458) );
  OAI22_X1 U4688 ( .A1(n2331), .A2(n573), .B1(n3863), .B2(n1992), .ZN(N168) );
  INV_X1 U4689 ( .A(n4461), .ZN(n3863) );
  OAI211_X1 U4690 ( .C1(n2848), .C2(n2704), .A(n4462), .B(n4463), .ZN(n4461)
         );
  AOI221_X1 U4691 ( .B1(n45100), .B2(n3197), .C1(n534), .C2(n3173), .A(n4464), 
        .ZN(n4463) );
  OAI22_X1 U4692 ( .A1(n2879), .A2(n2466), .B1(n2736), .B2(n3094), .ZN(n4464)
         );
  INV_X1 U4693 ( .A(n31100), .ZN(n3753) );
  AOI22_X1 U4694 ( .A1(n21500), .A2(n3392), .B1(n1495), .B2(n26400), .ZN(n4462) );
  OAI22_X1 U4695 ( .A1(n2328), .A2(n574), .B1(n3865), .B2(n1693), .ZN(N167) );
  INV_X1 U4696 ( .A(n4465), .ZN(n3865) );
  OAI211_X1 U4697 ( .C1(n28501), .C2(n11901), .A(n4466), .B(n4467), .ZN(n4465)
         );
  AOI221_X1 U4698 ( .B1(n45600), .B2(n3193), .C1(n539), .C2(n3169), .A(n4468), 
        .ZN(n4467) );
  OAI22_X1 U4699 ( .A1(n2881), .A2(n2425), .B1(n3388), .B2(n3098), .ZN(n4468)
         );
  INV_X1 U4700 ( .A(n31400), .ZN(n3755) );
  NAND2_X1 U4701 ( .A1(n1291), .A2(n545), .ZN(n42001) );
  AOI22_X1 U4702 ( .A1(n21900), .A2(n2101), .B1(n2742), .B2(n26700), .ZN(n4466) );
  OAI22_X1 U4703 ( .A1(n3306), .A2(n1273), .B1(n3867), .B2(n1368), .ZN(n4469)
         );
  NOR2_X1 U4704 ( .A1(n1245), .A2(n15631), .ZN(n3867) );
  NAND2_X1 U4705 ( .A1(n579), .A2(n2682), .ZN(n4404) );
  OAI22_X1 U4706 ( .A1(n2287), .A2(n3008), .B1(n38701), .B2(n1283), .ZN(N166)
         );
  INV_X1 U4707 ( .A(n4471), .ZN(n38701) );
  OAI211_X1 U4708 ( .C1(n2844), .C2(n3013), .A(n4472), .B(n4473), .ZN(n4471)
         );
  AOI221_X1 U4709 ( .B1(n25001), .B2(n27000), .C1(n3409), .C2(n54), .A(n4475), 
        .ZN(n4473) );
  OAI22_X1 U4710 ( .A1(n3003), .A2(n2929), .B1(n3083), .B2(n2478), .ZN(n4475)
         );
  AOI22_X1 U4711 ( .A1(n2113), .A2(n55), .B1(n2739), .B2(n31900), .ZN(n4472)
         );
  OAI22_X1 U4712 ( .A1(n2292), .A2(n3006), .B1(n3873), .B2(n19801), .ZN(N165)
         );
  INV_X1 U4713 ( .A(n4476), .ZN(n3873) );
  OAI211_X1 U4714 ( .C1(n2846), .C2(n1471), .A(n4477), .B(n4478), .ZN(n4476)
         );
  AOI221_X1 U4715 ( .B1(n2489), .B2(n27300), .C1(n3176), .C2(n53), .A(n4479), 
        .ZN(n4478) );
  OAI22_X1 U4716 ( .A1(n1112), .A2(n2999), .B1(n2475), .B2(n3087), .ZN(n4479)
         );
  AOI22_X1 U4717 ( .A1(n57), .A2(n3225), .B1(n2084), .B2(n32300), .ZN(n4477)
         );
  OAI22_X1 U4718 ( .A1(n22901), .A2(n3002), .B1(n3875), .B2(n1086), .ZN(N164)
         );
  INV_X1 U4719 ( .A(n44801), .ZN(n3875) );
  OAI211_X1 U4720 ( .C1(n28401), .C2(n3011), .A(n4481), .B(n4482), .ZN(n44801)
         );
  AOI221_X1 U4721 ( .B1(n2492), .B2(n27600), .C1(n3184), .C2(n52), .A(n4483), 
        .ZN(n4482) );
  OAI22_X1 U4722 ( .A1(n1029), .A2(n2995), .B1(n2508), .B2(n3075), .ZN(n4483)
         );
  AOI22_X1 U4723 ( .A1(n59), .A2(n3233), .B1(n11101), .B2(n32700), .ZN(n4481)
         );
  OAI22_X1 U4724 ( .A1(n2297), .A2(n2998), .B1(n3877), .B2(n1086), .ZN(N163)
         );
  INV_X1 U4725 ( .A(n4484), .ZN(n3877) );
  OAI211_X1 U4726 ( .C1(n2842), .C2(n2207), .A(n4485), .B(n4486), .ZN(n4484)
         );
  AOI221_X1 U4727 ( .B1(n2495), .B2(n27900), .C1(n3183), .C2(n51), .A(n4487), 
        .ZN(n4486) );
  OAI22_X1 U4728 ( .A1(n3388), .A2(n2991), .B1(n24701), .B2(n3079), .ZN(n4487)
         );
  AOI22_X1 U4729 ( .A1(n61), .A2(n3393), .B1(n1221), .B2(n33100), .ZN(n4485)
         );
  OAI22_X1 U4730 ( .A1(n2287), .A2(n2994), .B1(n3879), .B2(n2812), .ZN(N162)
         );
  INV_X1 U4731 ( .A(n4488), .ZN(n3879) );
  OAI211_X1 U4732 ( .C1(n2836), .C2(n3014), .A(n4489), .B(n44901), .ZN(n4488)
         );
  AOI221_X1 U4733 ( .B1(n2499), .B2(n28200), .C1(n3185), .C2(n50), .A(n4491), 
        .ZN(n44901) );
  OAI22_X1 U4734 ( .A1(n1025), .A2(n2987), .B1(n2486), .B2(n3067), .ZN(n4491)
         );
  AOI22_X1 U4735 ( .A1(n63), .A2(n29201), .B1(n2744), .B2(n33500), .ZN(n4489)
         );
  OAI22_X1 U4736 ( .A1(n2293), .A2(n29901), .B1(n3881), .B2(n1981), .ZN(N161)
         );
  INV_X1 U4737 ( .A(n4492), .ZN(n3881) );
  OAI211_X1 U4738 ( .C1(n2838), .C2(n552), .A(n4493), .B(n4494), .ZN(n4492) );
  AOI221_X1 U4739 ( .B1(n2489), .B2(n28500), .C1(n31801), .C2(n49), .A(n4495), 
        .ZN(n4494) );
  OAI22_X1 U4740 ( .A1(n2933), .A2(n2983), .B1(n2473), .B2(n3071), .ZN(n4495)
         );
  AOI22_X1 U4741 ( .A1(n65), .A2(n3396), .B1(n2742), .B2(n33900), .ZN(n4493)
         );
  OAI22_X1 U4742 ( .A1(n2289), .A2(n2986), .B1(n3883), .B2(n3343), .ZN(N160)
         );
  INV_X1 U4743 ( .A(n4496), .ZN(n3883) );
  OAI211_X1 U4744 ( .C1(n2832), .C2(n1054), .A(n4497), .B(n4498), .ZN(n4496)
         );
  AOI221_X1 U4745 ( .B1(n2494), .B2(n28800), .C1(n3176), .C2(n48), .A(n4499), 
        .ZN(n4498) );
  OAI22_X1 U4746 ( .A1(n2093), .A2(n29801), .B1(n2501), .B2(n3059), .ZN(n4499)
         );
  AOI22_X1 U4747 ( .A1(n67), .A2(n3389), .B1(n27501), .B2(n34300), .ZN(n4497)
         );
  OAI22_X1 U4748 ( .A1(n2296), .A2(n2982), .B1(n3885), .B2(n3343), .ZN(N159)
         );
  INV_X1 U4749 ( .A(n45001), .ZN(n3885) );
  OAI211_X1 U4750 ( .C1(n2834), .C2(n551), .A(n4501), .B(n4502), .ZN(n45001)
         );
  AOI221_X1 U4751 ( .B1(n2492), .B2(n29100), .C1(n3178), .C2(n47), .A(n4503), 
        .ZN(n4502) );
  OAI22_X1 U4752 ( .A1(n3384), .A2(n2975), .B1(n2503), .B2(n3063), .ZN(n4503)
         );
  AOI22_X1 U4753 ( .A1(n69), .A2(n3237), .B1(n2148), .B2(n34700), .ZN(n4501)
         );
  OAI22_X1 U4754 ( .A1(n2288), .A2(n2978), .B1(n3887), .B2(n1284), .ZN(N158)
         );
  INV_X1 U4755 ( .A(n4504), .ZN(n3887) );
  OAI211_X1 U4756 ( .C1(n2828), .C2(n2175), .A(n4505), .B(n4506), .ZN(n4504)
         );
  AOI221_X1 U4757 ( .B1(n2493), .B2(n29400), .C1(n2721), .C2(n46), .A(n4507), 
        .ZN(n4506) );
  OAI22_X1 U4758 ( .A1(n1028), .A2(n2972), .B1(n2485), .B2(n3051), .ZN(n4507)
         );
  AOI22_X1 U4759 ( .A1(n71), .A2(n2916), .B1(n3426), .B2(n35100), .ZN(n4505)
         );
  OAI22_X1 U4760 ( .A1(n2292), .A2(n2974), .B1(n3889), .B2(n19801), .ZN(N157)
         );
  INV_X1 U4761 ( .A(n4508), .ZN(n3889) );
  OAI211_X1 U4762 ( .C1(n28301), .C2(n1055), .A(n4509), .B(n45101), .ZN(n4508)
         );
  AOI221_X1 U4763 ( .B1(n2499), .B2(n29700), .C1(n3186), .C2(n45), .A(n4511), 
        .ZN(n45101) );
  OAI22_X1 U4764 ( .A1(n2729), .A2(n2968), .B1(n24801), .B2(n3055), .ZN(n4511)
         );
  AOI22_X1 U4765 ( .A1(n73), .A2(n2922), .B1(n1496), .B2(n35500), .ZN(n4509)
         );
  OAI22_X1 U4766 ( .A1(n2289), .A2(n29701), .B1(n3891), .B2(n1683), .ZN(N156)
         );
  INV_X1 U4767 ( .A(n4512), .ZN(n3891) );
  OAI211_X1 U4768 ( .C1(n2824), .C2(n2205), .A(n4513), .B(n4514), .ZN(n4512)
         );
  AOI221_X1 U4769 ( .B1(n25001), .B2(n30000), .C1(n1116), .C2(n44), .A(n4515), 
        .ZN(n4514) );
  OAI22_X1 U4770 ( .A1(n3386), .A2(n2964), .B1(n2479), .B2(n3043), .ZN(n4515)
         );
  AOI22_X1 U4771 ( .A1(n75), .A2(n2924), .B1(n2089), .B2(n35900), .ZN(n4513)
         );
  OAI22_X1 U4772 ( .A1(n2296), .A2(n2966), .B1(n3893), .B2(n1684), .ZN(N155)
         );
  INV_X1 U4773 ( .A(n4516), .ZN(n3893) );
  OAI211_X1 U4774 ( .C1(n2826), .C2(n1053), .A(n4517), .B(n4518), .ZN(n4516)
         );
  AOI221_X1 U4775 ( .B1(n2488), .B2(n30300), .C1(n3181), .C2(n43), .A(n4519), 
        .ZN(n4518) );
  OAI22_X1 U4776 ( .A1(n2733), .A2(n2959), .B1(n2506), .B2(n3047), .ZN(n4519)
         );
  AOI22_X1 U4777 ( .A1(n77), .A2(n2931), .B1(n3023), .B2(n36300), .ZN(n4517)
         );
  OAI22_X1 U4778 ( .A1(n2288), .A2(n2962), .B1(n3895), .B2(n2812), .ZN(N154)
         );
  INV_X1 U4779 ( .A(n45201), .ZN(n3895) );
  OAI211_X1 U4780 ( .C1(n28201), .C2(n2171), .A(n4521), .B(n4522), .ZN(n45201)
         );
  AOI221_X1 U4781 ( .B1(n2488), .B2(n30600), .C1(n3179), .C2(n42), .A(n4523), 
        .ZN(n4522) );
  OAI22_X1 U4782 ( .A1(n2929), .A2(n2955), .B1(n2472), .B2(n3035), .ZN(n4523)
         );
  AOI22_X1 U4783 ( .A1(n79), .A2(n3224), .B1(n2738), .B2(n36700), .ZN(n4521)
         );
  OAI22_X1 U4784 ( .A1(n2293), .A2(n2958), .B1(n3897), .B2(n1981), .ZN(N153)
         );
  INV_X1 U4785 ( .A(n4524), .ZN(n3897) );
  OAI211_X1 U4786 ( .C1(n2822), .C2(n1487), .A(n4525), .B(n4526), .ZN(n4524)
         );
  AOI221_X1 U4787 ( .B1(n2494), .B2(n30900), .C1(n3182), .C2(n41), .A(n4527), 
        .ZN(n4526) );
  OAI22_X1 U4788 ( .A1(n2723), .A2(n2951), .B1(n2482), .B2(n3039), .ZN(n4527)
         );
  AOI22_X1 U4789 ( .A1(n81), .A2(n21001), .B1(n1109), .B2(n37100), .ZN(n4525)
         );
  OAI22_X1 U4790 ( .A1(n22901), .A2(n2954), .B1(n3899), .B2(n1977), .ZN(N152)
         );
  INV_X1 U4791 ( .A(n4528), .ZN(n3899) );
  OAI211_X1 U4792 ( .C1(n2816), .C2(n1473), .A(n4529), .B(n45301), .ZN(n4528)
         );
  AOI221_X1 U4793 ( .B1(n2495), .B2(n31200), .C1(n3187), .C2(n40), .A(n4531), 
        .ZN(n45301) );
  OAI22_X1 U4794 ( .A1(n2932), .A2(n2947), .B1(n2474), .B2(n3027), .ZN(n4531)
         );
  AOI22_X1 U4795 ( .A1(n83), .A2(n3429), .B1(n3378), .B2(n37500), .ZN(n4529)
         );
  OAI22_X1 U4796 ( .A1(n2297), .A2(n29501), .B1(n3901), .B2(n1977), .ZN(N151)
         );
  INV_X1 U4797 ( .A(n4532), .ZN(n3901) );
  OAI211_X1 U4798 ( .C1(n2818), .C2(n1481), .A(n4533), .B(n4534), .ZN(n4532)
         );
  AOI221_X1 U4799 ( .B1(n2493), .B2(n31500), .C1(n1214), .C2(n39), .A(n4535), 
        .ZN(n4534) );
  OAI22_X1 U4800 ( .A1(n2938), .A2(n2944), .B1(n2509), .B2(n3031), .ZN(n4535)
         );
  NAND2_X1 U4801 ( .A1(n1293), .A2(n547), .ZN(n4272) );
  AOI22_X1 U4802 ( .A1(n85), .A2(n3232), .B1(n2748), .B2(n37900), .ZN(n4533)
         );
  OAI22_X1 U4803 ( .A1(n3304), .A2(n1283), .B1(n3241), .B2(n1032), .ZN(n4536)
         );
  NAND2_X1 U4804 ( .A1(n2034), .A2(n3903), .ZN(n44701) );
  INV_X1 U4805 ( .A(n4537), .ZN(n3903) );
  AOI21_X1 U4806 ( .B1(n2212), .B2(n22101), .A(n39401), .ZN(n4537) );
  OAI22_X1 U4807 ( .A1(n2302), .A2(n3149), .B1(n3906), .B2(n1277), .ZN(N150)
         );
  INV_X1 U4808 ( .A(n45401), .ZN(n3906) );
  OAI211_X1 U4809 ( .C1(n563), .C2(n14701), .A(n4541), .B(n4542), .ZN(n45401)
         );
  AOI221_X1 U4810 ( .B1(n3184), .B2(n22100), .C1(n1577), .C2(n26900), .A(n4543), .ZN(n4542) );
  OAI22_X1 U4811 ( .A1(n2875), .A2(n15880), .B1(n3084), .B2(n2733), .ZN(n4543)
         );
  INV_X1 U4812 ( .A(n12100), .ZN(n3762) );
  AOI22_X1 U4813 ( .A1(n2108), .A2(n46300), .B1(n1501), .B2(n15800), .ZN(n4541) );
  INV_X1 U4814 ( .A(n55), .ZN(n3905) );
  OAI22_X1 U4815 ( .A1(n2299), .A2(n3153), .B1(n3909), .B2(n1985), .ZN(N149)
         );
  INV_X1 U4816 ( .A(n4544), .ZN(n3909) );
  OAI211_X1 U4817 ( .C1(n560), .C2(n1201), .A(n4545), .B(n4546), .ZN(n4544) );
  AOI221_X1 U4818 ( .B1(n1514), .B2(n22400), .C1(n15930), .C2(n17), .A(n4547), 
        .ZN(n4546) );
  OAI22_X1 U4819 ( .A1(n2877), .A2(n1606), .B1(n1111), .B2(n3088), .ZN(n4547)
         );
  INV_X1 U4820 ( .A(n12300), .ZN(n3765) );
  AOI22_X1 U4821 ( .A1(n46800), .A2(n2588), .B1(n1501), .B2(n16200), .ZN(n4545) );
  INV_X1 U4822 ( .A(n57), .ZN(n3908) );
  OAI22_X1 U4823 ( .A1(n2309), .A2(n3141), .B1(n3911), .B2(n1087), .ZN(N148)
         );
  INV_X1 U4824 ( .A(n4548), .ZN(n3911) );
  OAI211_X1 U4825 ( .C1(n561), .C2(n2207), .A(n4549), .B(n45501), .ZN(n4548)
         );
  AOI221_X1 U4826 ( .B1(n31801), .B2(n22700), .C1(n3277), .C2(n16), .A(n4551), 
        .ZN(n45501) );
  OAI22_X1 U4827 ( .A1(n2871), .A2(n1064), .B1(n2095), .B2(n3076), .ZN(n4551)
         );
  INV_X1 U4828 ( .A(n12500), .ZN(n3767) );
  AOI22_X1 U4829 ( .A1(n4730), .A2(n2113), .B1(n3026), .B2(n16600), .ZN(n4549)
         );
  INV_X1 U4830 ( .A(n59), .ZN(n39101) );
  OAI22_X1 U4831 ( .A1(n2306), .A2(n3145), .B1(n3913), .B2(n1087), .ZN(N147)
         );
  INV_X1 U4832 ( .A(n4552), .ZN(n3913) );
  OAI211_X1 U4833 ( .C1(n562), .C2(n1197), .A(n4553), .B(n4554), .ZN(n4552) );
  AOI221_X1 U4834 ( .B1(n3409), .B2(n23000), .C1(n1576), .C2(n15), .A(n4555), 
        .ZN(n4554) );
  OAI22_X1 U4835 ( .A1(n2873), .A2(n15870), .B1(n2094), .B2(n30801), .ZN(n4555) );
  INV_X1 U4836 ( .A(n12700), .ZN(n3769) );
  AOI22_X1 U4837 ( .A1(n4780), .A2(n1022), .B1(n20901), .B2(n17000), .ZN(n4553) );
  INV_X1 U4838 ( .A(n61), .ZN(n3912) );
  OAI22_X1 U4839 ( .A1(n2302), .A2(n3133), .B1(n3915), .B2(n2806), .ZN(N146)
         );
  INV_X1 U4840 ( .A(n4556), .ZN(n3915) );
  OAI211_X1 U4841 ( .C1(n567), .C2(n2175), .A(n4557), .B(n4558), .ZN(n4556) );
  AOI221_X1 U4842 ( .B1(n1513), .B2(n23300), .C1(n15971), .C2(n14), .A(n4559), 
        .ZN(n4558) );
  OAI22_X1 U4843 ( .A1(n2867), .A2(n3295), .B1(n2728), .B2(n3068), .ZN(n4559)
         );
  INV_X1 U4844 ( .A(n12900), .ZN(n3771) );
  AOI22_X1 U4845 ( .A1(n4830), .A2(n3394), .B1(n2739), .B2(n17400), .ZN(n4557)
         );
  INV_X1 U4846 ( .A(n63), .ZN(n3914) );
  OAI22_X1 U4847 ( .A1(n23001), .A2(n3137), .B1(n3917), .B2(n1986), .ZN(N145)
         );
  INV_X1 U4848 ( .A(n45601), .ZN(n3917) );
  OAI211_X1 U4849 ( .C1(n564), .C2(n559), .A(n4561), .B(n4562), .ZN(n45601) );
  AOI221_X1 U4850 ( .B1(n3187), .B2(n23600), .C1(n1573), .C2(n13), .A(n4563), 
        .ZN(n4562) );
  OAI22_X1 U4851 ( .A1(n2869), .A2(n15840), .B1(n1025), .B2(n3072), .ZN(n4563)
         );
  INV_X1 U4852 ( .A(n13100), .ZN(n3773) );
  AOI22_X1 U4853 ( .A1(n4880), .A2(n1772), .B1(n1504), .B2(n17800), .ZN(n4561)
         );
  INV_X1 U4854 ( .A(n65), .ZN(n3916) );
  OAI22_X1 U4855 ( .A1(n2308), .A2(n3125), .B1(n3919), .B2(n3344), .ZN(N144)
         );
  INV_X1 U4856 ( .A(n4564), .ZN(n3919) );
  OAI211_X1 U4857 ( .C1(n565), .C2(n1472), .A(n4565), .B(n4566), .ZN(n4564) );
  AOI221_X1 U4858 ( .B1(n3408), .B2(n23900), .C1(n3281), .C2(n12), .A(n4567), 
        .ZN(n4566) );
  OAI22_X1 U4859 ( .A1(n2863), .A2(n3286), .B1(n2729), .B2(n30601), .ZN(n4567)
         );
  INV_X1 U4860 ( .A(n13300), .ZN(n3775) );
  AOI22_X1 U4861 ( .A1(n493), .A2(n2153), .B1(n3377), .B2(n18200), .ZN(n4565)
         );
  INV_X1 U4862 ( .A(n67), .ZN(n3918) );
  OAI22_X1 U4863 ( .A1(n2305), .A2(n3129), .B1(n3921), .B2(n3344), .ZN(N143)
         );
  INV_X1 U4864 ( .A(n4568), .ZN(n3921) );
  OAI211_X1 U4865 ( .C1(n566), .C2(n2699), .A(n4569), .B(n45701), .ZN(n4568)
         );
  AOI221_X1 U4866 ( .B1(n3183), .B2(n24200), .C1(n15960), .C2(n11), .A(n4571), 
        .ZN(n45701) );
  OAI22_X1 U4867 ( .A1(n2865), .A2(n1608), .B1(n1113), .B2(n3064), .ZN(n4571)
         );
  INV_X1 U4868 ( .A(n13500), .ZN(n3777) );
  AOI22_X1 U4869 ( .A1(n498), .A2(n3392), .B1(n2083), .B2(n18600), .ZN(n4569)
         );
  INV_X1 U4870 ( .A(n69), .ZN(n39201) );
  OAI22_X1 U4871 ( .A1(n2303), .A2(n3117), .B1(n3923), .B2(n1278), .ZN(N142)
         );
  INV_X1 U4872 ( .A(n4572), .ZN(n3923) );
  OAI211_X1 U4873 ( .C1(n571), .C2(n1484), .A(n4573), .B(n4574), .ZN(n4572) );
  AOI221_X1 U4874 ( .B1(n3185), .B2(n24500), .C1(n3276), .C2(n10), .A(n4575), 
        .ZN(n4574) );
  OAI22_X1 U4875 ( .A1(n2859), .A2(n3282), .B1(n2737), .B2(n3052), .ZN(n4575)
         );
  INV_X1 U4876 ( .A(n13700), .ZN(n3779) );
  AOI22_X1 U4877 ( .A1(n5030), .A2(n2152), .B1(n1502), .B2(n19000), .ZN(n4573)
         );
  INV_X1 U4878 ( .A(n71), .ZN(n3922) );
  OAI22_X1 U4879 ( .A1(n2299), .A2(n3121), .B1(n3925), .B2(n1985), .ZN(N141)
         );
  INV_X1 U4880 ( .A(n4576), .ZN(n3925) );
  OAI211_X1 U4881 ( .C1(n568), .C2(n552), .A(n4577), .B(n4578), .ZN(n4576) );
  AOI221_X1 U4882 ( .B1(n2721), .B2(n24800), .C1(n1579), .C2(n9), .A(n4579), 
        .ZN(n4578) );
  OAI22_X1 U4883 ( .A1(n2861), .A2(n15900), .B1(n2727), .B2(n3056), .ZN(n4579)
         );
  INV_X1 U4884 ( .A(n13900), .ZN(n3781) );
  AOI22_X1 U4885 ( .A1(n508), .A2(n3238), .B1(n1058), .B2(n19400), .ZN(n4577)
         );
  INV_X1 U4886 ( .A(n73), .ZN(n3924) );
  OAI22_X1 U4887 ( .A1(n2309), .A2(n3109), .B1(n3927), .B2(n1686), .ZN(N140)
         );
  INV_X1 U4888 ( .A(n45801), .ZN(n3927) );
  OAI211_X1 U4889 ( .C1(n569), .C2(n1478), .A(n4581), .B(n4582), .ZN(n45801)
         );
  AOI221_X1 U4890 ( .B1(n3181), .B2(n25100), .C1(n32901), .C2(n8), .A(n4583), 
        .ZN(n4582) );
  OAI22_X1 U4891 ( .A1(n2855), .A2(n3293), .B1(n2734), .B2(n3044), .ZN(n4583)
         );
  INV_X1 U4892 ( .A(n14100), .ZN(n3783) );
  AOI22_X1 U4893 ( .A1(n513), .A2(n2915), .B1(n3382), .B2(n19800), .ZN(n4581)
         );
  INV_X1 U4894 ( .A(n75), .ZN(n3926) );
  OAI22_X1 U4895 ( .A1(n2306), .A2(n3113), .B1(n3929), .B2(n1982), .ZN(N139)
         );
  INV_X1 U4896 ( .A(n4584), .ZN(n3929) );
  OAI211_X1 U4897 ( .C1(n570), .C2(n551), .A(n4585), .B(n4586), .ZN(n4584) );
  AOI221_X1 U4898 ( .B1(n3179), .B2(n25400), .C1(n1571), .C2(n7), .A(n4587), 
        .ZN(n4586) );
  OAI22_X1 U4899 ( .A1(n2857), .A2(n15820), .B1(n2732), .B2(n3048), .ZN(n4587)
         );
  INV_X1 U4900 ( .A(n14300), .ZN(n3785) );
  AOI22_X1 U4901 ( .A1(n518), .A2(n2921), .B1(n2744), .B2(n20200), .ZN(n4585)
         );
  INV_X1 U4902 ( .A(n77), .ZN(n3928) );
  OAI22_X1 U4903 ( .A1(n2303), .A2(n3101), .B1(n3931), .B2(n2806), .ZN(N138)
         );
  INV_X1 U4904 ( .A(n4588), .ZN(n3931) );
  OAI211_X1 U4905 ( .C1(n575), .C2(n1056), .A(n4589), .B(n45901), .ZN(n4588)
         );
  AOI221_X1 U4906 ( .B1(n1215), .B2(n25700), .C1(n32801), .C2(n6), .A(n4591), 
        .ZN(n45901) );
  OAI22_X1 U4907 ( .A1(n2851), .A2(n3283), .B1(n2938), .B2(n3036), .ZN(n4591)
         );
  INV_X1 U4908 ( .A(n14500), .ZN(n3787) );
  AOI22_X1 U4909 ( .A1(n523), .A2(n2926), .B1(n1059), .B2(n20600), .ZN(n4589)
         );
  INV_X1 U4910 ( .A(n79), .ZN(n39301) );
  OAI22_X1 U4911 ( .A1(n23001), .A2(n3105), .B1(n3933), .B2(n1986), .ZN(N137)
         );
  INV_X1 U4912 ( .A(n4592), .ZN(n3933) );
  OAI211_X1 U4913 ( .C1(n572), .C2(n2171), .A(n4593), .B(n4594), .ZN(n4592) );
  AOI221_X1 U4914 ( .B1(n3178), .B2(n26000), .C1(n3289), .C2(n5), .A(n4595), 
        .ZN(n4594) );
  OAI22_X1 U4915 ( .A1(n2853), .A2(n1605), .B1(n2933), .B2(n30401), .ZN(n4595)
         );
  INV_X1 U4916 ( .A(n14700), .ZN(n3789) );
  AOI22_X1 U4917 ( .A1(n528), .A2(n3393), .B1(n2149), .B2(n21000), .ZN(n4593)
         );
  INV_X1 U4918 ( .A(n81), .ZN(n3932) );
  OAI22_X1 U4919 ( .A1(n2308), .A2(n3093), .B1(n3935), .B2(n1982), .ZN(N136)
         );
  INV_X1 U4920 ( .A(n4596), .ZN(n3935) );
  OAI211_X1 U4921 ( .C1(n573), .C2(n3012), .A(n4597), .B(n4598), .ZN(n4596) );
  AOI221_X1 U4922 ( .B1(n3186), .B2(n26300), .C1(n1574), .C2(n4), .A(n4599), 
        .ZN(n4598) );
  OAI22_X1 U4923 ( .A1(n2847), .A2(n15910), .B1(n1028), .B2(n3028), .ZN(n4599)
         );
  INV_X1 U4924 ( .A(n14900), .ZN(n3791) );
  AOI22_X1 U4925 ( .A1(n533), .A2(n3225), .B1(n2086), .B2(n21400), .ZN(n4597)
         );
  INV_X1 U4926 ( .A(n83), .ZN(n3934) );
  OAI22_X1 U4927 ( .A1(n2305), .A2(n3097), .B1(n3937), .B2(n1687), .ZN(N135)
         );
  INV_X1 U4928 ( .A(n46001), .ZN(n3937) );
  OAI211_X1 U4929 ( .C1(n574), .C2(n2204), .A(n4601), .B(n4602), .ZN(n46001)
         );
  AOI221_X1 U4930 ( .B1(n3182), .B2(n26600), .C1(n15801), .C2(n3), .A(n4603), 
        .ZN(n4602) );
  OAI22_X1 U4931 ( .A1(n2849), .A2(n1609), .B1(n2098), .B2(n3032), .ZN(n4603)
         );
  INV_X1 U4932 ( .A(n15100), .ZN(n3793) );
  AOI22_X1 U4933 ( .A1(n538), .A2(n2919), .B1(n1505), .B2(n21800), .ZN(n4601)
         );
  INV_X1 U4934 ( .A(n85), .ZN(n3936) );
  OAI22_X1 U4935 ( .A1(n2523), .A2(n1277), .B1(n3939), .B2(n2946), .ZN(n4604)
         );
  INV_X1 U4936 ( .A(n4605), .ZN(n3939) );
  OAI21_X1 U4937 ( .B1(n1536), .B2(n2694), .A(n3965), .ZN(n4605) );
  NAND2_X1 U4938 ( .A1(n3357), .A2(n18001), .ZN(n4539) );
  INV_X1 U4939 ( .A(n4606), .ZN(n39401) );
  AOI21_X1 U4940 ( .B1(n2695), .B2(n22101), .A(n2217), .ZN(n4606) );
  OAI22_X1 U4941 ( .A1(n2262), .A2(n3004), .B1(n3941), .B2(n1281), .ZN(N134)
         );
  INV_X1 U4942 ( .A(n4608), .ZN(n3941) );
  OAI211_X1 U4943 ( .C1(n1469), .C2(n2174), .A(n4609), .B(n46101), .ZN(n4608)
         );
  AOI221_X1 U4944 ( .B1(n3287), .B2(n12200), .C1(n1856), .C2(n18), .A(n4612), 
        .ZN(n46101) );
  OAI22_X1 U4945 ( .A1(n1181), .A2(n2465), .B1(n985), .B2(n15830), .ZN(n4612)
         );
  INV_X1 U4946 ( .A(n34), .ZN(n3797) );
  INV_X1 U4947 ( .A(quantized_data[63]), .ZN(n3833) );
  AOI22_X1 U4948 ( .A1(n1524), .A2(n38400), .B1(n2089), .B2(n56), .ZN(n4609)
         );
  INV_X1 U4949 ( .A(n15700), .ZN(n3869) );
  OAI22_X1 U4950 ( .A1(n22701), .A2(n30001), .B1(n3943), .B2(n1975), .ZN(N133)
         );
  INV_X1 U4951 ( .A(n4613), .ZN(n3943) );
  OAI211_X1 U4952 ( .C1(n1462), .C2(n2174), .A(n4614), .B(n4615), .ZN(n4613)
         );
  AOI221_X1 U4953 ( .B1(n3277), .B2(n12400), .C1(n1855), .C2(n27200), .A(n4616), .ZN(n4615) );
  OAI22_X1 U4954 ( .A1(n1184), .A2(n2434), .B1(n986), .B2(n3283), .ZN(n4616)
         );
  INV_X1 U4955 ( .A(n33), .ZN(n38001) );
  INV_X1 U4956 ( .A(quantized_data[62]), .ZN(n3836) );
  AOI22_X1 U4957 ( .A1(n38900), .A2(n1026), .B1(n1224), .B2(n58), .ZN(n4614)
         );
  INV_X1 U4958 ( .A(n16100), .ZN(n3872) );
  OAI22_X1 U4959 ( .A1(n2268), .A2(n2996), .B1(n3945), .B2(n1085), .ZN(N132)
         );
  INV_X1 U4960 ( .A(n4617), .ZN(n3945) );
  OAI211_X1 U4961 ( .C1(n1455), .C2(n2208), .A(n4618), .B(n4619), .ZN(n4617)
         );
  AOI221_X1 U4962 ( .B1(n3279), .B2(n12600), .C1(n1853), .C2(n27500), .A(
        n46201), .ZN(n4619) );
  OAI22_X1 U4963 ( .A1(n1175), .A2(n2468), .B1(n983), .B2(n3294), .ZN(n46201)
         );
  INV_X1 U4964 ( .A(n32), .ZN(n3802) );
  INV_X1 U4965 ( .A(quantized_data[61]), .ZN(n3838) );
  AOI22_X1 U4966 ( .A1(n39400), .A2(n29301), .B1(n2746), .B2(n60), .ZN(n4618)
         );
  INV_X1 U4967 ( .A(n16500), .ZN(n3874) );
  INV_X1 U4968 ( .A(n4710), .ZN(n3944) );
  OAI22_X1 U4969 ( .A1(n2275), .A2(n2992), .B1(n3946), .B2(n1085), .ZN(N131)
         );
  INV_X1 U4970 ( .A(n4621), .ZN(n3946) );
  OAI211_X1 U4971 ( .C1(n1448), .C2(n1475), .A(n4622), .B(n4623), .ZN(n4621)
         );
  AOI221_X1 U4972 ( .B1(n15930), .B2(n12800), .C1(n1852), .C2(n27800), .A(
        n4624), .ZN(n4623) );
  OAI22_X1 U4973 ( .A1(n1178), .A2(n2427), .B1(n984), .B2(n1064), .ZN(n4624)
         );
  INV_X1 U4974 ( .A(n31), .ZN(n3804) );
  INV_X1 U4975 ( .A(quantized_data[60]), .ZN(n38401) );
  AOI22_X1 U4976 ( .A1(n39900), .A2(n2156), .B1(n2746), .B2(n62), .ZN(n4622)
         );
  INV_X1 U4977 ( .A(n16900), .ZN(n3876) );
  OAI22_X1 U4978 ( .A1(n2262), .A2(n2988), .B1(n3947), .B2(n28101), .ZN(N130)
         );
  INV_X1 U4979 ( .A(n4625), .ZN(n3947) );
  OAI211_X1 U4980 ( .C1(n1443), .C2(n2172), .A(n4626), .B(n4627), .ZN(n4625)
         );
  AOI221_X1 U4981 ( .B1(n1572), .B2(n13000), .C1(n1849), .C2(n28100), .A(n4628), .ZN(n4627) );
  OAI22_X1 U4982 ( .A1(n1169), .A2(n2459), .B1(n981), .B2(n3284), .ZN(n4628)
         );
  INV_X1 U4983 ( .A(n30), .ZN(n3806) );
  INV_X1 U4984 ( .A(quantized_data[59]), .ZN(n3842) );
  AOI22_X1 U4985 ( .A1(n40400), .A2(n2153), .B1(n1493), .B2(n64), .ZN(n4626)
         );
  INV_X1 U4986 ( .A(n17300), .ZN(n3878) );
  OAI22_X1 U4987 ( .A1(n2271), .A2(n2984), .B1(n3948), .B2(n1976), .ZN(N129)
         );
  INV_X1 U4988 ( .A(n4629), .ZN(n3948) );
  OAI211_X1 U4989 ( .C1(n1436), .C2(n2172), .A(n46301), .B(n4631), .ZN(n4629)
         );
  AOI221_X1 U4990 ( .B1(n32801), .B2(n13200), .C1(n16320), .C2(n28400), .A(
        n4632), .ZN(n4631) );
  OAI22_X1 U4991 ( .A1(n1172), .A2(n24301), .B1(n982), .B2(n3293), .ZN(n4632)
         );
  INV_X1 U4992 ( .A(n29), .ZN(n3808) );
  INV_X1 U4993 ( .A(quantized_data[58]), .ZN(n3844) );
  AOI22_X1 U4994 ( .A1(n40900), .A2(n3236), .B1(n3022), .B2(n66), .ZN(n46301)
         );
  INV_X1 U4995 ( .A(n17700), .ZN(n38801) );
  OAI22_X1 U4996 ( .A1(n2267), .A2(n1044), .B1(n39501), .B2(n3342), .ZN(N128)
         );
  INV_X1 U4997 ( .A(n4633), .ZN(n39501) );
  OAI211_X1 U4998 ( .C1(n1429), .C2(n2204), .A(n4634), .B(n4635), .ZN(n4633)
         );
  AOI221_X1 U4999 ( .B1(n15940), .B2(n13400), .C1(n1849), .C2(n28700), .A(
        n4636), .ZN(n4635) );
  OAI22_X1 U5000 ( .A1(n1163), .A2(n2463), .B1(n979), .B2(n15840), .ZN(n4636)
         );
  INV_X1 U5001 ( .A(n28), .ZN(n38101) );
  INV_X1 U5002 ( .A(quantized_data[57]), .ZN(n3846) );
  AOI22_X1 U5003 ( .A1(n41400), .A2(n3232), .B1(n14901), .B2(n68), .ZN(n4634)
         );
  INV_X1 U5004 ( .A(n18100), .ZN(n3882) );
  INV_X1 U5005 ( .A(n4910), .ZN(n3949) );
  OAI22_X1 U5006 ( .A1(n2274), .A2(n2976), .B1(n3951), .B2(n3342), .ZN(N127)
         );
  INV_X1 U5007 ( .A(n4637), .ZN(n3951) );
  OAI211_X1 U5008 ( .C1(n1422), .C2(n2208), .A(n4638), .B(n4639), .ZN(n4637)
         );
  AOI221_X1 U5009 ( .B1(n3276), .B2(n13600), .C1(n16330), .C2(n29000), .A(
        n46401), .ZN(n4639) );
  OAI22_X1 U5010 ( .A1(n1166), .A2(n2425), .B1(n980), .B2(n15870), .ZN(n46401)
         );
  INV_X1 U5011 ( .A(n27), .ZN(n3812) );
  INV_X1 U5012 ( .A(quantized_data[56]), .ZN(n3848) );
  AOI22_X1 U5013 ( .A1(n41900), .A2(n1023), .B1(n27501), .B2(n70), .ZN(n4638)
         );
  INV_X1 U5014 ( .A(n18500), .ZN(n3884) );
  OAI22_X1 U5015 ( .A1(n2263), .A2(n1041), .B1(n3953), .B2(n1282), .ZN(N126)
         );
  INV_X1 U5016 ( .A(n4641), .ZN(n3953) );
  OAI211_X1 U5017 ( .C1(n1417), .C2(n2708), .A(n4642), .B(n4643), .ZN(n4641)
         );
  AOI221_X1 U5018 ( .B1(n1579), .B2(n13800), .C1(n1855), .C2(n29300), .A(n4644), .ZN(n4643) );
  OAI22_X1 U5019 ( .A1(n1157), .A2(n2466), .B1(n977), .B2(n1608), .ZN(n4644)
         );
  INV_X1 U5020 ( .A(n26), .ZN(n3814) );
  INV_X1 U5021 ( .A(quantized_data[55]), .ZN(n38501) );
  AOI22_X1 U5022 ( .A1(n42400), .A2(n1024), .B1(n3379), .B2(n72), .ZN(n4642)
         );
  INV_X1 U5023 ( .A(n18900), .ZN(n3886) );
  INV_X1 U5024 ( .A(n5010), .ZN(n3952) );
  OAI22_X1 U5025 ( .A1(n22701), .A2(n1039), .B1(n3955), .B2(n1975), .ZN(N125)
         );
  INV_X1 U5026 ( .A(n4645), .ZN(n3955) );
  OAI211_X1 U5027 ( .C1(n14101), .C2(n1484), .A(n4646), .B(n4647), .ZN(n4645)
         );
  AOI221_X1 U5028 ( .B1(n15960), .B2(n14000), .C1(n1853), .C2(n29600), .A(
        n4648), .ZN(n4647) );
  OAI22_X1 U5029 ( .A1(n11601), .A2(n2435), .B1(n978), .B2(n3282), .ZN(n4648)
         );
  INV_X1 U5030 ( .A(n25), .ZN(n3816) );
  INV_X1 U5031 ( .A(quantized_data[54]), .ZN(n3852) );
  AOI22_X1 U5032 ( .A1(n42900), .A2(n2101), .B1(n1495), .B2(n74), .ZN(n4646)
         );
  INV_X1 U5033 ( .A(n19300), .ZN(n3888) );
  INV_X1 U5034 ( .A(n506), .ZN(n3954) );
  OAI22_X1 U5035 ( .A1(n2267), .A2(n1037), .B1(n3957), .B2(n16801), .ZN(N124)
         );
  INV_X1 U5036 ( .A(n4649), .ZN(n3957) );
  OAI211_X1 U5037 ( .C1(n1405), .C2(n1197), .A(n46501), .B(n4651), .ZN(n4649)
         );
  AOI221_X1 U5038 ( .B1(n1573), .B2(n14200), .C1(n1069), .C2(n29900), .A(n4652), .ZN(n4651) );
  OAI22_X1 U5039 ( .A1(n1151), .A2(n2469), .B1(n975), .B2(n3286), .ZN(n4652)
         );
  INV_X1 U5040 ( .A(n24), .ZN(n3818) );
  INV_X1 U5041 ( .A(quantized_data[53]), .ZN(n3854) );
  AOI22_X1 U5042 ( .A1(n43400), .A2(n1525), .B1(n3015), .B2(n76), .ZN(n46501)
         );
  INV_X1 U5043 ( .A(n19700), .ZN(n38901) );
  INV_X1 U5044 ( .A(n511), .ZN(n3956) );
  OAI22_X1 U5045 ( .A1(n2274), .A2(n29601), .B1(n3958), .B2(n1972), .ZN(N123)
         );
  INV_X1 U5046 ( .A(n4653), .ZN(n3958) );
  OAI211_X1 U5047 ( .C1(n14001), .C2(n1478), .A(n4654), .B(n4655), .ZN(n4653)
         );
  AOI221_X1 U5048 ( .B1(n1576), .B2(n14400), .C1(n1069), .C2(n30200), .A(n4656), .ZN(n4655) );
  OAI22_X1 U5049 ( .A1(n1154), .A2(n2428), .B1(n976), .B2(n1605), .ZN(n4656)
         );
  INV_X1 U5050 ( .A(n23), .ZN(n38201) );
  INV_X1 U5051 ( .A(quantized_data[52]), .ZN(n3856) );
  AOI22_X1 U5052 ( .A1(n43900), .A2(n2917), .B1(n550), .B2(n78), .ZN(n4654) );
  INV_X1 U5053 ( .A(n20100), .ZN(n3892) );
  OAI22_X1 U5054 ( .A1(n2263), .A2(n2956), .B1(n3959), .B2(n28101), .ZN(N122)
         );
  INV_X1 U5055 ( .A(n4657), .ZN(n3959) );
  OAI211_X1 U5056 ( .C1(n1395), .C2(n683), .A(n4658), .B(n4659), .ZN(n4657) );
  AOI221_X1 U5057 ( .B1(n3289), .B2(n14600), .C1(n1856), .C2(n30500), .A(
        n46601), .ZN(n4659) );
  OAI22_X1 U5058 ( .A1(n1145), .A2(n24601), .B1(n973), .B2(n15850), .ZN(n46601) );
  INV_X1 U5059 ( .A(n22), .ZN(n3822) );
  INV_X1 U5060 ( .A(quantized_data[51]), .ZN(n3858) );
  AOI22_X1 U5061 ( .A1(n44400), .A2(n2108), .B1(n2741), .B2(n80), .ZN(n4658)
         );
  INV_X1 U5062 ( .A(n20500), .ZN(n3894) );
  OAI22_X1 U5063 ( .A1(n2271), .A2(n2952), .B1(n39601), .B2(n1976), .ZN(N121)
         );
  INV_X1 U5064 ( .A(n4661), .ZN(n39601) );
  OAI211_X1 U5065 ( .C1(n1388), .C2(n1487), .A(n4662), .B(n4663), .ZN(n4661)
         );
  AOI221_X1 U5066 ( .B1(n1571), .B2(n14800), .C1(n1852), .C2(n30800), .A(n4664), .ZN(n4663) );
  OAI22_X1 U5067 ( .A1(n1148), .A2(n2429), .B1(n974), .B2(n15900), .ZN(n4664)
         );
  INV_X1 U5068 ( .A(n21), .ZN(n3824) );
  INV_X1 U5069 ( .A(quantized_data[50]), .ZN(n38601) );
  AOI22_X1 U5070 ( .A1(n44900), .A2(n2151), .B1(n3375), .B2(n82), .ZN(n4662)
         );
  INV_X1 U5071 ( .A(n20900), .ZN(n3896) );
  OAI22_X1 U5072 ( .A1(n2268), .A2(n2948), .B1(n3962), .B2(n1972), .ZN(N120)
         );
  INV_X1 U5073 ( .A(n4665), .ZN(n3962) );
  OAI211_X1 U5074 ( .C1(n1381), .C2(n2205), .A(n4666), .B(n4667), .ZN(n4665)
         );
  AOI221_X1 U5075 ( .B1(n3281), .B2(n15000), .C1(n3326), .C2(n31100), .A(n4668), .ZN(n4667) );
  OAI22_X1 U5076 ( .A1(n1139), .A2(n2462), .B1(n971), .B2(n3295), .ZN(n4668)
         );
  INV_X1 U5077 ( .A(n20), .ZN(n3826) );
  INV_X1 U5078 ( .A(quantized_data[49]), .ZN(n3862) );
  AOI22_X1 U5079 ( .A1(n45400), .A2(n15301), .B1(n1222), .B2(n84), .ZN(n4666)
         );
  INV_X1 U5080 ( .A(n21300), .ZN(n3898) );
  INV_X1 U5081 ( .A(n531), .ZN(n3961) );
  OAI22_X1 U5082 ( .A1(n2275), .A2(n2945), .B1(n3963), .B2(n1681), .ZN(N119)
         );
  INV_X1 U5083 ( .A(n4669), .ZN(n3963) );
  OAI211_X1 U5084 ( .C1(n1374), .C2(n1481), .A(n46701), .B(n4671), .ZN(n4669)
         );
  AOI221_X1 U5085 ( .B1(n32901), .B2(n15200), .C1(n3326), .C2(n31400), .A(
        n4672), .ZN(n4671) );
  OAI22_X1 U5086 ( .A1(n1142), .A2(n2424), .B1(n972), .B2(n15820), .ZN(n4672)
         );
  NOR2_X1 U5087 ( .A1(n11301), .A2(n32701), .ZN(n4188) );
  INV_X1 U5088 ( .A(n19), .ZN(n3828) );
  INV_X1 U5089 ( .A(quantized_data[48]), .ZN(n3864) );
  NOR2_X1 U5090 ( .A1(n1232), .A2(n15550), .ZN(n4189) );
  AOI22_X1 U5091 ( .A1(n45900), .A2(n3398), .B1(n2148), .B2(n86), .ZN(n46701)
         );
  INV_X1 U5092 ( .A(n1234), .ZN(n4119) );
  NAND2_X1 U5093 ( .A1(n3302), .A2(n1136), .ZN(n4139) );
  NAND2_X1 U5094 ( .A1(n2679), .A2(n546), .ZN(n4194) );
  NOR2_X1 U5095 ( .A1(n3216), .A2(n1617), .ZN(n4118) );
  NAND2_X1 U5096 ( .A1(n3212), .A2(n2215), .ZN(n41401) );
  INV_X1 U5097 ( .A(n21700), .ZN(n39001) );
  OAI22_X1 U5098 ( .A1(n25301), .A2(n1281), .B1(n586), .B2(n1369), .ZN(n4674)
         );
  NAND2_X1 U5099 ( .A1(n2535), .A2(n1117), .ZN(n3965) );
  NAND2_X1 U5100 ( .A1(n1096), .A2(n3966), .ZN(n4607) );
  NAND2_X1 U5101 ( .A1(n4676), .A2(n4677), .ZN(n3966) );
  NAND3_X1 U5102 ( .A1(n2695), .A2(n2211), .A3(n2209), .ZN(n4677) );
  NAND2_X1 U5103 ( .A1(n1288), .A2(n1242), .ZN(n3758) );
  NOR2_X1 U5104 ( .A1(n1537), .A2(n548), .ZN(n4673) );
  OAI22_X1 U5105 ( .A1(n3968), .A2(n2219), .B1(n3086), .B2(n1911), .ZN(N118)
         );
  INV_X1 U5106 ( .A(n38100), .ZN(n3969) );
  INV_X1 U5107 ( .A(N939), .ZN(n3968) );
  OAI22_X1 U5108 ( .A1(n3971), .A2(n2224), .B1(n30901), .B2(n1908), .ZN(N117)
         );
  INV_X1 U5109 ( .A(n38600), .ZN(n3972) );
  INV_X1 U5110 ( .A(N938), .ZN(n3971) );
  OAI22_X1 U5111 ( .A1(n3973), .A2(n2223), .B1(n3078), .B2(n3333), .ZN(N116)
         );
  INV_X1 U5112 ( .A(n39100), .ZN(n3974) );
  INV_X1 U5113 ( .A(N937), .ZN(n3973) );
  OAI22_X1 U5114 ( .A1(n3975), .A2(n2228), .B1(n3082), .B2(n3333), .ZN(N115)
         );
  INV_X1 U5115 ( .A(n39600), .ZN(n3976) );
  INV_X1 U5116 ( .A(N936), .ZN(n3975) );
  OAI22_X1 U5117 ( .A1(n3977), .A2(n2219), .B1(n30701), .B2(n1911), .ZN(N114)
         );
  INV_X1 U5118 ( .A(n40100), .ZN(n3978) );
  INV_X1 U5119 ( .A(N935), .ZN(n3977) );
  OAI22_X1 U5120 ( .A1(n3979), .A2(n2225), .B1(n3074), .B2(n1909), .ZN(N113)
         );
  INV_X1 U5121 ( .A(n40600), .ZN(n39801) );
  INV_X1 U5122 ( .A(N934), .ZN(n3979) );
  OAI22_X1 U5123 ( .A1(n3981), .A2(n2222), .B1(n3062), .B2(n1076), .ZN(N112)
         );
  INV_X1 U5124 ( .A(n41100), .ZN(n3982) );
  INV_X1 U5125 ( .A(N933), .ZN(n3981) );
  OAI22_X1 U5126 ( .A1(n3983), .A2(n2227), .B1(n3066), .B2(n1076), .ZN(N111)
         );
  INV_X1 U5127 ( .A(n41600), .ZN(n3984) );
  INV_X1 U5128 ( .A(N932), .ZN(n3983) );
  OAI22_X1 U5129 ( .A1(n3985), .A2(n22201), .B1(n3054), .B2(n1912), .ZN(N110)
         );
  INV_X1 U5130 ( .A(n42100), .ZN(n3986) );
  INV_X1 U5131 ( .A(N931), .ZN(n3985) );
  OAI22_X1 U5132 ( .A1(n3987), .A2(n2224), .B1(n3058), .B2(n1908), .ZN(N109)
         );
  INV_X1 U5133 ( .A(n42600), .ZN(n3988) );
  INV_X1 U5134 ( .A(N930), .ZN(n3987) );
  OAI22_X1 U5135 ( .A1(n3989), .A2(n2222), .B1(n3046), .B2(n1905), .ZN(N108)
         );
  INV_X1 U5136 ( .A(n43100), .ZN(n39901) );
  INV_X1 U5137 ( .A(N929), .ZN(n3989) );
  OAI22_X1 U5138 ( .A1(n3991), .A2(n2227), .B1(n30501), .B2(n1905), .ZN(N107)
         );
  INV_X1 U5139 ( .A(n43600), .ZN(n3992) );
  INV_X1 U5140 ( .A(N928), .ZN(n3991) );
  OAI22_X1 U5141 ( .A1(n3993), .A2(n22201), .B1(n3038), .B2(n1912), .ZN(N106)
         );
  INV_X1 U5142 ( .A(n44100), .ZN(n3994) );
  INV_X1 U5143 ( .A(N927), .ZN(n3993) );
  OAI22_X1 U5144 ( .A1(n3995), .A2(n2225), .B1(n3042), .B2(n1909), .ZN(N105)
         );
  INV_X1 U5145 ( .A(n44600), .ZN(n3996) );
  INV_X1 U5146 ( .A(N926), .ZN(n3995) );
  OAI22_X1 U5147 ( .A1(n3997), .A2(n2223), .B1(n30301), .B2(n1653), .ZN(N104)
         );
  INV_X1 U5148 ( .A(n45100), .ZN(n3998) );
  INV_X1 U5149 ( .A(N925), .ZN(n3997) );
  OAI22_X1 U5150 ( .A1(n3999), .A2(n2228), .B1(n3034), .B2(n1654), .ZN(N103)
         );
  NOR2_X1 U5151 ( .A1(n11301), .A2(n1538), .ZN(n4001) );
  NOR2_X1 U5152 ( .A1(n26901), .A2(n9250), .ZN(n4675) );
  INV_X1 U5153 ( .A(n45600), .ZN(n40001) );
  NAND2_X1 U5154 ( .A1(n1096), .A2(n2216), .ZN(n4678) );
  NOR4_X1 U5155 ( .A1(n543), .A2(n2913), .A3(n2), .A4(n1), .ZN(n4676) );
  INV_X1 U5156 ( .A(N924), .ZN(n3999) );
  OAI211_X1 U5157 ( .C1(n2691), .C2(n1132), .A(n588), .B(n4682), .ZN(N101) );
  MUX2_X1 U5158 ( .A(n1133), .B(n1803), .S(n46801), .Z(n4682) );
  NOR2_X1 U5159 ( .A1(n4684), .A2(data_set[1]), .ZN(n46801) );
  INV_X1 U5160 ( .A(data_set[0]), .ZN(n4684) );
  AND2_X1 U5161 ( .A1(srstn), .A2(sram_write_enable), .ZN(n4681) );
  NOR2_X1 U5162 ( .A1(data_set[1]), .A2(data_set[0]), .ZN(n4683) );
endmodule


module tpu_top ( clk, srstn, tpu_start, sram_rdata_w0, sram_rdata_w1, 
        sram_rdata_d0, sram_rdata_d1, sram_raddr_w0, sram_raddr_w1, 
        sram_raddr_d0, sram_raddr_d1, sram_write_enable_a0, sram_wdata_a, 
        sram_waddr_a, sram_write_enable_b0, sram_wdata_b, sram_waddr_b, 
        sram_write_enable_c0, sram_wdata_c, sram_waddr_c, tpu_done );
  input [31:0] sram_rdata_w0;
  input [31:0] sram_rdata_w1;
  input [31:0] sram_rdata_d0;
  input [31:0] sram_rdata_d1;
  output [9:0] sram_raddr_w0;
  output [9:0] sram_raddr_w1;
  output [9:0] sram_raddr_d0;
  output [9:0] sram_raddr_d1;
  output [127:0] sram_wdata_a;
  output [5:0] sram_waddr_a;
  output [127:0] sram_wdata_b;
  output [5:0] sram_waddr_b;
  output [127:0] sram_wdata_c;
  output [5:0] sram_waddr_c;
  input clk, srstn, tpu_start;
  output sram_write_enable_a0, sram_write_enable_b0, sram_write_enable_c0,
         tpu_done;
  wire   alu_start, sram_write_enable, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, SYNOPSYS_UNCONNECTED_1, SYNOPSYS_UNCONNECTED_2,
         SYNOPSYS_UNCONNECTED_3, SYNOPSYS_UNCONNECTED_4,
         SYNOPSYS_UNCONNECTED_5, SYNOPSYS_UNCONNECTED_6,
         SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8,
         SYNOPSYS_UNCONNECTED_9, SYNOPSYS_UNCONNECTED_10,
         SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12;
  wire   [6:0] addr_serial_num;
  wire   [167:0] ori_data;
  wire   [127:0] quantized_data;
  wire   [8:0] cycle_num;
  wire   [5:0] matrix_index;
  wire   [1:0] data_set;

  addr_sel addr_sel ( .clk(clk), .addr_serial_num({addr_serial_num[6:5], n25, 
        n26, addr_serial_num[2:0]}), .sram_raddr_w0({SYNOPSYS_UNCONNECTED_1, 
        SYNOPSYS_UNCONNECTED_2, SYNOPSYS_UNCONNECTED_3, sram_raddr_w0[6:0]}), 
        .sram_raddr_w1({SYNOPSYS_UNCONNECTED_4, SYNOPSYS_UNCONNECTED_5, 
        SYNOPSYS_UNCONNECTED_6, sram_raddr_w1[6:0]}), .sram_raddr_d0({
        SYNOPSYS_UNCONNECTED_7, SYNOPSYS_UNCONNECTED_8, SYNOPSYS_UNCONNECTED_9, 
        sram_raddr_d0[6:0]}), .sram_raddr_d1({SYNOPSYS_UNCONNECTED_10, 
        SYNOPSYS_UNCONNECTED_11, SYNOPSYS_UNCONNECTED_12, sram_raddr_d1[6:0]})
         );
  quantize_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8_OUTPUT_DATA_WIDTH16 quantize ( 
        .ori_data(ori_data), .quantized_data(quantized_data) );
  systolic_ARRAY_SIZE8_SRAM_DATA_WIDTH32_DATA_WIDTH8 systolic ( .clk(clk), 
        .srstn(n32), .alu_start(alu_start), .cycle_num(cycle_num), 
        .sram_rdata_w0(sram_rdata_w0), .sram_rdata_w1(sram_rdata_w1), 
        .sram_rdata_d0(sram_rdata_d0), .sram_rdata_d1(sram_rdata_d1), 
        .matrix_index({matrix_index[5:3], n27, matrix_index[1:0]}), 
        .mul_outcome(ori_data) );
  systolic_controll_ARRAY_SIZE8 systolic_controll ( .clk(clk), .srstn(n30), 
        .tpu_start(n29), .sram_write_enable(sram_write_enable), 
        .addr_serial_num(addr_serial_num), .alu_start(alu_start), .cycle_num(
        cycle_num), .matrix_index(matrix_index), .data_set(data_set), 
        .tpu_done(tpu_done) );
  write_out_ARRAY_SIZE8_OUTPUT_DATA_WIDTH16 write_out ( .clk(clk), .srstn(n33), 
        .sram_write_enable(sram_write_enable), .data_set(data_set), 
        .matrix_index({matrix_index[5:3], n28, matrix_index[1:0]}), 
        .quantized_data(quantized_data), .sram_write_enable_a0(
        sram_write_enable_a0), .sram_wdata_a(sram_wdata_a), .sram_waddr_a(
        sram_waddr_a), .sram_write_enable_b0(sram_write_enable_b0), 
        .sram_wdata_b(sram_wdata_b), .sram_waddr_b(sram_waddr_b), 
        .sram_write_enable_c0(sram_write_enable_c0), .sram_wdata_c(
        sram_wdata_c), .sram_waddr_c(sram_waddr_c) );
  INV_X1 U1 ( .A(1'b1), .ZN(sram_raddr_d1[7]) );
  INV_X1 U3 ( .A(1'b1), .ZN(sram_raddr_d1[8]) );
  INV_X1 U5 ( .A(1'b1), .ZN(sram_raddr_d1[9]) );
  INV_X1 U7 ( .A(1'b1), .ZN(sram_raddr_d0[7]) );
  INV_X1 U9 ( .A(1'b1), .ZN(sram_raddr_d0[8]) );
  INV_X1 U11 ( .A(1'b1), .ZN(sram_raddr_d0[9]) );
  INV_X1 U13 ( .A(1'b1), .ZN(sram_raddr_w1[7]) );
  INV_X1 U15 ( .A(1'b1), .ZN(sram_raddr_w1[8]) );
  INV_X1 U17 ( .A(1'b1), .ZN(sram_raddr_w1[9]) );
  INV_X1 U19 ( .A(1'b1), .ZN(sram_raddr_w0[7]) );
  INV_X1 U21 ( .A(1'b1), .ZN(sram_raddr_w0[8]) );
  INV_X1 U23 ( .A(1'b1), .ZN(sram_raddr_w0[9]) );
  BUF_X1 U25 ( .A(addr_serial_num[4]), .Z(n25) );
  BUF_X1 U26 ( .A(addr_serial_num[3]), .Z(n26) );
  BUF_X1 U27 ( .A(matrix_index[2]), .Z(n27) );
  BUF_X1 U28 ( .A(matrix_index[2]), .Z(n28) );
  CLKBUF_X1 U29 ( .A(tpu_start), .Z(n29) );
  CLKBUF_X1 U30 ( .A(srstn), .Z(n30) );
  INV_X1 U31 ( .A(srstn), .ZN(n31) );
  INV_X1 U32 ( .A(n31), .ZN(n32) );
  INV_X1 U33 ( .A(n31), .ZN(n33) );
endmodule

